��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��e�ik3�������w$����g|��J^]��)�[H<Y��O�h����	�O�_b�[ջ
�l�s+d��N9EP����N] ~�������[�k���;&�(�f�˥|��X%�8!��cYUc<���������F�Ʊj-�����Kx��jj�m.��ތf>�?�5w���e�Z$����)\{-��7� ��;p�������N��,R��X��<�z'0w�����E��e�y.$c��8�f����OY�I��p��4Q�"6?��h�8eEL�pN�� I�|���iD��Ut�w�+����|�> 8ACT���f济$�ߓ��Mldi�
�T:�^�PL�Z�c�f�ѡ�8%mW��f�t�b�'F��c�k�mH*Ӓ?Z�)�S>X9g���Α#j�P��`�6<l��\�K��-�
����3�`V?�	tS�B������$xg(v.��E�me�,����k���0� ���8q��;�^&,�+��O`5����u8�1�a���Tw9��������Ǆ�|�y5?\7/D=	^�p�$ޕ�7y �B���N�nL�k\�"�q��[��� �)���!BA����x���u1�p�L���j�vrƏ��ѽ<LRD���,�"��!�5
Fe��%1-t]�����U��o����9Pp�R��*bGF'����Ցo*̟<��f�\���&6���Bd�R�ݓn����r� ��������dR�a(h�$�D)d���a��%��t#O�`�m{��y؊�5�%[�)�q(Q��SGC�ܑQ������@eo~�~ՌL%|����@{��_�\H>,|6����m��9P��,���ޖA�6Eb�i������^�����wX������q�=��9��-�m��և�"��rf�����lFh���5m��������'&�F�?:%Ռ��!��OA�a��cQ��6�A+Q�Д�H���5��\�I$㲆�w�Oų�b�z<�.˳���/ �}���ɑ�d����i@���*b��K3�ڪ@��ϼ)|QMS�= �y"4����SX$/Q��6�,�%���b�Iv�k3z�|P��T�Kr�jBW�u�2�47WD�3�w�?�'̌ �HН�@��g�E�F����\���QV������&u�2&����e�gv���ʺ��瑓O �[<��[+��I��i�8>@��w�0�t�GUs��
��pLS��|׌VJ�� [����c�hS"���"IwL`���K���^�v��Kb#-�;@<?�ctQ�Ui��6H��*F_7�cOD3-�p���X\5�OX�Rj���q�'r�
ž���Sߝ*�L߅/��7��$K���XU�4�V�
����(��	RǞp�&0���&�J7��6pQ)c3��[��A�z�Z�k�rk�?DH �p�|>�p�;�t�(4'�ZEХ��RG���P����u�Ú�Xd!,T+y��1�c.Q��R�W�Lp�C�2�r���[���g-�c
�Wg:��{�zs�-w�-R�r�ղ�� pwa�ejӼ�Ƥ�='�>*���9��!����<a��
ŞB4�X�-L���#��u�	��	�)�	�y<{�+�=�#gD� ���ذ�|�?P>ވ�I!�G��E�)�E]��r^uv��%��������P%�{:�)'�;�2�%p��4�/��<�Ό�|�u^�u�6��/��P�V����)T�^cY���j�1R3$i$���� ��]�٦�"!/:��ny���>+%�$���2���;�"���A+ Փ�I^���6]�|x��M	7�e��7�%W9���O2O�F�N��ܐFbx�e	��!�Yr/���)����N��a,x>	 m�:�h��%�މ&X�V�c�nPP�_���4l�e^�@��0��ݰ%�Dl9<����W�۞j�ú�(B�1���s�9�
�g��ܚ_)@��A6	T)]d`��L��=��m���En�'���Z�+�<d@��˸����2PZ��פ�iQ�>�N�K�1��fe��-���=��1u�ݪ�\�'���䅯��
�jiV���5�=��]�(���/9���aRC�C��=t�Kx�l�Τ�-Vc�%K�{`�U�!r�ۻ�sekV���\c읫��e��XS�f�0+������	��vL�ܬ��䩩����K�o�����Whi8�����:�qi�����
��
�OsS�/�+!{�Ё�2��<b� �4��qK7��g��O@䦑m 2������k���wU�q�X>
��yԮ?����5Qy�O��Z�F����'���NB��"7�qk��B~/4έ����l�
vԫ�P\]���b#�5�%`�q$����꼳�-h��p�ͻޝ=�� �}������c�XF*�;�=�~JEv�><"Ʋ��ȑ*6�[���?�+]l�a��$Zh�ԅ�!gHYL�@k��_"��y���f�ڼ	"N:̊�A��}G�v�U�]L���H�0��T��	*QiJzڽZϿp���T�]`�(���`�!�w�����
W-��h� Ey��A�*���[/��W�N��`noY��)"�>�-ጱbKQSnAj�|N%��>��������2��`��ȃ�&:#�-V��0�`��X[JL��~%�vZ���J�B�Yc=�\��[���|��9�B�4fbE8S-��hM��f��55w������2׋Ϧn���˛ǜ������B��xټ���H���T����N�Y�P�{Y�N�:�^h���mf�L���6�#��J�pމ����X5&W�jxpQ�ѲI`�M���ʄ]��{�r��)���x�(�9���:����3S�º������$���'�u�c\�����������}� �o/�&�f��߃�3ܴ�5����ש�������<����Ь]�
��܍���]q�Z8 n�A ����f��zw�;f!�U���̧!��1'���n�q�g�� ǚ�5�8� "Fy��T9��slBCeQKЈRyrG���Sc���m�1��:��"�6G�V��chz'� �S��wGΈ�-^jvl!k�ۿ�C�ka�R"B�<�{2u1��q���o�D	�E�/%W�hz2����cy�ܫF?}��!���j�%�ȿ�l�8�h�w:-w�T�
4��������C �Oպ�yS�bLoQ>����;Z1���*K��e#JN�¦���}/�4㬜+��1�T�����&�BX�|���|[�T�;���A)�y���7FRo��RNL��Ռ�}H�\��������0	Z!X������H����L��'�D����.�X>R^'�C"���H�F6vɜjJ?��>�|���b����}H zȌ�ŧ��#��Ѝ_�9l�"�٤6�?�ܒT�ᨁ���ۤ��4�R��\-}{�f�"X�u�8�	S�	�����|
sw�&h����1�t7t&��Yx�8L��Mфf�}��qT��?��j�-�Q�JN�$�6L��;�Kְl[�v�ߪ�KMJx�e�D���A���C �:Ql�$2C�����Z�bh��
+|t� ���N��赋eyLO�3�=���1����Z���N�Y�k�­�(�`%"�L>iN��9�!�G��%g	�CT����N�ӏ��m�9!�m��Zagg���Њ�D��!��P�K��1d�L�����SS6�؞PsnZ/̓���	�}��]�.���*Y��X��:B�ם��A���T�Ä_���7�/��賿�1ݡ<y�X\_.����b��v.�׶+�M`dY��Wx�B�7�#tc�n㬜&�UL;o�s`BM�����wȯB>�Qg34�$�r��)�K���L ����؛�iV�N��l<�ύK3v�ݮ�r���2F�7t��ѿ���?�"�IU�"�w��/�:*�@�$�ߞL'bu���Pˠ`l�Ѕ����̐</�l���\��^�0rԦ�H[߹�>�,������`۰���d�~��n�U�x�8R 1���<w[S���A�|�ξ�6<l{��$�"������W�|�X�5�U�� �U^��4P�U6!��U-���:}j�Ѵ=L{M|,]J�O-�3ܤ~�,��H�a��|_�[�.:Zy��~�Q7q5=n��u۫��Z�9(�ʈv{l�ݠs�G\t.�fZF&d<t/B�8=���9�*�3�qR�=�%w��|y����A%��W��Ybx�Go�vd2z~~e4p1~� �CeqWQnj��'W=^7N������-w(Y��t)r	T�(�m.Џ�L� ����BJ�/���~�0�q� �g}~t/�l�'s�hhe۬�a	oG7�Ԯ�9D`�c��sߵ�f2��- $J�jB��Rv �<���P}�nH#���]��պ�Yv_�yñ(�Ͱ
��!$�H�0���a�����L<�p������%D��4u�׹ե��s�O(�-���bV�4��u#�@N�P԰I����H-��3s�y����_�IH`���:r�9Q�?e@��wmo%�I�?vB���{�	@@ΞG!o�gs�]4��>�9�`�̆V/qa�ݠ��m���GŶ����`&�#�ܶ8e����M(B��u�8k<�}p�S�m�C=�Ƴ�  1g���Z��M��/@h�*�5��tFp�Um�uK�w�	�JN����J�4���o�Bu��2�{ȹ*^U|����ˇ�z��g����^���/̰2��"X��q��M_i�Z���'�l��n�?@ե���Y�8+�;�T\Sv��*�A|��������6�[+��ͻr�N8 v�Q��a�ܢ$bڧ���N�=[́�tWt?��]��4�xk��ޕ~�	��{X7^��i��U��(���m�{�\1**�MqJVYK��~�=��TM�p?�	2���.�:!^�7y��M�Ä'%���H���){B�f|"o&r@N��F�+� �Z�q�F֨��;����?��Þ�s��48�
K�ct���tfR8�Ͷ��x�&!�����z����^q1��?�
���`���3�	�xc�?��}3���ٞ�Q�/��'�g����� e�Jdܡ�y�b|D4 `_�P����V��]{_m!%�r;��N�V�  �;1����Νc�jc�x؋��U	m�0٦�/tV Y)��B�T��� ���_��i�㬿��1F̄�`�S&�^�r�G��J��T9�Z�"�>��Q��y��Hjh�7��Q����u���ٱ
��5}�)	t���H�������iv)`)v7�ڌ��g3ۋӇ���M��*z��~�^՘�c�U��z�G^�M��?��Ϩ�Q��{�Z���±�����|�2�vF1xJ?L�T>��".l�[ą����!�/?)qdQuQG�
���)��Q������q�9�@3�P�����z����{k'<%�Iħ&"��N[��*@m�Gоx�{���W�ɧuo���`�4Y%XHg��"l T�*�cr��6��ˮ6xjБ�m�aF9���%a @f�"c+O������10�����錎mY�����iNm�n�V�����?��;��\��+u�R!�s0o�̃S���v�}8t�2A< -e���.y7ҧ-�f��8ɽ���\��w�,�����9��H\�kA�7���)������wec��=�7�
2H<w|gm;����ыM��r�p�f��Z�:X�J����HO�p�s!�kl���{�����09-WVrX�l6b�����榼xm��B+@a���h]��S{�����b�6��·��~"��L�Jjitk|����=^��Kv�0�	|u��\4�h<|��e/�]�9a���W�{��(@t����u�R��m[#B�0�~���M$"���)�q9��\�溶y���k#��I���A�jc�ne�7i�~}�V��Z�
��!u%���1`��4���99rkȼ�a�9zdZ�F��jÒ�D���S�q��qi�&���I��w�X*���.ْ0"�^��6.�z��F^D6�%B]���i�B�Z���8������L�� ��C@_���VWZ�����+�nS�Xw9@������K�A��! &5� � ��Ƥ�hG�E��
cy������]h�	Lb��.�2�=����p�pY�q�.��.Av"q���u�m꽐X�9<�1]l�Q��!���l�$jn��\7C��+�S�4UD�\oz��ٴ�s�>ܕ��;�d�xn��\������E�x�g�5��z����* �[NYq{2֧���]+T[D<��j���b�;�e�s:�^^�Z:�g��kJܟ�(vϢ(��Sc{ǚ��&�zȰ.�V �}���eI�<��{��9��7Iʋ��dG�k w�X*�0Po*��a&��K���֤σ��M_U�a_:^�h��
IWm���B��������pK�gX�<��I�1i�t˕���<pxP|a��v�wH\`$�D�nt��}�!N0H�P����Ez3|/��wk�L��>%�x����ᨧ���"H�����ZY�tW~�C��ʜ`��W�j�n�|���2�x�[0����2S��Z�b^3y���c��/��`�E�s�zJ��t�С��&*򱶷{���D�{�P<��
y��H��w�<���潯}^�X%tnj����Ž�cR���d0S�m��Z�̵Iz�T�6_��gq����:i���ٸ��d��|�ڀV��!�7�*ݕ��g �ٔ��:�����I�~��3���6�(1��-�X9��.�V�`�!9M	�����Z���� :�&\�8�@��X$sg	C��"��m}��q�:��NK!E4��	�p��],�DZ���F�OoV�Pq�C��"/��tlPP�Y[с�����<LM���&-$p�oLo�2YT�gqw�y4>�������Ir��|����g���n@hԝJt������}�<GX�����z.���A����S�ܫTL�{˷�13�خ��sb�#���4�#�7���ߛY�p|	}�˱��� �*$�W^h�h��q��J�6���f�/r�H/Ǳ�b޹[�����#r!]�KXc�}TU��Q��(Hu�������zJg	�N,�4�\��B7s?��"�| "M��A�)���V �{�R��XPǑۻ��Q~%�V�u�{�&���L��Ɋ�;���:��@�R r*S����ik B|ë�+0�,���t�����ePЏ\��5�r���?�~�:<N��'I�߰��OL�&^EH�J�`Jq9�� ՠ�LA*X �d�Tg��BM���m'#�$�T'w��ǝǓ���BY��P���B���/yub��XX9-�K�V7ѵ��&�ܒܸ��sG����S9�Sø3w.8JW�*P�C�� d�rk�r�RJ������Dce������#.�I�EPw�x���mHD����K��Cॡ�^�U霗��Ș��v+q~j�x����mE	-y%0�����~Ќ{r�L��~�7	>h����F=�3=e�ZkD�{�z@�|�(1Ӈ/3�u�)���sđBY��eJ��z��K�{�,wݖ�R6od��_�����u��[�2Y�nw:խ���8n��ǟ�f�>O�ݖq~UF�B���&L%I�~=��aA���Ơ�X���Q7�X\�}m�@��n�Ⱦ�O�Z?9����� ���]�,m��U�x_~�����X\^<�݊BA��c.�ͪ��;����&�\@�]9�.VjT��0r���uD�y�h�19S��������	6��r]�M���
q��#�p�j~yY&6���cx������/
7�y�=�/R$O��4Z�0o>sn�v��F���sJo���;�_E`�+�A1�}��-!�q�V��6DI�W��nH�Sd�܁�#��/U����(�J�Z���*8�:Se7�Yx�xj��O����X�ٳ���oіB�k=?r����w��K�U\�8��
��'��1	y 0�H(�S{�l�'j�o��/���hP"O�Fb����l�Ԫׅ\�M����Ƭۙ��e�$,��Pf��~���5�H<#-g����`q�i=�<m�Ja�	=B\���$lf�e�A 7�|������p;$V����>Q*/��N(P���_m�.U�:�F����$g���L-љ��"�w�������u�47�,�d�&����imɫy�����	8�;����d��[�zPlii��e�<A��qfu�w �FWo���χ<;�f�Q!�n-��-]z�od7�Oۤ(+ʆ6E�3����h�a!P����\e��F�Ɛ{�L�y���JM�%�1���Q[�[2ւC��<$�j17t�Ic �Ayo-�5:�[�_E6o�����_��y��n�)�VGY���q[8����NZ�3ܭ��,d�J�e#- P��O�-�AI�Z��m䑾�va��y)�SF g�27�J����u����H�Y�Y$5�˛a��
�s��k�oj�IU�E���N�T���K������`;�>��*bL.�4c�B|�]������f���Z$A.�~W�BF`�a�0��iת\��#ǚ����u�e�oxBS��-�ǝn��5�Ud�W:N�]�&Ё���i~fD�j��Oܿ>N=��M ��@Ҵ0�Oʛf�M�&��($ե���9(��\���g�6�����!%ؖI�ƹ��}�ϥ���d+�i��ȨU�Ez����{�?�ıXQ�Nj�{l'��@�tt�(d��UF�87.�§���9"[ʬn'ݭ����t�J�BFT^{kѧ�����I9��a`��.WwKQi�~�)臟����l=|<����ٟ�-l���m�̹�|����ZٺL��BV�y�(�O_�B�+��$�����P�A�c����I6�s� ���[��u���zu�
�j�e����e��=��8�"l��	i_�w�?��P�Z֘"�Η�S��6oYW��O��u��0�E����<r;�j"0e;�h�ky[��Z��,�] FgGS�Ufal��7@��e�>w�+p�_^/�����כ��*�@H�x6~X��f�A���~	�`j�r�<*����_�~9`�J�@L46�&Z���<��..�b��1�;N饫aE�D�S�/L�I����`�Υ�&5�Ԗ"=k�U��ī%�*���rh�������P۾��>̮;��@IYU��+��l�KV��$�t"~S��r��"�x�_�l��O��mP;������z�T���,�Sn��؂`��aN�H��h�1�V;F��n=��,���"��p4���-�E�醙a>�-�f�6�e��1��L��I�<�wc�`�Qr�N�pa����bt���#�/�>�����[�6C@s_g e&4�ǳM����1���f�6�i���標
�C97W�6gR5��w��	]�T�w���$,`��RxO�~�|q&��3d@�#�-���fqJM0i���s�V2��p;�,�U��H1#\7� �4�� �vLP�Y�d�s�n�1aRv�lk��֛zQ['�8� }S�Sȃ��c~֔��?�7�}�䯸�T���eB㰪-{�ifg$��$# �ji,�܏p4(�'>���a��3�r@�H�b�R2b���-�A{*�2�w��?��EŮ�sl����2E/R'r"0�����q�-��ɥ,�0{����X%�j�d)w��G5�H��21�Ѵ��*����OkWBܒ�A�.W(Ҁ;��h)���,���''硿�eP8b�t�3'#��Ͱ��X�.�	^#���~�fMZ�����<����~�N����s+cO-y��
��k�;�zӷ�=�X����m|��Z��N�_�"�%�n�ֈb���,a�n�Իo�O�^�E��EӀ&t�^�Yl|��$���
�(���g��F�#e���!y�"9K9�`At�+a<�R������~;�A]c�Ae����]�;�(��<sы�D���t��m�myY:���e���`�3<ڨ �0_HCt}��)�T�lE�K�FmBli�
��>ޤ�?�+�AI~�����62�>W�4��H��P��8�e�߯VE���잦ش��>��!r�3�HƄ�aC`����f�����D��d�.!��ʗR��ȳ	t2�W���vբ0Av9|��wLAɤ&��%יl��_&o���Jw���D_��(,�z��ҭ���α���B9L8�66���L�Ѻԏ��$���W���h��AN趷�X/����U�OAj�YX�۵�~T�_a���DQ�Yt�k���#gC�:�:���U6�ǫ�aS^ξ�C�; �b3�#iF�"����<�gf&�3�W�H�Oqw���.@���(�����%rI���"E�|ݕ?��tx��f����N�=8���Nv���E6;�Ul*��l�V���R��-��S�>d�v��!`@�Q`{�͢��Y��F!� f�D���Q�jo�K���^6��rL�z��1������z+�vt���	�Z���ě�81�
2�N&���]�tЋ�@a�9v?�Hm�HGd�%���M\\�zs�]�n)���_|r����'Ⱦ�`���h8s���Bav�-w`�`$�լ�z�v��dͽ��Ij��[[J���=
#I:t��d��k��8]�<x��Pe���x�H��OS�@���{v()�M�X��+��Vn��
8�5�n[�2c�zz��"����Q�+Ne�E�)D�h�H�5��N��v�b\y\&���8�j�Y\G�2ګ��Ui���\�ٖ0j���������AS	*e�M��D10��<XZR��F�`Z3�&�<
n�)̠�X�a$�R��G��M-�o���+�u�(���ކ3�R��A�@��%c�cX�P�+0��!Wۼ�����AVS�k����J�g	�KA�P-D�!|x/�����?Uy�_�@/�':�H��?v�S]���  ;��JQN��2Z�>}����n	��u��.~<�YBȈ2�&��
�wq�&4�5�=3ٸ�X�?1��gu8��^��H?��Ȥ�p���F�2$��[���}�܂��;*p֭����YD��9V�܂��<!��͙��t�Q\�� W�$&[}�l���<
.Ph���oM{�a�_j[��ffǬS��M~p|��tM�t����
��,��v�����_S�M�R��uؿ�/�{Ȓ���>qh�j�i�6���"V^�tD����tr6`�n�`[�.��Wh-�M�!�~�݉j�w����K��g��z�F8�No?s��e��}2h������I(�-��/͝�}X��ݡ�z����0��7l�=��D[��<����sNb��p�]�ϕ�i�־bq�z1r��Sا�j��Q����Y�� ��-) ��b8��M׹�D�A��
;L�r�ly[*��J��R��o\=��K^�NH{.�.I�WQo���pH�ۓݰ1��}�DW^�G����D���%T������1�N]�x�w�Ň}AVW�f����Ҧ�kRx���Llh�u�@'gw�\��l���r5���E����V$��cQ0m�HgN�y��4��Z��3���`�����+����$^[��Z�{�_��5��8�������ag�������7�oS���Ѹ�f�Կ�S��q�NK;�m�oY�z����wq��SN$&�HƎ` ø��`{" MӮ\�[$5Kρ'|Г�,�ӝRF*?�o�"q	!���Wp�E*�{�pX=pQ�eWNo�}O���<��"rjj��yS�w	]�`}�����ެ�����|�Â��>��	��hܝ��t��F�'6�x\�����`�f��)����W��`y��)<[W�db�?h8���B=!���S�$��fq���` ���hz�.X�K�6�V��'�B3n��nIm�-�fF�{��w��������?� 	ⅷ��7�q��	%��_X�U�`�A��J���fyz5o�@ p���2*�� +�ЄL���}U=��0���,��lK�����њS����ڛC�L�)|Q�� �7e���x ��A�`UЉV�#Xt���<��I�S��ί�N{���to��GcF��/ˤk�T��n��̮2�@�ة"k=��( kְL�J�~�HE>k�"ܬ�����RjE9�w"1$1�bc�v0]��v�嬮1'�E�osi4����T�n�� �VN�V�	1�+��6�.
cJY؈?5����Ǜ�/�=�6U�z>�[7>�x�4�
h�N�����蠞��oÌ��iBz�b&h����)��i�����mdr��TԴ�e��F �]��O����9���I�^x�j����'Z�q��;���2�b�+�]��B|��f��P6�%�WXHB�i��5JK�ںE^w8
�r�w������J�K��$�\�򤈲-`�>[I��?�R����@֖2��Ġzb��ڼ��-^�qN'wOG�|�=z}öN��ʚm�S��<:��"C4k�j�x������+Ô�W(�<m�*�}�|VǤ���������Lb,of�����_r�3���^�1��c�������I��@$؏��qfb���$�$������H�u�#�U��/�X�%��=>U�R�z�S3f$)�_�颢��������qFpg5�a1O��8��k��$����>A�a3����^� �q���w$a�n�\�Z�L����Q������a��2Q�~�罱AR��C��1�<3vP�|�G%m3�x�k$]�"�i���U��Ͽ���sAF���qұ7$	2B�i�̡@E�mcE��t+�."W;%b��HʞKe.._,����\��u-���l8��p��a������uK
�1Iv��@�aU7�8��9V&��̽��̀!���DeOU�v#]č9�i���MOa3b��L����9<Q�lqv6RӅ?鿉/
�${�pJ9	�=�b����'����f�5ylT��5d���X}��Bl�X�f������R�c5���� c��=��TC#��h��SS�k��֡5�*����Wu�}�;T���,ȸ�'��U��(_S���u�����p8�|ŷGS�t�ż��ay���"��fpN�T|�(�'�)�����.���A�'��K���i\��d�1��Of���?L^���Y#�j�v��GZ_E��z,kt�9=>��@"�[�UY��R������Rn����i)��Y9^��j)q���s�A����Q��"�e��{T0�v�����u�P�l��z�f�\�km�\�OQ���뿰#�����w�ڶ�zWn��[z���`�#�~V���5J�C ������o /�鈄c����T�e�ը4p��>����&�bQ�������E�P^�Y�s�ߵ�� C�L���J�5ch���܌�%N&"���/���KA�'��˭@m���D٧���Q/(���������̀��Dp1�@2qne(}���F�|y�Qn�8�g�'�¿�jR��aBSw9���Q�(�G4���"���M���P���~΋���]'�ydh^�����;�ܽ���N�����]UM�e�ׁ�ځ�$mgO�q������\4��VP�Q�Mqwd�+� g�z�ƭL�C+m�+z���r�=�U�*_ft�$��v��NL����/��5�%��Lɳ+�R� %�r�[+,ݶ��Y�~���ֈLE�| �$	���4}��V@��m�IӟXϗ�o�Z	�z�sdB�:�iޣ��g���?��J$q�����YШ�E�0u�h�9mA��I����t���-rRa�z�*��ˠ���Ӌ¢б��M�gf7�DC�#� 2��:���o�xTHR�ܣ}[���^�L�����x��
�"�ϧ���/����貱e�,��*<(�~I�ZҒ�-�O����.g�h7���R3��'eRrd����~�����n�04䟞��fp(&��H#�ф c�)� M��S#3bg�� >����5�	E��w���7條{:�U�׆����"�wo*�p���Ë��JoYX��1r�l�"D[xު�O��Ŧi�L�¬�"�)V7�ش:�G��kXq8݀�|˖?�$���BH�bb����4>EBu��YQ���Pl?
��Y� r��	�r�m���!g��Ypu*=x)*��y-�����2����|��k������'�Wz��.R&pj؊���:	Ylc{�,�ȤQC�哏�aLn)�{�uo�?���:�"4A��fű[��U8�]�����༰�蕮$	,���E���t;��i֤���ӿ6W7��VSLD����烿0W�[�����$յt�����&eL�N�:�g�����ea7�R�/��g�1Asj�$#�;��&V��=9�hT^�!�WـtI6=.�G��L�ק������X��d�>��o<�Eh��C Ҳ���Ĩg,��e2�f_��)�9xeD�R��@y���-u�)	�[m��	n��I��F���m��%�qt���yf��!�ȱ��vg�M�f���;��8Y�xV��4[_�f��l�b��ߺ}�x�jF䔑.��`�?�L�������r�͇I��ק�@��\�o��O
|\��ɳ��lx�S|T�[s�����+�la$
�����2Oe��?�{�������}w�^���SN������PX�q G��kh=��BVP��pkiRoߏ����ɛF��>-�;��gN�I�.<:�Vs��E�yQ�6T����硜P�`U�̠L/q�P`��Z�^?���z(fb�����Y�������
�ر-䆚�MgG�>�m,��Wi� �j
��r���~Σ;̦��3�@�ե[�]*9�8�KU�i-��A`�Lb9J��kZL1�m}�e�kݦ��غ׺&T��Π�T8ոζ`@���<�ٴ|�i#)o�%6�h��TO�ϜU�!����e#�\�ܮ���/!IOd7C2Rs:�O�OR�l�%���S�$B{EU��Xy�՗��n���-�O�� �v;��'�.����8h��ݛ��jUnl������?mt�G�݇�%⺄�\��.Q<�& QF|��:)�ꩆ�¨H�ՙ�Azs�g�	�.�� c�����ED~ߜ�L�Y�ގ^y�u������uc.ix�f�D��-x�"r�,�{��s�a:Q���S���7�:ֵ��� �*F��uP� �
ۖ4S���\�r������;���]�f���<�����\�s�����s�B;Q���n���,La�_vd3��rP�
��h�בrb�(��
Gr{���խ�x��zy�[�w	H������Ŭ��U=g �4��w���t�P�x{�V҇�4��;��?��*� �������6p1��$׀@������g9�D����y��eJ�8��`��;��llZ���0'/��͙i��n>��o��ϺRF���Ќ�T!�jR8��I���50 @�ѝ�cv0Ně��l��kM�ؐ-�	2��~�H�t�;������-��wЈ�FF߽y�˜�k�L�
�}v(�W9��(G��*I��3��$��K�l��K��AijA���m9��� �]�ù�h~>�r��+�)&R��M�-�pa��
{��3��=���VP'rl��B���33b8n�6�IIM�"�?�V\NU�*�����*��4���,���oE���a�~�����	�T6�e����>S�Q��!���ަԶ
���)�H���h^e�^�7r(������w��4w���&��d��a{�a�����D�2��F_�U�uzJj�(�h��I��oxYw��i+ G-DZ@�@t_Ik���r�rEp���h|�!����R	����`�4ϫƺ��zʞ~�ӿ�Td�j�l(� ��`����+�1<�Ͳ�F��$,\�Dܿ?����F4����&=��!��6����%C�0KHǲV%1�al���^���Y]��̗y�����H����X4�q�J��5��e|Z["��IYk�YPv,�)ꥦq쉵�f�t��h\vx���U]8+0n�\�܈�3�Prx���ĕ
s�	�.?��D->=�9r[CֳSr���%�S�b3��kD�
k�[O�<I*�O;�s�N����d�����:�+�y��UZn��A"b���wF]��P��~��!���,�Cʪ�~9!�`�c�0	w�l*h��7s�yӸ��/����
4h֜#�<�����@^�1w�[�O�I��R�iYG���~�"�+k���Bcdj�"Um�z�HIC�S\����8E���+��R�z}���XAW����� �>�;2�_��~����3������dPl���Md�LE������^k��tl��&��>&�)W�����*j�*�U/m�F#�U�5ǘs����J����{�Ɣ	�R;�gIY.�w)
��J�^X;�yS��MÔ�6O.��Vv���0U�"{%�ށ�#"�Ư�d7�8����yݜ���Kc��s�x��:���;V�E8��	T~��j����HO#p#$������fqNT�Uu�i?�.;`i{k�5�}C�d�s/*�-����������v�K�-�:�	+&ŮT<r=Q�x����Ň2f������e�z�45�lO_�\�;�w&��	�%���U	u��F�_��iXy�C�-�`8XF���Af�bIs��QX՚h��o���}�����Z��?��	��磾�Tf)�m/>�x��e�ߞGD^�����.�60`��ׇ=d"��Q#�"ޅ�C�9_��5� n$��R�t9�+�z���o��
�b���T�[��7�o����H��0"�W�Y/:�_���[�������AH�TΒ�g��^�����4eO]X�i�S�����2�K��Q�����EzhK�2�V��R6+��ޯ )?��ex��d�o�|C��@y	����b��@�{���i��wبUcS�r�.�Մ���FbX��E�e��"�K��!>����UûҪn)4u�?�	hz�,ì��.���������F��ʂk��+������Y�����}�hw\����&�l6E���.AY�Hƒ�#+X���0q~n��wc�&0�%�{�պn7����P��.��kr����p���8�e�d� �1 �r*��Ncu�B�����������/�� ����֜=֮Ț Q�Z�*�f_$g�Ή� W�\?8�����}1��fE�$h A�d��~��ǔN�8���8��n���0U��5�}�z��@@muew+YL�S��8�cAV�kڻ'�|��hH��9{���������[!\�@�+l���{�����o/Rq�x)�q&8�4��Kr܅��wB�U:�w�����s�4�j�H�z�N[���U��?k�Fb�9�yi�nB��<��l���(�@�da�l�v�`�&W2ta>�%2��s:X��3 �Yn�B���?�����,��t�e�]a:�hIB״��+W�*�"U�v�*�0���9���).��-���򶈮-�;��uP����E�{��p�md��l�ŧ�'�)��O[�[;��1����7��uR5�!c�
�<n�q>��2
׊c��O����_V�4	�4�L���l��&�\W2�����52��C�ܦ���q33�1�b+���-�F��T@nx>�6���h�a�?�qY�2b7�C@)���%D��q��������@�A��?�g�bz��+�)p�7F�-�ާ ���K-�>��/V�\�Y�=K��YS��e.)���dam���ƕm����y �؞��I���6`������N�Wr��!�����rM�T���d^�cJv(}�����<��Ԥ/���#��HxD�#nwh}�ERx�!�A��!�A�G���V�C���x�$��&����kϴy�E�j��O)�(@�hR����:�K���Y����e�2���Q���V��M�|��U���Յ��6F)~�B��K��)*��1���Q��Y~FZ��t�m�������ar�:��\6?נ��I�4�5ذ�x	\�c!/'e��)w�߲
�d�s|��ԋG��!��½F�Mp���sv�p�y>Hz��w��o� �Ώ��Mv(XoZB�f��*H��8����7E�뱈�3����;���WJx���Dna�w�ڢ���R�/y��-�%ǳTU��[Oi.���a+��߮�,f5w�ߊ�id�W'{���(:T��S�����ʳ���u<�q�5�n�)�aeqf�<��t�u�&��x}�R�e%�Nc�L]��ؠ�&�ӏs���_I}������f�4��`�ZV��A�`�;�a�����Y)U���8�}�Y��>wp/ ��>L(�Q�4G�C�z^%�o@�@���4Z�>#>��c�����>�XVR@0`|W�x���uyhu��1���G& �d����F:&�#�Tx�S���(X����P�<�xJ�xb{O�ҏ��+h�_;_h�_A����,gdV��>HD=�K���Z9����]���z��D3�*�x����s#,���<k�r��%�3ֿ��,����X+� _f��]NC���yrU69*�bv,�����;]�v@��3�G� _�!$jɫ�J�TT�|�!�hd�tT��N,kv�&���;<g��A#�i4<�qM//>"P͈�����`�����(`��ڷ=^#����B�b8��f�bL&�0�T���+̠'�֖�
�o[�#0�'�qvr]�b�02ACq3���R�6-�x�)���$��J�����/ 8�r05izΞ���U�)��&Lg:`��#[lu�ƞ�s&�r1 �_ٕ����������7`��_�2��ӀB����Y�I�=��V�V������L/����Ӆ@����n�b�����n��bj8M���l�}�s�$�[x ��jS��l�pU��w��ٔWLhV������,P�ӥ)���� ��8���w�b�p�OT:�����X,p����ō�6��5��4����9����"�C�ۣ��PD۔�L3�aY\�ቨ���u~=b�6ж#R�?
L��?�;�G��ov��p�a���)���p	$'��;m�+D�9Ǖ��@�K�d�8�qs�#0�[�^W�y*%z�У�7Jf�.#�>
��-D�?�H(��q�>&^l���1U�A�R���B{0F�&�[qQS���B�օXf�OMID�0�7YP��g��viG)	Ҩˮ�aSx���[$ν�!��6=�=h�{��Nl���ן�fHdDK�}t4ْ�'@jŨz�^fKz��Jf�r�����J�}KKd Oh�/b�=����\�FzW-�w5#S�\<F�t�,��+�͍���Z�d;;m ��U<
ev9�iz9A�梮>S���x�e]�N�kZ�^�7�x��IX7:ؓr+�[G3IJ�dx�/��s��z�{��+L�A>�ڿy2���%��uzs"A�B����ːH�>5�fC�Jtiȭ��6�I�ZEr�wV��unϦ��x���QWM��N�=F��\��dSB�m�k�ا�2�Ol/�� pW/~lG[�}�#����F��!����0��������|��7s(���-��Ae�=t	i�C����${f��^�o����cX�]w	�K���3�&��VJ�^uQ	_�u�ّx��ٟ���k�K�&��t
kB���K���At׿v����@�@+��_���ɴ����L�.�԰��j���.�ELl�\�ܝ)mZ��SwT�`�D�ޢN.f:��鹑�e�%ޚp��dJ����}4\Q�"��#s
#|�oϱ��O��p�ю�L,V;;��?8���'9&���x����b[���~Di;��#��]񰤑�ԩK?�m����'~ט�������Q$NU�x��e(^-�v�����л�8xi�q�zƥ�Ъb ��J�\i>�15�//bM;�ɒ�q�6�|�ׯ����yY����<⎠�α��Do�V����c���%1�jWn���,�8�5�	�`���ȢZD���)LR���
f�y�jK��o]���0�]�MX��&�'R,��%�Q4��Q��WK��/N��~x�OD��V�_.�1λ���C�~v��?��gN��b��̂�(L���ƛ����V���=+̠�>؝��K�}U��6�U����e��*�ĝD~��{ՠ��s��Ig�8�'��=t&*U��fH���O��Ի�-<���HB}b��|�p���"��%9��X�\�=w�r �rm�o�կH7��,I����ɓs��f���&1���]��Y�=F��D�ם-�[\�.��%{^�K�5�8����z�r�m=�� �ף�0���"�޺���DE5��u���q��	�o5�����,�N�)�١��ق$P��2b%V���i"���������lE���A W��[ڵ���������w\�x� y����\��I���a0M&<v��hbw��@z!]�d G�Mq6h��|�q��f�Z�,Q���]��Y�2�|9h���[|w��
%Ac��d���%:�˥�o/�1Q4V�p��Gf��Ȯi��� �ue� !�30�"��W,�S���aKQ (�ƕ���6����Aޝ	�g��(س�
*�����o=���`�Gn[����]���׎�r0r/��tm��y�P���/T!�ǀ-JXȕ,������(��C؁�g��c� 1˶#�o#�$�ɪ���{G�ܜʢ�gf�;�.KR�m��p���T3�f;�.���ck���7�R%Հ��Yy�"��r9�1��������)�
�n���I.)���^R7�7�����i))A��2=��,R8A���ðX�L�&z���K(��Tw��T��R��*���8���R�<W��&9�%������H��~L�2�%Wr�9��1�j��#���J�0n��� �>0��\��d8 I+]B�s��T�J|
�,[�We�TZ��
��F<���n� O4/�W�`������P���Ry _�_�T
k4d�K,\�pj���b�Z�K�C֫q4��$�X����3��}53T�&J�c#ǟ$X���V�����#��ac}�/���Nu?k�8�H�ál̡����0�ԯ�S��CE|UP>E��Q����a� nb��~M��`{/}m��ڛ�у�h�U<S#�"�+A���d���:�5e��v}��0uZ R
���\��1Uj�3�����T�.;�Et�	s,��\IfEKY�(Ip�[A��ca���s��6*m��yeV~q�
�����C�9o/M?L���Q���ej�w"gWb������D*��|3�U�dl:z���
�7���(�U���d���s`�`��ZN����d^�{8�u��_an�������j/��miOc�:�8\��!{<F����O�d��+0u�O���UѬ�<���&h�<�Ϧ�-ֽ���O���2njT�v�/
 �����Y��,ȫ�|��m
.�s3.p��#nE�zw����2�b�����l�ۂX���]�:p��xnhY�^�g^��4&c´���!�T����{k�(�V%\!��$2��7��H֜0�j�����K�>���GDM��'���C��q����x���D0->����6��O��i߻��6���"ٯ!������*7�Ǆ�`�-ϗC�q�<����"i�0���T*�m��=s�H����$����b_X�ܠC!�/O×"�~+�R��*ȗ|�>�G���܋�g���5�U0vѤMz�6��s��BlRY����0�х������o��Y�,tSLX}��j���rյ`�3�kO�3�
�R-h�뵝^��.�*��4���c�hT�N�v���������q��b�u��`�)S�_�?�GP��(�L����W���kP���������9�=���c�Ј(���Bn�1������ރ���s�㵴V�D-�GԾhK���3@%�N=P�Z�R�����L
�Q�H��a�j�E�R����f����;�<��R�a��5{�-�ƶ��q���N�ɋ��ū����Ƞ�xD��X� �1bv�{ߞ�w�D��F]���Q�U-�?y�`��,�KA�������R�=�f��,�m(��6�@���I;t�c&����5k�I��7{����{1r�}�*��G�ْ���nB��������$��"�6DU>�C���b���՚����pnK���o�NԈ�����F�R:Zs`WyJa
nFVN��#5�y�q��6�Q�a>5��8)��5�j�F=��jVY�j��
�|��X�|9s����������1�VR�j۩�'��W�!�̀�[�L?&i�9[�$�0?���N��, J�� �[��a���`�4_�WQ��Z���U���F��:f��[���o0,�ԗ�l04ֿ?y����Fog���屄�:�G�����`a|����w-E��0e������c�v�U��q�# (��
c�08�v16���"���F3��!����ܙ��*�4��cI� ~v�c̠9�"*t)X��b�Q��A��?wk���y�q�¬���#ߧ3�i�J�[�u��	I�(�9t��Ɛ}�y�cq�5��tT�(�Dc|؁ZV���;��&����[1�a	�U�{���W�NC��R�j�*A˩�iI؏�H�m��_�[Jg�E�3h|�Bǧzw��F����}��:هci�!0��7�a�	1�l�Դ�ʛ�T�!g���v��a?�_}��/UɁ �����? ~_��P�y���rpf}�+���� _w�� ���Q3Bd�n�?�
'eh7������ܖU`&���3|N&�g�rt1��rb��$��}��o�_��0�~��x�tiq�;�"���Vw�ICD�F5Lc�3}W !����.���P��\ع��4�����)ΨL�9O��&��������:���j9t��j�)�v�0�bk4���p���J�+Z��U��C�b�jj�G��3U։��.���6�Ȣ�ED���LJ�(�����`� �]Tc,��{-��,q|����r4�${��2E��e<L1�;�y>^9��%(L�:��\5��C��<�\d����[�n�	��^�U�87Gi�l67ѐ*�fX���\�@�J��D���3�6o��CԿg��h*u뷞sӯ5 ��WD�f ~^<�bL�{��-G*���&$�^�����:~ك&Z���7|�O �/c��rj��������P���w�e�~���"����+��`+-U���b���o ��.��9CÿH����u� �lI-�*"������daS-���P��)\dB�����G�(��oM�qt��T<a���XH� w��O!�Ef�\���`��d��;/�=�"mv}T.�~l�ocyk��({Q�Ȑ�>%Œ3����Լ���������:�����`[";>�J��ƨ�tQ��k���)�X>|2��#u_%^���z���ʡ:���ǉ@Ђi�? ��nP��S��SY��uY����<�_+��c��ASA�`8H��՛wziL7
B��n�w�+��
&ǸV�8��ZpgVo�mɄDo2ࠪW
8Ty0n�����?Ĵ�V����=ױMu��>������D&8 �j��$l��(��$ƙ�c BG2�?M��'͎@���S������+�g%�lF��]�-�5�4灸S�iA��PqxTo�c�@�4sK��,]�R$ec�U���x�x�7��ҿ�cqp�5RO��'�~�E&�a��u����Zk��u�{� J��J��+�{�PV��W8�o cKTB0����2N|.A	4�jR�]D�Q<�o�"~�������<]c�ߎ ntPN3���L��Eʹ�o:j��j��yɥf)���Z�:�T��h�{����P�^�M�#3�w� �(�}�l&��m�y?����� 9j-S0|�?�N�	9�π�j5\*4��v#a��a+���m���a�D����v'�\r�c짋L��8c�%̜e�	A��	���m�p>g'��D���07�*��T�<�4�e���8 o�7pSmyD�tr�['�]".?/�^q�n㴎�q6�IC����y��)��	�I,T�G��ۊ����	4=yP�&���fX����W��ʗ�}�����ϟu��>��D�d�SG,�+���۸������?��*I1��%Q=��2&z*l$Qۻ���O���}��U��2r��$T�>� ���S:������65��:S��N����*��y�煄Tռ1��ͯ-̫D�߆PI�l��R*μ�[8t�Qc
�ӛ�x��H勋��������-�A�MC�����JZ�r�v��+�㶇�r	b�H��e|�L��7��hs���<���8:h�?w���<T�_H�B�^���K##��f�X.�"�����=�M�-1a� �KB�S#��4I�P�8���Jд��9��%Jy1�W�esf�N}�<�1N���_%�Wp�[���ڵ���Bد%f��Dұ�1�9�bRI��'N}7?��fŢ���U8����O��,�1��ћ���$M1�m�F����� o�j���YS���Oѻ#մ��E��*���Bt6Gm:��w {iI���
�`~-<@��+FLۈ/�Nb�2����R�u����)?��Xվ��D� ����^����!2(�\K���?w�����9�+�ҵ��
ފ�<t�C���ХH�-m�vO��2�V�2��:^;���]3N\�h�~�*�J䱔�5d"��~�֧�_�{<�9$޷���
� wZ�U���+���0dɸ��p���F�P��\�~�ײ(<���JA�adÛ�V���.��Kj���q���L�_]��B��Щ������� ��o�_O�`��/���4�@�Z@���:�ͫ�</�v*[A�d
�>��.�;��2�.�KyL�Q���m����S�.c��JEXI�ώlB�����h=x��E���*�F���d�|�m)W�y��3�Z���+b~p��D	4�lpԦu� a��yE�8J{�9����@;Ba��H��B���B��>�7sw�!��E�^!Ö�6t���|h(\jM������^��̾@!��c���M?�ٹNs�2��?��X����+{;Ā}Ik�15�|�r+���p	�mí��5T�jn�U�����$�+Q6�w���($v��6fN��87o�/Q�^B3+����mt�-�Pሩ�]�F�[~���wO���.;�m�b� ����<�_�	xə��Č��$L�'�n�4�Iʣw�c1��=�Q�u�����A�;Gk'���;�-�w1�-��T�[�-��g�}��֣B���!�L���˭s���UC9����v�ѻ�Tt��+ ��"���k�x��@���zq��+�sd?��]�j��V�Z\*��&�,��EF�Q�oK}O��B���o�!���{��'�V�cS������ K�ޒf�۴�F9�e�0�rD��|���A��o��/NׅCu^3�le|�I�U3vޭ^��sҧ��P�+�\еm�	�Txn����D�J��*��������KNyH��3r����o,�'���9�nl���}���yY�bI#Ń.�2�=��I��@ypն���bvg���C���1l�o��nc�4�9̵�Z�a��_a,�f5��ZkȔi���vND�-C���w
)t:O\z��.�既9��#l.��MA�p.Áp�`?�Z����撦nT�xZ�ny*��ʍ�՜�$�D�UX���1�^/�%������j��8�&tK�`�-M;�1�'V��+����A-4$JjY��>�c	 ߷k�j̸4�ώ[\o<6Ä?J^T�b��kҸ4!v��T��X�v��;t�o�{��
E懰:�k���I�Mͨ-7Պ���Q��4�;�4K��g�.�"�F��0�6��NV>�Yɰf�o���a�f&0�sa������~���n)�WQ��+>wf��l���dzYFa�� �dd�t�P �����a��mv!xMl��������L�(��!�� P}�ٗ>S(�d�ҧ�k��9��T�t0	�1�Y�Z�Pjy��ݘK�g��D��QY"��O��"�c���z/��� ��&��@��@���Ʀ��Z�"9Yƣ �$�	�E����G+
��j�G���0�������v��m�݉R�7����5]�A����dG�������":��Y}�"�������^mW%���}CAw�� b�_����R4K��э���qDx�lU?��e������%��Uv���8w��j�������xwDH����^$#�e#�CB�J��;�BҸ�K3]�t�Ʊd�[��� �T-�W�R�^1�FN�	�i`����v/sR�dc�?T�A�=�t�<�3VzRh���7	0��x=�j��Q���j.�L�}���d��-����NI���5zU+F���2�t��g���	�B�&-8r�\׆���2|篓�����w��
4Y�+��'w컄�
�Q3�=�xx��M7�Ğy$�w�g�e�4"�T�
�x�y�`���ϼ��L�y���{�m	0�>��Y� I��y�E�b�R|B�D�u
��woP�
�S�K�<�e�]^�� �5�T��o �	/Xi�|,��56G��Z-S���T@{K���D#928�)��{I���{n�ǔj�i]�Ms���r��[y�`��4�N1�腰w��_W�/b�Ǡ�����g���C�c�Za�_f���&F��r���J�U�\j��?��k3j��PyI�RJ��)u����;��ފ��gAbw}c���~(wZ��V�����:YSx�B��\���L�wI-*s].G oj�LV
A�3�%��B�B����C��2���f갘��<q�V�"���0 Z��r��w�tm�/ɼ9w!?��+�l÷/��p�Z�Ȳ@�Ί?^ "M��]Kz��,������mb#s���ם�Զ�V1`I�`�/�G�aB;.��P��6�<@�>�!2g�V����o|:��P�R�;�P�:�c�4���tŷaL�(m�������"�T�GBO�g�,PFXE�G1!�ݿޠf^���ъ#��%�黤��}K�%�8Ǫ>	����������9i����M�-�F��7$�����#u�}��V!zl�����C�Q��8Rq�(.�;w��K$5	��зPq�c`���)ZO*72��!X�_���@P8�I
`��Wu�s̟���zHЧk^��X�zL+�'�R,� �@�Ly�x"tr��Wˬ�\��u`�A`G��u��{D�>�f�R�8��HضS���nB`�OL�0R��T
9d�.?�Oe��K��l�1��[�sW�hv�z�`�-�h�%��Bq�;b������kmg��.  .�\'���R7W
,���s\<#z��"m�j�jX��	227�e����<`w� n �f�FM(�M{��5��Ւha��u'%?4Rɒ�C3ftv�~9�у���	��^Vȏe� ��W4��$�M�Z0צYm��W���6�H��sϑ�@��1þN��T}O�Ѷ�Pmv���/r[��s�����O�5h]!�}�
F����/aڡ$"��X�}��T� RbZ�:���8i��D�7d_,ǡN�(�V�gh,�^a��Q�ļCr	Q�̟��b�������-�ET0��F�����m�5���4m����5�{������R�
�^5󕲌A�m S'�������μ�5 PEe[N}b�s�6ɠ��H�4��y6~��!gf�"�a��s���ә~��nG�&��e���?V��I�<*$��rb�!�g�W��~��C1CGXm��kD"�]�5d���/�[���E��oC�"���p�s���J��׆d�����@7�כ����#���Z���s�h��M\��;��aK
����>u��	�7���D~R��?�ӱ�8��5q���H
�S���o�� ��c�A���RYO&YV'�M�S =v[���Ӥ4'#�Bsq^[A~D�ˎh�9P	2kkV�}�?$�8��>T��6������ګ��`Tv�~�m}8���1ý�uMm�_Z�ͱ�S��B�8��U0�i*l�8�z�X��ϸ�#��T�͞���=��D��&��۴�������!��.F��+�:qr,���[�!����A�x�~D��qb�7�݂�=�}�Z^\�O�:p�61�"���Ǻ�P��T݅" g��|�	&�n� �S����0~��X�����顐���7i��l�]C1g	B�H\�L�?,�m�}	�#�S��-�J��+��`�~�UOt��"ޱa�p9]˄c��r"K�(F�Q��~�\i�3��;��l�D�R6�7%��=���36������t@�P%��%F�s8�I����la6�+����`UYyT-�R�j�jPnغ������V�S��ˬB"y����%�ò��� ��eP�,:Fxw�P7�i[&3Ū���Yu�OC�7���2���1a_�y@=�Q�+��A���e���4�(O���4�D�$	�<��X������(��ޯ;��C�%1&��Tz&�iz��߄��soa`̓�,"~��N�+�pw0Ѓz#U{'�
QX�F<j�/�J��\PB���Li!�]��ǡ�g(h��>�%�PۅH���B�u�f[}?,;À�j�N`��ɇ��^��"�Zz�A�14�N5�A�n�Jd�t�V�WF+TJҽC�����G�ّ����gv�C��{�pR�����Dز���PѦL5���~*}4�Us���$�xԠ�Bg�jr{��0\h6�Rf���[�O`��)%>	~�����g6��ی�2�[��G���SU~Q�v��԰�`�z���K�;tPƦ�P;Ӗ��������vB[�.%e�~�� �g����)K6�3f�D��'\�����/%�憯1g��ڧ�u��?���R3w4�?H��r�w�߽9<���&�,���pے�ˢX�!I����Ffh���g�!~��x�^t�|�2�B��V�<�>sȼ�e0r_n�f��l0����Egڹ�
�=�����yΚ���j��/��������]�Ju�nxme	��dW�*FE>�wa����J���X�(�.9�� <��`�3�1�h��ߓ�тM{6�&���#�V<��QZj
�~"�dP�ɧ&��Dr�<Uv5H�&cfo��ii�;�9Ě{<�[D{:��Ud6��h�B3.��%R��#�Ͻꖻ�k��!8��8{K|LQg�z�9̄�K~��9.��N1,x��=�^n���;a�}0�+_T��[ɮ� ��Β�6@V*�0?��J�4��n�Ł�(�fB\���1���輋��n~��?`G$~�3&���l�k�����m�s���My��g��=Vg��7�w)����=¯�?�I��mM�Gr��l��Sz)�����}��F�͊�Y~Ј%!��\�Fֆ�b:H�F��+N��T�(���-尊^w��4ᵯ�3�c���������"s��3���ܘ,��N�u3�̟CìqV����Xf3u!���T��F�-2�J{��J9'O,w�D�/0�9b���b�#�" �e�{P
����ks*�w�&q� �T'?ˁ.<����!�_Yf�P�
@t�<�&�E���?�&¾y����I*��ih�z��� �5��<��D�1ōTq��9�Y|dw���c��e�ZA!e�&��RRl�6��~l�Α\�rսlBxܥ,���;/��i@L�ܬ�~-�9�=g�Ƣ�s�W� 2F��$d��7Z��W�8/��"|���^);��\`v\��+o$EY�n
(p��ȱ�9����G�#q����|Y:�2�A���i�����S- �!D$���<Wzډ֏�GYu�zn�ں�ت����Bez�����
�bN��<&~?�u�Q}�}^*��`+0��
R���<u6[������_��Y��jLZJ��&�mHU�Q� �}���Ff�d(�$=�z/4�|�_S���&�Ϧ�@q~�B�Њ,����L�ўu�$��a��yqKf���|�"��ظkX�&+��"����2Գ\��*4��L�	\y���M� ���y��'\H Y
�6�3�[b�c��Q�D��T���p�m��A�E��&:^e��t�֕��b�u*���e}W5�y;;o�O����lR��o�~`����vP?��(��B�K���{���e��w3��>!�� �kd�vi������soE�#�l�
yv�+|��	 E�m؎x*݌Pe�g��V�s�oI�s�k�37�Gn���O�(9A�n��"���4�O��Z�I�ڧ�"N���|dE��"t=(AM)>�U�|����o�t2�{�O����N�D���<ʺɥ~��(\�58��x��-�]Gۿ˸�LP����E��p~	}4Z�G:ڑ�t%�P�d��1
!�]�m�_��8Ҝ:|�]V�K��2�
(�2_2����X���Z�@�97��\7�VՍ�V�
���R��{k��0騄0�~.�a��{�	W7��s-��ޓ�~��P&�H�|���F�R8zoq8��a-�M:�wF<�gl@�z�}���*WUS���������Z�B1��S�[8�n����Ν���:̩j+�x9#�#�#sX��
A�_�V#ݦ��=�
N�C�vR�V1ލ���P �owN��w7:�J/�m��j
nK{�������V���g:�[�t�%���ܙq��g�BuhS/w���tQ�-gT �jrѹԡ�8�g���v8��� �G³���4��݋��������g�f�(tjY��|��ۯG�אIE���63����~�y�[�4ރ�����HZk�^��>/���>VQ*���/��NS��/,��j$���þ��-�~�&5$�^.�"�.Gr�F�9ٓ��/E��g�x�����Z�&��J�V�����B�����&X�/��n��U�(���󮾞��d�۟�p���i�"0��&�A;�Q��v�z��3����0u���]���3���!����-�[ɷ'�dPa���-��$����Y�ѱ���Qw1�#�.��Tqrr��eK�@���܅d�۩�R�c5�c$�Kg��LTW6�(�B:�-�(5�[I��~�JL�g��5��UņTN�"T�7-�n�J�5��q��HOx� �q�p��8g}��t������'�Q�Ɲ���I�m�@�9��t';E���=��c�i4b�`B$���Z����������@%���	l4��?&S�31̬>|	�<n']�� .���l���@�lp\qU�eۊD���
EWn+�1	���{"F2�8�v6��X7�O"E�"��0yM��SjV�ɰ��u�ߺ~����rq�巧uo�l�)�o�o����w�hR��,�63M���ő��X2ҭ����!Ǻ]��2��E�ʺg��:��C^p�=��v��`�}����+�̫�����qI�PS'?ۛ*L��%T�(�)��Q�z�����W�i�?=g6�X����X_KSF����UO��o��C(2/�<Auķ=���*<3h�S�Uc �\����#^/�Ҫ5!5�i����~H`E�k�k$9꽅�������y4p�u�UknJ�Gr�N��e�x]��ǥ9��we�w`�/��$U-θU�Hd�t�b�`i��0�M�#6&$�q�#�7�kR�f1#��X���]δ͏����<2��ޏ���1%���d[6+�&�ă��i������;�^c�vԬdn�/^�� 9u{ɀr/��W�������;a��O�)�hJ�	^)�]��x�ߢ)������,R�&Ӟ^��p����bai��PZ�T*�q��˛�J8��]�w����\s8j;[���:�.u�۹�&_J|ٟ|^��� ��+;��~�f��� �M5��N*�s��6 ,�p�<s�@t+��v.'��SxΨS/c�����|�`z0N��m	�7E�9�����u�+�� J���/R}ͬ���9׶P�Xkr�%�f��[)��oOJ"Yoi\�l��(��H�h�����m*i\ߖE
E��'�Z�u�荸_�s۔��)V��l���	��%xo��*U.<������IFr�gO��Y����#I�x�����$t{�HE���e	��X�u%�b���pX�c]��ۮ,�D�ް���})~NU<��4���9�����IW���>�t="ZdR�q�qG��F���k�O�@�d/=q�ZI����M�ɠ�.�a�*���^��OA���scpWъ����:�E����=��w�po# U��L�~����a��Ɇ�w���6��g�3��2�w���ΐy��b��gX��4�F�^�TG�_.X��VLZ�Wk))ԦX�|�M&��=�?�}����5,�]��	�`-�q?Č)�zJ���Jh�g'VX� ��*�eZW��	��;�#nD@��rw�5i���y���������l�H��ȷN��F�9G�n=�f'l�MGT/�i�d]
�!ZD.j��L�U���A(��əe1�`(05�9�pT�:��Y���u�y��6KR'��<;ƪ}5�i�&����'�?�81������ź�/6\�G��Ҫ�Kh��w����sq���7�?�Lz�������TU60�+� tc&hg%�d�k����l�q�`MNf�9�r��&�}�<<ǿ��T�CF�	.�=Xr2�Ӣ�k��v���QQ;A��lA���0�n����?A���5��
��h��hW*�}�x�Z�S����e����is��.����s\�O(�����vh%�3hxg��j���,p�	4bZ�l�:���`��-.������{h
R�OmP7T�a�7�OMo,����j9R����1h#f�F��8}gEF���$���:�
���M��̉�22���Q��`�ౖFp�Ap ��ԦϘ~,�9��3>lb�6�p�������IX�|�_����*���3DF*��[V�ֹ��ZM��D_$�N8�Ъ'.�f��S���Y���Qj�'���~�M���3�Aݹ������5�[`x���������L����&��D�&��a'�p���{5�,��ѩE�=��"� �]X�k��c !��&'�R�P6b�^z�8�SH�#�25߾@��Ҳ�t�D!��ɧ��e�H5@3���D��F�����4���x�[����ɍ'�w�_��F�I�H�=����ׇ�����U�z,럌���;��)�ڪ�^���TB�C�8�w�	1���ٮ���sO��V���$ZΏޓ<�*�u��ӡ�钔 $[�`���QA��(t1�J�
SA��d9q*�Q<p�t��m`p��͡���9�ĦvY��I[O��\]�m�d�|S�1���+�o%kU/F;G]������\'�|Hg�5���߆
n��}���K�4�U��>5�5��@��zp!�&�]��<�5m&
阱6|�����P;�h�T<'[8hވ6��T�'�7�T�����K���1`\�ܓf��}��"J�Q��eZ��`��Ko��/��ƾ^�?�j���	���#�T�)�IA�J���j��窬�g�A�#T7X{ag�Z����Ê˳��BG���T�].C�Lώ^�2i���i���8�<T��L�B�b�C������ŦxeQ���"l�m�Wn��[��I�V1����&<���:+�4�a���n*�q�^Hf0L��pC]K��暖"MM�۔�}��)�1J��x�"ү����;�d߄
w�a<��Z����ת�����x>�]��=�@�2��j}DY�1P�*4ud͉�j��˞��i�S�b]��6\�Y��c0+���ͽ�b"��`��� �ܑ�4)��'k�=-��-�v>�;�R�1��M���/�'�x�U1�v7�j���m펯���T��np��~�.��=��EI�~D�c�a\3̧I�p`b_(�q���4=lj�Dʢ`���?�-hH��O���V���7\
��5�z,��ݵ��-ɇ%�>JU%Ѳ(� ��
�tF��V��{���5��RJ�~��p�W�tñ���n)5v�Uu2F"�V0UU.�%�W��Q�C��j �ޖ��	������TBD/���~H���ZMN�����S�Ӹk�i�Z��M��}{y|Vbhч���s��o�]į>눴��Y�	K�<6F�Z���ܒe{�2u��>8�\�QX"Y$h0j*D�\���^�:�Y�pƬ]��N�:8�a0��j�|��h�����-��"�n��,V�kۈ��!Ot�}{�E˗��ϕ�B�j�$��W�Y0�
�5�������GN�,�i6Vl�*�ߞ�}�/1N V6�.u���/�/��;�n�e�RX����_r�4����Q(��k7)a~*A�wQ{I���n���ɇIG#E>�6#&[$�����u�~?�䒞0����:��w2|��2�l ��K ݩ�����]���wm�|t�#]B�a�u�Х��Im9Mv�7';g).�I�n75����c#�c��=����[߈O��uu���F8�:}~���$�d���A��w�}�koKM��'-X�,�� <���5�_���E���ͦ*N9���.ܕA*���<hњ/)�)as(��,�����dy8l�ŒL����	ŵ\8���p&5�����Z�~��z=�7�`b�D�K�C��I�.��TV��|��B��#��W@k�G�#w�E�}()��7��Y�@JB�:i�~>0���4x����A=�-qo�*��Y�%��L�D��OŘ8�)��^�2�8�ZSsY>T�&�.�m%�³���&&>9Gz��u�Mo��A��������w9,9���U��X���˷Y;����������n�Ü�Z]�O��,��J��&'�v���i���$u8�GX��*���^@t�p���JD�ҿg���[���M!������.ml�������//g������� OGUUB��ܩo�A�>�Z�o/��A��k�����%��b:��B���YWA`�\��gȺ�|�LD���W�2=i�
�v��Cc%����)�k���H�G�u�=2���.�098�߰��\�ʏŝw�m�,��"���sK�ءp�IX;�/��ZMU�+��>�s.yR5��~{��z��C#�6@P5YU���F��-��p_y���&���i��V�,��
��Ɍ�++��B-�n�.�o�}��N�r��@�v������fDf�t��<�\Z��ן-�W�G2F6X�)�TJ��9
����3�:��'��v]&��`i�y��z���K�c�|ʎ1��Y��׸�\h��T�R�D��f 1��2�U�k�����,�EP�^Jc�|X�ä�� WI-'�! �gPK�ڭ��F�f*���f]	Q޽=t���,������� p�� �ek_�Hݝ�^V�!X�VoNt֒��z(����(�h�uPW�P�*�vV"�ې�lS&a&�o�?V+�_�>�`�fl�)�t�Mہ�m��Zǽ�6�à�U'����r��c��(�����M�n��{D��f�sLT��^b���TЦ	7�l7%P�
^G�F����T���0G���x>�_R��\M��հsOe�:�[(� ����3�����\D�,K��}������߮��-1����q_��6O��}�>��$��D����Y-�zX��ܹ�8I�q�.��՗�����Z��P2���GGS�.5�B3R��Jވ�j���+����^9u��n�=���P|a\ ��/ 􍑞a'�/�E��Ĵ�;�oWeԲ�H;�/7�~Bf4w5�@�+����d�{���Z?�@F�S�[��� j}�b����fq+�4:��l,���d%��9J�³��
����V��(k�#z��l�hB����,��;l/8�9�Y��mi/�]t,����a�3=����B�n�[g��[S��m5A���֕zU��t�Z����� ��+~�
��ߗ}��g��̌�/f��xύRW�-��*�-~D�z�
������,�*���|%�trU�Ĩ�˻�_\�)<P��,�o�ʱ����l��Nk|�̜��=�}6N�,�<1��h���aOsM���>iD�\ͬ���љ���k,"^J7���B=�@�o�����	�xC��K~���?4m����Wd ~n���J��i����	�R���B42��-ę�#_���ۼ��«��}{�R���5Qa��K@�6Ʉ�����̈�sz�$�UT:��ⳉ�����ͺ�rp,�?\���XQSbsO��雠��!�����q
�b5��Z�����}^��r
���\�l_�9�I@�p�
��5q�u��7Ĵ������,Wv�T��_���aN��~�0j�.
7(7K��\����'�|�邀�r�G=��J�*���7�'�KD唣VŴ��.�T�c=;|R��Q(}��wB�d��A������~�n[�F�A0�N�Z(p}ң��\�r�i*��1�?�m�JRxju���|1��g�Z51�\JQ��\r���og�l���	���t,�-�F������Y_��oI>ͨ�Ī`�kH��$mJ+G�֟Q�׈[ba�gȽ�t�f��|���YF`��EU�8��PU#��۠��xe���6L}��XǄ!�ďV=� �FgVx��Z�	@�R0��(����i��8�-�z���`pPtS����P���)y�����P�t��>o?��вblL������CnI?N';�2s#	��4�r6�]Ӛ[��e�=K]�[l��KN˱�M�	`�}���Y��T�
��qQ5���%Z� �o����|h7���juߐ��8>�g�ٻ�t�j��Nև�A�+�[�!��M����;p�f�<O�{ �$�����gQ�P�]7�[,wt�:C�B��es@��~�nА@A�z3���7g�à���R�f����'���a���"7�+�e�$ܵ(���ia�iU�;^���h��x���Z�ԍ�=}̅�<�Sӏ�֊A�1D�߄���ɯ�9�tw`e)ua�Z�f���rǋ�(=RK���<������\����)�O��P�UG��΁6#d1�2���ݏ���#����dl��8�aMĲ��a�KI�� gj��'��P7���&CJ�����T��1W�����+V����5��y�9}E�7����� .�
[QP߾:���:Ъ���j�i����!�/E�U�,�o��`�~Sq���
ؠ�ۅ�*���cr��<�,
9����Н3f
Yr�]���{�`�c'I��5����[��zgܐ�;p}Sbƌ^��bB�w���v�!���#s�%��>��w�֭�(�b"uO"�YN� �����r[^y_���*�yw���.�Z"�m,������>	4:�c�t[b��]��Eޝ�g�ń�*���e�q�O�D13�7f0OחU�kg��8��V�J����݇�3�{��9y���b%&�L�ji[�ՅvҖ����}�sxx�K|#[�\��E	l�1a-�����#i�^ѿ��rV{�#���������j�Jƒ��h'ʐ��8dN�&���ȰBQG'�'��0�k�\H3_���W�����Ii���n�]�u��d�~x�CU�}�~�t���ܧ`˕@BX�{��1��r�*�L���0�P���5���� *��Mz��;�#���?֍kxF�J\UP�����\��< OQ���˵HQ�o�3Z27�&�d!6E��L'�A�;pވD��@��-Y=W�%U�V�Q�Q!�cI��W��Ĉ���oq`���r����'���__¥(Iq�1��.e,'���8��.E)8���o�MdB;�Hj��K�<��򎬗�el �ችEǃ��]тN@��:��0vP�� �e����a2� 	�t�����{>�è/`+�����3i��a����h��?bzn��X[�'�X�Rex�`��G��Q���P\�{�1q��o��U�'�?%�,�o��`_/Q������d�}�.#x �缨�4��.Q} 6 �b%1�kn<�uMWү�b�g��4�P��4/�w�`��fh� ���Cs��ņpp�
{O1;ࡨ�����N�0���yW��g3,�@�����k�J�Om��^��/��t�J{s$偕��r"�(������'��T=x��G�ta���V#�(�����T�����a[�w	+P�ʧ����h��������/+�OK%Bf���2��إ.�)�a.����홄�.P�C�vO��TJHo��YYd7�SAT�����]h`m���6����5V˖�5?D61�'�B!���X4�|��A�Sk+�D+��w��Sב�*5�\5`SE�ūɢ�N(G"�����4MH�U�������R��[�7�β��s�伎[&Z
2��m-�Y�/Š��C�F7j�l�m#���k�ԣL�#bY�}7��w�:k>�gFx�Rhu���%|���޳T��"%-��RB���7OI���؊�l@��d���*%yd�ࡾ�8)$4hQ�M�O*���F���l7��[٘՟���eX8bn�y���/�_�QF߸�u�!3[9~Y��͹����y�O����n��#�}b��`����h�m�;�/�|ŭlAn�-�x�,�+ks�v�bh|g`�Vɩ�՞Z2��#�V�i����{���p���yϤ�X9p�䐬��hק���X< ~S濬^��T|�3�qn�J_�h_j��+�m�b~Lz+��`��hٵqE���*��N��K�Q1q�<�B2{ԩ�&`�tXt�R;X=j��*������"�
2��j�&�r��	Y��$IN8��XN0r+|DsC�x3@�}ң=���S|ͤ��=�c/W�~ ��z�2"na+R�1ҝ����$��tWڎwI���j?c�!��$Z�L�G%��:O�g4uZ$O��"Z�m�k���՟�cv2���g}.���ǫ��al6O���;�F
B:�e[��q����=��ô��7��n���Y���� �m����Ct���8D���Ǚ�/��U��VW�)�=��S2���<r��_�������·���m����1������	fJ�J�3&�H2	RG:�U��z#�Ƿ����s(3 \�=�x�~�	
.�J�{`0[�@9�w�I8�C'��~L��EKJ�x�	��"���Y}���Ci����M���,�6RSpx�o�M��NUP�q�$�ӷtu��Hb׈��Dx(�T�|	:0N�@��% v=�W��ŀa��*̫���`Sf�|�]���Ya�挜����'�S/s* ��O�3�	�R�`9Wy}�B��]��'��	�����
@}�Z3�,iN*��6��L(.=2{(0��<k�U��5ˉc�-֏h�\���Q3?���l�����Q��K���Fh6�.��c���7��6G|FZ �$��#:Soy���(����@� �; �d8�Ƅ�T$]a�*��
z� Ǿ��C	��zYv�;̧^�(΋c�	��{r�EYo��C��Z�,��,��M+\�:�L�X�^i^��s��vg��(#�f����%\���!5omX�\�R��WqK�*h�gR�^漄CY���Oď;�������}�3P���94L����zN�J�=���'(��C���bpI'vOO{~�*_F��׊팚�͆�e<3�d�P>];��?��C}�c������ʁ08��X-|0�G���U�b7F����H'�Iv���]]�&�D2����$!�h�3s9=�K�
,�[�y�r�t�Qb�y�7@�������7�I9�	���~i��>1_���n��q5`�B`	YG�t���ݦv��T �^jNyJ0b	H�܌��ϯ�5B�>B;�f�mKMoK�?%@~��7<�qf<���B(�DW�^[��eD�I�!�='@�ү/���4��]�0��mW�)�xpa�w/I��Mtי�6;}s	�������T� !^ � ;�r���IQ�2o;���gۜ���8�<��4�23���Cs#h������e�$��4���˹a�r�y��}���ec�6�'�SL>� ��VBc=�tg@ƫ����ݝ����4��~3�_��GӢo6�Ѕ����f���ھ��a��ݹ1���e'�����Z+K�l���̎+�Z=ԟ�ڤXm�'�k���T:p��%���m���o�QN�}/�\R��X��3s_V>�Hv�����@�a`X0�V�Y�!M/�6�d7���q�4[�&�
�`C)�_��@�c��0�����_!Qʜ�b��.�0d�� �9��ՁR�l������0w�O6+�}�\�.B<��=VA� �]{�AE�vZ0�doK�乼g�[ũ���\��aM�r�R�-��tO�l$ a{(�w(�	�1�5���W����ؓ� Q/�{��m��2�v���1(iS��f��ޭ�q�(���ZC�ږ<��|�fJˡQ���n�ߊ�|B�y�D��t�5��[�����8�U�2�I޹�}�K��S�Te|�W�'u��o~������Ga��{i�3%��r�=����zǯA
�s@�������/�̛���+����&p+�%c��Q4��\}�Q��!^���1�!�^��j$2�G8)�܃n�k4��,�.���J6NMü�����'1���E��0w@BBR���l6�Y� 2O�ؐr5�5�C����VUEf0$4g�\�ݟ�&����;G{�1}�วw}�nÑ�ƢR�3Wtju�Xn�%��;Ѽn���}��EȒ��l��>9�1&����%Em^`��^(Y�Ҁ�*�k��	�ͲMцl���F|l�FL?C���BbGA`��Ԏ��ǌ�pdLR:���Ǻz렜S���o�!�rlu�|o'���xҮ��/��j�d�m��LN�9�Ea��m L����.~���)�G�wk��鉧�j"`�S�L,�{�QeKD����;�%T�y�|~��1Oσ��z@�j��	kP�J2fU�1f�5*��K���P>3K^�)�����3�F~��8�m7p���C@���{8ϫ��^|�Sb�k��>��ڑ��r��Ѭ7Ћ
�ہ��[>]��V\��w���>��[}[Ϋ��z-�\�-�	�!�ؐ��� ��(;��Dhqq�&���1ڕDnRF�=�����>\to_}��_����1*�<8��娢��a�,�a�ԍ�ޕ��"��u܁v
���$\�q�>�0�R5;�Eh���^s�I}�Vr���a�;
�%\8�o�n��Ɨ&�)D�����:
�E^�o�y�Vˬ�,����>��Â���"� [2Wh��T���X�5����t�;�x�YvZ�s93l�fɃv�q!��3a���e��My��-�\�@��R?�yN�5�[EqH�k�L����+�kqB
� {�����JSM4H'R3!���?�|�)!?��/g�?@��(�`�u�te>9m���Gs�6�ݘZ��Ͼ�9��Tp��?�Y6#+�\W���3��Y庅�ѩ��lw=���ѽ�5�A�f$Z�Π���r�A����#7�5�]��O)d��?���Y�%��5���9� T[�B!o	��&�l���K��K�vU�aY/2G#�Q�X���XtA[� �#��=l��O�T�
��=-�����/g_�uhJЖ#�O" ���u_vц�Ψw���e2��0����_R���EMlZ�?��\{��g��I�}�
B���k�a!��rw�썪c{�(�,�����!��=YX�_c�ɤ�e���l��Q*[kc7_P���|�I�LA����b0���;:�d��<QS97��Q)�p�2��o����+G�-��Ӥ9������#�֐�����s�
�Yz �V;�ª��a��I���NJ҈��oi(�E�|(+��H���C�z���$�V\�@s�^0�ӂ0D����W�G��Gϙ|X����#Nl	��罆>�ԙ�^�����K�(+Ynb�ncXvTQ�i<��_�S*�©�������
4�c;i�������h*�KJl�,�Ln)?�s�^Ft�a򎟃��Dg|�d ��,'L~n���ј6B�x�<\�6����l��$~\��	�.a���?��!N '�$���' ��A�[�{�y�#5~�.N�TX��r�B<e��X�D�ʃ�폗%�W;���Z�r�O�l�}yy��Yʑ����X���g#|ဪ���|�fX<��6#0����{Km�j�O��L�ew5n(�Q"�6�Q��~��VPo��#�P��LL  [�C*Q��"#7ω�9N
�k��md�b(G��$�`?Dcs�<#�z)�u+��+.��k��[�������`�B|\?��U5)t#�y?Ԃ��&��>�qF.�{� �U�oUt�#tO�R�d�N'�g��w8���k�?��N��N��6��8�������U|[3Z��#�Z`���3T~h����?���c�9�����Z���U"K��Z���J��a�i3E[��l�X��1ў�c�X��z�"����|��+a��m&�P��f�J�ɹ��՝JDC�zb�_��	��	��h�:Gw������PĨi��%�t��]��� P�3�v��H�۰*��(d����6��ۈr�Wd��̈́���RH�Z���ƙ�|�������߭�M��鿢wpc[��*A�n����	K:P��d��^���P��)"9�l�D9�t�0��S�U镇Z7ք�b��
���Nױ��Ku�[��q����Y��BŻ���C�QL�	Ĕ|8�5/S�(q� gr������ l�����@a�k�`����( ���̮C��İc��L�4��i�or���n��g�i�]xl��ҎӘ�wx�Q弰����E4Ⱥ���вAƓ���-E�2��c�!d�|*�<ţ� n*ˡ��G���ԇ`�D��ƾl�b6��3ń���#��`�0�oR=��@{����ib�$� r�p��{�PބP�(*{J8���_�k��N�x5g�����f>Q�w�r���Q݅�A���+�<�ۢ�-�.M�&��"�x*&�k�*k��O 0}x>c��ŵA ��7��i��g���J3�I9�}��˞��?�P�9�L�r���s��e8���ᡇ���5z)���f6(J�˂�@����J� �/]"���쓩�ȿ��O�/���WZk��3xgrZ"[�����$�a�&������n�J�4T���M���^G%�Y�;�[V=ʩ�CP�}����_�I�l��Rڑ�7q���².���H�m�N����U����?jv�_⃍GÑ��JIհ���-esq ����M����(E*�P��#��S^��_(P�X�fo��:]�H.m����9�	��9�/R�0s����y���a�[""b:I�ۈ8%�}?����Yea"��U�X}������O��#��.K/�`����Ս�^͓�.�{��
zeF��f&���W�6A+��<��h,�$,�xj�5�,s���:�.�y��oh���'�0�9x�u����3�aؖ+�|G�s sW�.,����:�g5� ~�-�F�������'iWpA��4�ݮ)mI��|ƨ1��R���.lE0 �q��e�J]�Bt@e�z��iN��5�#K+#�r�> ����!��.6B�2⯸W�|?�
e�P�j݂C�63���^8݀����dnz����&CF�2��%�6E�b�����_y����r�l݊e5���i(��0������dV�UE�Q��W�
-��ok�xN8B߂�V]5 ���=/qQ���w��ٶ����m,��S
L��~�geW��uA���.�U���Cx$0���+�{���g���s��a �Ym�-ŀ��a��Zx�}]HUbTO��I��*�8����PZ�\7t+i���3qf�������x�}�ᴯ��Cx�LntrC��Z��4_ 6���*���{��|oYO�sHB�>Ҩ�jdo��#�r��G'��n���M�$}��?�=���Ś��t�p׋��?���uW֪r'����Ż}T�c����I<�ͯЧ96f�k,øMW;���ʙhy�Z/����#bHmqWͺ\z�AN�l��?���.�eq(�~��%�H�AbJi	fŘ?(4`d]>�,�K u���E^t2=�T��H�� ?b��ҕ�W���%�{{�l��ۚ���s�0�����PI�[K�,1@�\���vQ��8^�{RRCi��Y�?���%��������@z�tjR�*�|Τ���TO��)\i�<�N�Ug����M�4�4?q���o'VA�����n�^#� y����;,�Y��P�Qj�����RÂ�$�^�f�XAW�7��πق%TH1ظ�P��u�&��vǝ��.v (�/�◞��>����^^��%NwB�
@3���n��ع�%���3��>@���p�?q&�+�7�]�W���>������0�̚��N@�]���jdl�;݅ߥ�k@�O���wΆ���/jSu�y����o|v�ۣ��ݑ�����-�R7�L����}����h�x�����$P�I�hr�s�bL��Dub�2v+���W��6cknШ�L;���zr2�����Ɗ�aS2��8c���U~�(,5&�]�b�S��Y�b�9]C+9~ލ�;��)����:<�B��Z��_�re��
>�|�紒� �=4K�&�����߭߻ux��Yз1Zp�����s�g6d�]��
�x.����U�P�r����^Ӷ�C���酮&h��,7 ��@�4��P�vg[RC�.cfL�{Z�7�=�:���9|�K%���D����T4�l/�륊�/�y��+���>4Yb#��c�=%m�jR;(P��}�ր?:-���&�. ��uʊ�Iư�����oG�t���{x�G�Ļ���޹6����(�07�;�^2�����G��ن�H�ؖ�O|�Al}��� ���s�/1���J��Ʀ(N���P�{���ZF*�N|�d�����b�0����lh��9*�LF+�!ƽ�WUJV.(�{j�x7�Zx���Bb?��
%�=:�%%L���Zb��rN*/[4D�z{C�2��;�w����:��64��@��X�NP&M��LxI}������'T��Tu#��Zu��'�:1�<ɻ=�σ��:C\<ݚÜ۶��+LH��P'Ք[� I�$
�i�aRS0|W���c�3�������Q_^�߬�J�\ ���z�lG�VU)�t�*ϔʂ2��^��:(��������u`V�y9u#L��lK9��=��I��y��>��.z�1�ƞ#�vu�!z��r�]�0|x�N��^Ux�:�z?{"�b��%寸Gԡ�Y�^B�1���m�HѲ�O��w�W�1��ϩ^]_�7��f�����ߠ}���{K���'���ĥ�� w�@�eW���᧳J��J��QF��B�� ���|>z��Z����&Ej1����cb,8����m�s���A�S��5�ؠ�_q�����,���Y5��u������f�*^���[T�qlQݫ��P��W4<�'6�c�(����T��q;G������WZ� �e~'2�z0Hƛ���s�n�W[E�ҫY4L�=���y�ˤRB0����:�.��_u�Ǫ۪���k������9��;��ޜ����i�6�<fL��āw���<QEҘH�+�=$���R
<��Sm�qL����i޻1���F���C��fYr�H_[��S�I����Z�v�3��Jy�g^�`W����tȲhT�πP9��4�k�r��������"&��!r)��I�(a����bW���ўi���W��O-֣���E�'H��P-��z�[��
@��A�?ц$������F���ε�����3<\f�Y�`���r��ں4��Y7,f<�D��^��E
���Y�wV��Ngȵ�פ`�����q�y��Y�ܤ�J���8��BiA����MFR,�/�j��|�${g�@���@d.�nu�A2��G	T*\j�Q~���� ��+{4�N7J�1R7�"��Vz��n0ߖHK�8=����_}���a�s�H�M�������p�e�c�z�*�w6��o�[�C��#��s7�άM����Ǣ�"�)�����1iAщ
!�q:��R�w����}0sCY�PE[!Xu�̭�r�ب~nMi�ki_L�O��6nn��:Ĳ�� ���[�f�~�r����C���U�H�F����7����R�ޗ�׼9v�;{j]�:+&&,fGu��$r૔��c�f2�r�P�n����騯ݷ��C����?�~6��=
8KA�0�d�퇨�M�f�`�Wo4cq�d������x�#ƕ7xNm��T-�v��F5]�i�TzG;'�,V�A�`����;��������j`5�BK�� �fP��}b�Q8�_nhjr��P�^��/2'-[�r�2_	��l�8�a�
W]ܻ!)~6|Y�8U����Py-�����0���k](�!��-a ͊��Fe���X�9b� *�$�����!I�xm%�W$ޅ�#̜j�e���ÿ���\~��<`±��������!g�W���K]�3 b�dG謨������.LO�fO�nU���Qے���!��H8Ϭ�e>��5�;	)RF&�f�C'Ϋ0�6⧚?Hq5l���U%H�H̃q�p��kģ�=b�0�ղ�]�Fw�_��"1�������M�7(`,�{�;�/f��_m_ �po�X,�Ԏ�۪T�ҡ9q����V��8AqV��F�����Xħm^��h$E�v\�(���ӑ���[�P���̦�lG�R���^|Z�LjY�����6F.\Υ�u����^ߍ���t+�T��5,��u��e�T��Ò�ZZ����Ŏ�1+v�@��bL/NlZht��e׳q���
2ȱ���g��:�������V�}W� z�b&�0.<��u�@�9'i�Uq��3X-�� IrE����z�wDI^�!;$��ؔp@�ܢ?�jp�0滤-l�2��L-$�� ]�
hȢ�����Mr�¼�w�54���{$��0�Bl��i��!}�*���������O��G>h&>{���%�D��F�K3��Pq�9�}0
�D?j3��$���4�j�/��"ױ�X�N��hm9�/�p�=�8͑.WxW�-�Է��s��]� ��'Ucp@X���q�]~���2��43��N<9|,8�f�Y?��x7C�y m�V'X�$�Ԕ6T�QV��D�$F����ޛ��vYƠE�_N�z��RQ�����2;v�UUs�yUf���hy�r>�z�J��h2dǮ~�aø%1�e�Nа%�oB��P��2ظ��)��f���m����ī���	�;�s��)w ��C�a�����=�������&F��^)��$Q����嶲��r�+��k]��c������K/���* ��bGvfI�I`DS�A?�T� ��ߪ�;e����NY��~�[�� x9:����t�;%��W��tV<����牃�#��r���i���w�Ԍ�2!�v�p *���N$<���M�UEX�#ِn���E\�p!����f�Ε�>���_r�Z��|<�LI�j��z � >�S���Q�ݟ
APK� ���X��zr��܍�����ξԲ�1��Z�D���b%[R=D�6�.d�ov�_bG���s��_Nֆ��tE\bV|��&�o�/����7܋"X,Ęy٢C�<I�<�}$���T
���oe,�ÅQ	�=7r������G������|6�$�}�3���D~�1BM~UGkvCc69z%�2$�b(�L��]^z�#�m����hwh��Z�P� �"�g�Q[HQY��B�翿���s�]Շ��d�};�43�KW�B�����+�1�\=�J�� ?��=9]&g����8f��l:@�@�ps��=S�&�G����P��!��Q�.8����RlP�ڇ�z��g�3��A@�8,~�� �N�ɴ��a#E9o�-���T�P�OnLS�����`_��3agϺ;�X�؍����v�TŹh��zjȌ�ۗ%���̋E�c�����I2�� �� R���O����.�������K0T���oT��P��	�'���t&P���3�]�G����ݯ���B��2�Z�Jn��w?�@�����M����Hsjd��%ruk�(:+�,�]������)���ZP�D~�Ƽe^��/"����<�qO�;��mA���{��!�kR4[���e�F��_8�$}9�� �Z �s��� (,^���!�&�)��u��z���������'J�f��|�&�MԵ+�o���Giq�����lpR3�:��|��vy�M4j�=l���
��cds2hg��^�t|�T����f1�i�@8�
b.l> ��8��M�t�IIv�>#!������P�I�:�-L1�������ʮ��l(c���H��u�*��$8��:��7� ř9����E;Z�������N���4�q,����7Ԧ�]�OxΞo�ό�lL4,Z������I+	?��E(y,5oP7%�����@����ŌkTӲL����ʟ��L�y_L��������������6\��'.F���_%8_,D+}���mJ�7GO9Uo��E��e?�fmc�eB>������$�xԂ|��]���~�yx�������-�C|����u�z�`��-|�uQ��_���o.;-� :��6�X4v5��s��y-
� �n0Z/�u
�T���#|f(���ౣ��w�� �Z��>YV��|��Ё�$K	�=���L�gɄz�t�6����O�_�U_�b�6�_��p�����T��z���<�&��Bu�G}^HW%��"�¤�wg�Vdh74���V��>������㷡}8���*�Qh��TTn��^��2ɓ?/����t��9����r�8��E�#��"|����p�h{��`����V�%��3�`�B���ɄKl�ާ'�ҧ6�5=��7�t?�y��(*��f2NG���WD!1�:g�Y�>��!}�t1�!��p<F�Ll��6�����ls�h=�ذ�, 0��V9/[c�R���F�x�Y}+�Q�e��+��w�P;��(fo �@V|͐$�T����&ظ���4�v��5c
�'��M�)(���]`н��cݛ1Ἥ���V�@�ʎ�WpU��U��s?�v�5k�[1|��� ����ڽ�Z�+��jk���5b�e��a��8�n?��z�(FB��k��P�l����e�[�A�~C�7�˷$�Wx<`u҉��rk'y��Z��Z�i��HJG��i��/�>>+/��oBp�Q౟/����a�P�6�eP��@y�|���VQ}��.iJΐ�=JѴ���V%M��ů��m�u�<���P��.�'�F̓{�HlC�H����XP�/�|F�U����f����t/Pu������B�:9����=뗳�-�{��E��N-�R�!G_'������y���v�?k�<�{�u	J��@��x���E�ֺ~+�$ov����e>����m����JMᬏ $o�굔˼��G���ر�s�#	жc�Ѻ"Vt:��Qh��j����W��
^�au����>�N�P���A�l��H��2�W3�1(������ݚ7�;
�R��a�����4�������s*�تR�,)l�
��ϝ�
�)��T%K�#d�f�?iG�շ�[dѣ_j����s��@P�:œ����4���^VE
m��p mPx>��Y����X�D=e�z�����LNN��(��x����8��ޝ��0�r��XUXI�݀�ʾ��� .w�Oi�!��ٮe�B��a�xI���r�4��7Ҿ'B��A D���+���N�j��F���k(�7̬3�	��C�Y�����4��]�	���\��n|X�vV��������*�#e��1�ö�]W/3˪���^����赍���Ы��E_̹�ɢ;�F��"��R���W{�i��i�����=����}����3����6���]q%KXSC��ð�N�gR�uOS��ヰ��Kw�P���Dr�-�A�j�U/Į<�g��<��7_P����k�=�� X�R�HR�����U��G��~�Kʻ8���Q�d'l�Ljސ��q�u��R@ ���;}���	U�3S���!7�vQ���8�Pӝ���,�`:��h���J]+��4c�Ũuҟ�ST� &o�m�f��x 9�u��L	@�f��}t%F5Xnk��=s>����	��1y��P��|i�~Y[g���{<�c���؁ ȟ�e�ڊ������.l�}S�ɒ(A �/i��_�4�J+������d[�-u����gTE^�h�c0��|2�@�_wo���I}KkS�*MŘ��0Ckh*�v�S���x�X/7&�[����&�tޢ
��;`>�ɘ�-@�e�a��� ��抶.���b�] ʍe!�q����f�O�[�6��'fC��`�29�o}�����N j���E�fK13�X�~��'�Y��c�P��X�}��K%9��^_t���wb1��E���tR���S���Xn*_�~
8\Er��	 \�#�O(Z�tS��S��kL=������.�)Bs�W"�>�������h���)�S�/�{����E���ex��f�r8��L5�6�ǀ�����{5Y�K�+��(se�T��--!�l��F�j���e^�ݸ�x�+6�b&�e��I�k�A��vv�l�q4��[�%D0��ح�mD�6ߝ0�r?iuo��~��nak�bk�? ������S8	O�C��7P�҉�����s�K���.3��D��.:U��W�`*�T�[�ؖ5LY�
�91GY�A�~���@��@�)��2)!�'���u�C/[n��L~�X@?{	�c
@Y;c�_��^��h�$<}?���s9:�Z��E8G���1v�C�toh
M!<�+�����ª{^z}��:�c�-�p#Z����5����jP�u�)��K���@�_�.;���`^my���%�͔^`�:��g�]%�9���LCՑթ�O������?��=�Re�&�~��F��v8#YCz7�l4ό��V�J�_k̬P�g����5U�j@�q�O18z�#Y5E�?�Ɍ?�Do���Zv�]@+T. ���J�g���CׂZ��_u�TŞ� ��߲gӷ��w�L�{�?J%~24F> ������8W���M'����%���J�!$��/`n���q��؜J�Clfy�A p�y�̾TV��.FBJ�cLt�B��+�G9fNͨPiC�u��W���R�F)�3]�04���/`e/�����r ���4u��$�U96�3*��g\L�]��ӌ��J]�ɝ�9�%,0�Zqړ�n��)K�� ˉ6-��^n#l���-�yr&�P1HC�������}����˩�9+�R�05�Y�?���aR�)�](��+bg�Ȓ�@��E�LpNƈc�/`��o`i���f�4ms�}�C�B{�Vy���p�()0�̈�AQ����O�d���L'�H<�u� �Tn�a������[����Ws��+�|�$x��gdk�����A;$��F3�>89�A�&�5�K7�9�-��TN����pױfk�^��PI
	(��о/�@*ዻ|��&o� f��C����K0p��"x�:J�y���I�2���0+'�7w�����1���]�8��@��)3^A�A�x|:٫!��j2��j�@�3��Ӓ?�"���p�FQ��f��l��Mb�k�s�Ђ� |�)�e�?�����)B���ߒ�ۧ�~��Q���y4ݭך�R�ܻb��z���}A]�GH�в������ݩՓ�e���B��xQ-f٦/�4�2�	��b�8��x�rr��"@=ށ�����Ŕa4T)sP���� ׇDۜ�՛ɏ� .s��b	q�G��W����D8�X�:Aѽ�>�D9���fy�ej�ٝy�1͛��nҘ����_\�6��!�뿩��n�Ktz�S��	~&�V����lio�W,`���t�x��_;�Q��PzTc�7�TI��K���������vlAw�Lou�ԟ
��N���2@L�)�\��C��fHW��(��o�V��]e�4�����	����Ar�v �Os'� \�D�I�ҩ�캁2��¾ ׳�h#��p��|�ۣ����9�R
 �9l��\\q|��Hz�~g���{(T�s�`|�G��n�*�k�5�>�?��Ը��yQ{1��|�2��V�czܕ1h��?������&9fU:�,Ch�a�E��	�w�[-��P^Q��D�u(�|������`{L�~4�h��3�Q��ك��c�^��Ӗ����M��!�x�|�r���ѮM<�����̡>�xI�|�'V�Dc��؎���!����+g�[�{0�&ߌ���M%	��sr�ajbJQj�9�V?���+Ґb���8f�U�e�;=�B�
����k� ���L�u��F��
<̡�J�\�znP���UB�f[HW�N��p��uo&/6���jQfS^xMB�XK��;��7���J�Ra�J�GV���V���'�ae�_=ڵ8���\qh¯�� ����Ӓlz%"�`$�L��g�'2�N����n��콬!���^�O��3�S�a(0˕�z�����>�Ă�����g��'�  �X+�������2��@��W�J}���EKWu;P맡�����Ṇ1�Q�VgصR��`�L���k�4Q���ك��d�_Kuou����*z��� c�H �f�����.�	aH�?ƍ��v����O^�`�����rsr KX0P^f
�?y�+5�j!U��-[��p�@8ȥz������t{���"ЯZ�����U�3Z9-mN_��ŵF�c����|)���,o�%l7&�����g��A�X�r��Z���l�Y�V���6�Ţ�k
=Ʃ�԰!z����܅-�fº%� c+'����J���H�d�f��\�
�|���0d�����yfjG3v�"����f��>��Hy~�7+�7.���w8�4�6U�{vN#�_�c�ڍ��#gׂD�VJ7%e�j��F=�����r_F����\i�;R�"�7�<���,�*s?�b��Ǖ�1(��܉�U'&�ۡ%�ישn��
��!d~��\`V�$}'a��24.��jT�^��Q�ٴ~�U��Y�n���M%Ӽ �,��߈3�Լ�o
f�eS�$�1�3�ywq^ț�7��Sr��βܩ�<śE���-�29]�m��Gr����gR6����B���D&գJ�!�������Dq}{�<Ų+Y��ꪈ������+�����'����2�l&��6�]��cs�ϓ��-��-XzNjߵ�z'��{ޱ��"��燊�8�lnbۏVߺ��^4�bҎw'3Ȝ�WO���G�?Lb�1�>v	�AQ.�����v˙���Z[��+xx�t�����WG����Lu[G�㼜l��%\~�Q}����p��Q���.��$i�_�5_T(�񒊅w�Y�a��(��e1�9�8%~�sN-3ch~O|���ĂR�6��s9Y��p�L�;R�.$7��`�.*���Ht����Y'.����4����L=�OWY�-1�Uy���S� R�-Ǒ����/�5wv��j��:K���)]�r�\������7�l����]4%EO�� ��.�����hh�m4�W��C��2�/��Z���>�D����F]t����M&&�et3G ��#9���7Í<}�ٷ�H��#�-,rű)~�k�u3������#L#{À���E������6N�v@�>[�<�Y�k�qm�0,~�gk�L�6A���| �I�de�E"�De�EIea�hQ�M�j�(舏 ��9��3�`�4�����P"����*��`�ܔ6@s���U�W=E
0�g����\��]�L�qQc��Wk��>��4�LgU:��i{�2h�f�(��� n��E���S <��ˬ�;����
p�fVR驷o��C������2Љ��ӴO���AM�A �z%��k/8h���<3�o�t0�9{g���G�����f�Կ{��&����~�D2�i31�����+���v5Ϡ�-(�Q�O������K���.�*R��)>S�w��>��ѵ�� �g�fO��G�
��`Րo+�ҥ�-�����\ Lh�/k��t�3���n ��[���FH�_�;x��ËӚ��rL�"5�(Ϗ�|��Ľ{���0�+T僈G������c���+`����V�ZV��*sl���k���M��$���(�����9U֟��������%#��̿���#��H2+R��*1��̟��ۯ}J��f��Y!a4��W���<ErqMIk�/����J<����(v�L���իU�dItJ�?��݅I,w�;�Xg���L�Qu '���^Z�/j���)�҆1����o�SZ8�O�u� ����Ѧ��#����/�b ��<楐x���")]��%�i5q`BnN&bB�<@VS�	鎛��csN�)ǜ̯��ʃ��*����%���{���`��*qOt.�HS����ָ.�R���
;D%��G�R�Q���KS.�-�CF�
�&X����w݃iup�����h�QC�pCm���]Z�k��v�Z���"V}���p,1I�{vN-�����nX��3̟ �kWcMR�^�5��*eb}�#��b �ޙ�
�2q���w��9�mw@�����;|��+�V���K���Hu�8V��_��ˊWQnӲ H��">f��d+�ԑ��3�;�������>|R�ξۉ�6A��rW��&l鴻}�w^�g�#Ӈ5"���J?g�m�#�d1H|�����sY�8,���69��'5�S��6�������vF���bp��1�IA�2���{Z�1#���l�֯2V�W&T ��c��2�g;�l�HJep ���(ѼУ��lV�{#x����o��VӟGH����/�}��
�B�i��7���$]��Y6FSFU���6�w���a�����
[���ߓ5��4�"|\E�����5�Ʌɢ8���;�|WK'���߉�`�[����)�}�K%��SN����ߣԬEGp��4���E��U1��ζ쫚L"w�<��
���������rW�D�v��j��H{k�/s)a��c߻؃P�y�َ�9�q`�?��
v) ��NE����e�E��3ȹF(���=6�&����Vw��m�.��{��RDԴkeX�����Q�����Ƞ�)[?�%0 i�Q�Ǻ��1�����r���@�Q��~�tXJ��i�%Gsz���^VbQs/����s\]ށb��+1^N~)��O�9�Y5� �����T��X��.���-� �&ɔ��(Vna�H�M�G�Ε֥�x��,��ZDvfX�a�r��魯��5����fR������W~ـ�[B R�*3��F������tf)�f����z��%��AykqO5UuBϙ�����(���jH+�ʥL�Ȉuȭ��h�7���@@���E��?���~ A����ܖ��ݾ�i�d�������"��7p�$�!�CV�vdU��u��K��Y&��Y|�
?��ׇ�)q潝�ӵ~��r�OL�����-l)���+���/fL�/����u�f� ��x#��V�yU��KN�(屷�n�;�t/�MU������L`�C/$�Ln>��d8νE��?��f�)bە0� 1���!�H�E�!u�l+խ�3��9o��z/˖0����'Aה�Z�ې�0��?�T�(Mvz��^���Sqm�QF��Ru�EI$�5��h�!v���k7��uK].χ{N����ٵ8�#�W�o�@�T�X�ߓղ'�\�2���~ޚ��=�>F�D��A���C*Q4ݧ�S�y0��@b������	3S�v�]�#�<l`�7L�\p7Ls�)�����=�6�Ak5v`�^��@����7h�#�����RB�qUYu{�	D����U݂v`|i��6%��N���qNp9�1�V��!+tFok����F U}āch�RG!e%py��ŋ�tq�/� �d��ي�O�4�]�����O���l}#�@�gVofcP:6�]��U�3r����;�AJr�*#ۯ�LOG_`^��cݴ�"�a˫�.�gHM\� �1	�����}�|ߣ+��X3m	r�y��b^���b������]I����M�m��P����^J���83�k��	#�?�����LS�U��8��R�t���E��h�إ���
��P�%(�B70<G;>C�Ţ���!W�1<LfJO��>� �Pw�SV*ǇRI�x����{�+��O�MT<!%y�6 �B�ҏ�`GC���>-�\b.���jC�K�Tܐ��5�[g0C�p�D�.���/�]V�>���u�S265ڝ�,>�"@�N���f��,.K��&."��Hl�����n��O��z�|`�
��4�J�f���B`����GU"0����:�OF���Di�/�ʖ�p��g��GS�Q�>�w#e<��.��v��5�pK47j^T ��0���,es�ט�h�dD���V�����W�Oӆ��P�Χn����}r�d ���b��jQ�x���?)�s|������LUya�Q&9�RX����-�ŮQ��N¶�ή9U���f����_����O]�� �*�wU6J �fX�R�7�/�v%�rB)_n�@[>}��+���s��=�/�����h�,����$\ �G��z�ǰ��#���'�_G|nZH�Wv�)��l���6�2�d!�1�w�^��,ĵ9P:\�Ń63������P_����YP r��}�Jv,�C�͏&&�x=W~u�=�g[U��Z�1*��U�yWQ�Ϙ'I�־���:��:��d`Y��FSKkO��u��j*��
�i����FA�Ȫ�|v�a�`�`�s����!��Pp-��\��{� /u���M�G�������i�\��`[�k�q|���}#��2h�ڸ?�O�*��}�/Wt���}����-O7�Ҭ��+�#�Q� ��Y�NV�\_���~Р�%+���wz��g�6o*�ޱ�%Ќ!B�7J�u�(�w&������vK����gx������(�>i�5q%O����R�M��+/v{U�[YX{�r��l�w�@���i��7�M�0-�pIb;��_/�l�l�V&� �r������5�?]U�	A��������(C��q�o`��-V����	˼���=4��K#���7uQN���߸�����N�M�u6��.�>[z�Z✷�S�����\���a�ә �>�׶�l�$���慧������8��땨x�����OK��i�Zj�������w8�ޟE�@C���M5ݎlV4<L�¼x�&��U"[P�	|�ʦ�+E?Z)�S��6,z1V�`�#à�q.Z�\��q�>d�����IL.Ajv+��!�#�-i?��R�A��~�B�i2�L}���%�!9:*�-����#qM(�B���g͢
��C�.��H�)j�$R^�xn�cc�Ӷcu�]�ƳH�=Q��KN}W��V�Ę�(:��"s��U%y�P���υ_?nCƢҞ�k��K�kk���i�C��6��l����ͻ`��C%S�t�+]��ǆ��a��)����Z�����%�{�J"���J1l)	M�� G�ۓZ!pk�L,'��.�4�P�w����5F�!��	�r6[�d���~#{#,!���f0)y�\�?��v�S���H���&"/�K�t:�A$�����,xO����r����.�n{)l�ay�m�!��I	���]tү68FzX�
��:�+���}p�g-a�G���3��d�^U!nB�� ���`�o��B��ڞȁ��K[=$˞��9
o���
�^m���33hZ�2�#�+w����7��B0�����A���'�%|��7fc��ߜ9)����x\�a1ssƕ�Щ�y������˔�B2�������R�y'bՀ.fc}�^<P� S�EB ��[�p��M���8�pl�&�ș�ئ���C��4[����zr	�`�S�ޢ޼/'f���W�:���Pqɟ��l����s��t�2&lkQ��нr)_:Xӆ��Ǯ�s�g>��֍q�����Xc�{	���On��NG	��".Zg)X#s^���Ρ��d�վ0|���8�C�3�X3��	�~.��D'��ǲ~&�C ('=�R�㡤{���_�?u��c��>|RQ��}�m�-�+�<ΌFCxUv�lm-]t7XNX���������;�q,��Ȣ���v����:S���U^;�!*y廚���Y�yp4Tb駔$ 7����)�� ɯ�����ΌO�8 �]1B?�eLEF.h��n{Ձ���h�=x'ǣ��<��Cٛ�	!���Y(�"�jѣi�8���*�xy��|	_�U�3Ƙ���W���ַ������H���"O۱F�Z~���¿�sϜ��b��Ķ��^C�M{��r�*��®��Pʘ�FxjSs�s�xYFB��s��l���}oR���;5�!s��Ӌ����PT�`���a
��m���:����;F�.�<��i�r��y��L�Oz��h\�O�QJ�����N>5`�6O5A�G��i[��St��S�Rt�6��l��D�%)Fٴ2#�#n0��d�����N�n�����i�<K܉DC���3A���}{��0�;�#,�'��ϊ�}�1��8i�)kw��UT(�� R����'ȱP��G���K���^\VQ���eE��G;�}|,�Z����q*(�YU�YOY����r����h���j��}t��I�����┿���q8q�~��" �!�a����	�	�}����rR87H�o��ϲ�Z��,!��v�Ѯ	6f�Fw:�t<F�ﹳ�E��s5ն\�=5$_�T�|+�;�6
o��g��gq_0��0*�9 S�w��U db~�JY)�L���)���'�,*(�+mpX�0���)��	���Ug�D�r��%��É�^1!��R�t:B�3cleΧ0(/T*`��=��~��n���A�l��Ґb��D�
FƞZ_��0>��V��>�fg��DJ�������@+G�o<��m`G�Dq�~`jWP7h�#m�C��
��e�+Vϔn��57��EJ��z7�W�΅��9���RM�9�7�I�v�d�G�&f25yFV��j�9���H.	��,�<
����� �Ձ/_	�E'�"�����`�v��P�k�沤�d}иm����	�$�<��NN�	oB���Xf=j$��\�qdK�݀��P�E���e7�3�3u}�X�x�xV��T*0��Q�Mvϔ{z����o������;><��H����yNDܭ�q�ĦJ�b��>�:|ΜO�[�/( ������7�}�C�3�%�+���0[I%-o|L�k���K�~F���	\9�>�mv� BZ�S�P�U�H���b}E�e}C�f���)�m��Lˆ�w���~��a�(k�1��`��:u�g�,O��w8�q�Ӈ#]��ՠ^#?��?C`2������f�Ne��J3�1qG=�̖�!��]��"��3�����~}�,"d�ծ�B?�<c�]��ۣVx��쮕��m�X���vfܾ+�e��c>5�+@�VMY�T���8;\Y�)�����-U�V�� �.Jr?��x;�B�|�I[�u��|&+,8Z�æ�.�Tg��{� ��d��FNSm�`[��Į���{�4�z1�-8�,�Ku/��Z��x������?��L��+��Ɵ�j7��nPVoP��=4a(�	����	�;qg�}-68���
	���'XĒ�)"r��m��:M��:�L`� �`�.E��.�2�o��F;�»;�S�!	���[/-�ƴ�͹ ��դ۸}����_��hx�����h˾=uj9\أ1�go������ཙ�E�G��K̴���k��a9w;��->�H��-�dLD°.`�9�L��6�"7	�u�-�f�yQ���hZ�kB���� ہ��1J |�����W+S}��)�Jh�6{kHB�$��X>�Y�HM'RZ�q���0�Z�C<C��
���~�ىm����o�%��>����(Om0���\���d�=$���w�D^��/1qD��Y��"=|�mޣ1Y$]�r��bF__;х=j;��=ʹ�R�/da2�S�������z�Sm�#aU-7���23F��' �Xؚ���9|��~��^l��sc7#�J$��	�yư�
����0�'h,���9ߊXYv�˯.���x>^u��M�l2aI3�6���N�M�|�(/1����z�������(�Z7m�s�b�AR��v���.(�� �){��HPr����v�"g��ˀ|_�
l�3^j9V�f��5�i��,	�7J�Į��3�˞ST(�=]�<X%f�D��ϵ�I^C5����e��u����g:��ǫ8Y����Ӏ
� ������%�O��ZB�nG"4g
�)��R	�ّ�)���w�JE�����N]Ƽ7�\�3?�j_�����T�� }�UQ��I;��ꇵ�x���P��~���K�q�ॄS���H���:	� �>E�f&��n*!B���s�c}��3D���z��\�W/��,&�'�v���`sX�V"6~�ڹv�:��G���q�?��l_��+�^��?
q�
��;d�j��̃��C*�aBd��O��~��k*�*/����ϣ=�k֬ܠ�G�Ι���؎N�I��cF��?d�z���ڠ�G�W���2�;��IY�����
L|��4���΍�����e5�}�л�YN���۔�Ҩ�B0�y���.�to/[���7N,�p
	��{R/����ކ��?�e�_ʊ��:>fP�.���eo���ld�J�-�D�j�� �Z|�DK�p�t�����eR�CD�]ߢ#l����z�_K�!f���`3�2�&vV���Z5F=+��(8����0��Q[�|�+����q��k+U�,�oL_�7�)�'���P�SeB��d���c?]�A�6����G���o��̺w������A��H�֌s:�Z�(�RО]Yq+-�'�d <.T\�r���{!׹��f�.��(�=t>~�#2hGa~@#�7_*��)��WMH��8aV�h���E8H�ʂ�Q����������.��?�TU%e�rY ����ȉ!����=�>��)Ű<��<p�&���A(�l�7H�`6ݑ.Ε?�a}�f��v���e41)B
�q=�YZ<B%����6���r~;}�~%]�̆��i�\f�,<��#�m盋Ľ���s��NqF��Y��&�vi�*�N?Kkv���K)��I��A[(�@���V��B�c2�`B�s���ΘV4[�7����t�J��h> 2���I�L��V�:Ga�_�)��,\ŵ!?��=I��T�Z��I%�E��}��%?�`׏AK�h�k����''��}�<ֵ�?5����?*�����7a��ӫ�ć�M7��'� e]��7��)_UDP�Z|�|���-.��f@���Y���(�=K�:�q�c���ZF�[.�&���V��o�z���L���}���C_�6��|Ʈ{�ru	��f�9q��ja�v�����0~*�&+͌�WڿWϢ�Բ�7�~�GDy�9a
x$��g-c�ձ'�F{C^:R��>�O�w,�ɪ3�Snϴ�K������n;  u%?a��R��@ÊD1�1�T �&���}���E5ޟ�"�r	�����K4��,�mN����li�!��/0\pәb�I.�ؤr�ى4�?�&���������FPER�RuP�Y�K �nSF&���L�o�#N/�3�]����=�(��5��	��}W�C�}J���f���dCP�5�ȁ< 5~IC u�nzsF�Q����1��U�O��=l3�d�h05���=� ��w�L�Ҹ[�(i��JzU<S�7 L8.mxo�GP�����`��;Ŧu߫�s�j��Q��V2C�+�Q�-[(�ZoN����
���߶��!)�wq���_���{JG6; ���ڱ����L���ͿA�꤁jr���n��آi *4�c�o���u������jo�Y��^̸�[e)�>u��<���&���Sp*V�+�HtX��������\��
�.�<���.�]+H%v�����w��X ��W�5�������}k� *�
����u��b*WEsl�D@^$�W���(���Jݞ�w@<1� ��:�Bh���&<������T,���YN���Okhp����_�����׫���w�w��W]�$����?��>����v�\U�l,�ʔ����ڲY���4P ���0 nl��c�$�%N�d�`yC�$�@���-Vw>������s}#nC�h�Mb�M�p�H�w����5��B*�
�ȏ�T�ɀ:�`�h������p����=g�&��9��R����57V�&�v�kC�ܿ�T��(]}���g�<�����'�ϺTV�=,��#�y�1�v������l
�$�Y��	��BF1��R���j�#<��9��g��v_5�l���'A.;����p;����kc��b,[HT~����J���y����HJ����?�/�E��n~�(lљE����q>�݌F��n2�:Ĳ��V�������T�:V��ݍ�o���~�Q-���B��r}���I����\�xu�w�w�Q���-c�tA��$�Ҽ3��g�25�V�B��Ə{
�\��E8��+���K��`lS%�C�������?��t
�=�r��1���V��c Un��`����Ƽ��^���M�Ua��ؒ�՘���1Ȳ״$B�E�;���S%����OR���\#�:Ţ\]��N\�3� ?S
��#�d���Rs'>(�l_R�'F:�_� ��@4��H5��V�]��ZSit����`��9�*qn��S�`���6����f�
�F52�;�o3
<��9�k�)������>U��n�G�]�LXƻHd�P m�D`������B��2��W�Asѣ�
sTKR�פxf�,o/�:[��}r-9�1�pv�!W���k��BS�9�R�%6���H�8{�ؕX�X'�f�m��P<JMo�f�w2�8.V'���	�Kg������i^�80��S��C��l���fO��sOƇ}��ъ.����,���Z #�tL�5e�'̐2�V��]k����e�l�����J�WQ�i �C��z���J�j� _�,cV��_*�UuK���,cDh][Xe.��.����\�/]������-8�������";��vYBM��2�m�	�r"cTΆ� '|�����f:���eo�ha[�6����eS��ϒ�(���6�f�Y��S���'�U����P��4
��>�/�
�̳��nʨl�ָ�̺�	\:8ĥd�p��d�#ha�:��8M΋�Н��>ϴ�*P�V,)��}�a�<�xM"�'���X�-ݣN�j0��@�S5�� �aF?,!&�Y՞��7�a��|�ܛ���J�%�:������kS�^t4���ȸ��;���V�����"<\u �Geq��J4���b���^��+zA�҆rtq�0�`:��1&K"�h�66��<�m�TnhI�>.�,�l���牔P���}�@��/$����'��^�.��E2�]�f�Y �?mݓtCڼb��F��E]�k\q���r��,3���L8�!!����L��+:����9[� �%� :�?
�-��	dBk{O�[!���wk���n?Z=N���ɺa#���$���/��Ξ��3�������NA� �d��|�J����[Hw���w��9��G���Q�u�BC2�"I-~�[�@��rLJ�An��[���?����W��YǕQ*r뒗,�7��6[(�+b�oi^�^0��Q:�K@v����o��^{cX���q��h�_w�P�Q3?��~�3X��������E�&��=���IqɄ�=mB"� *;k������{}E �����0 H�E�XZ�	[��#��s	dBc�~9��^�߹����������CR6�p෍>Y�)WSL�u��~eCi L=�k;�k$t�$C��A����E";��6��W��J-�SfW���op7$�
qQ;Y�{A�t]D�b2�h+A(A+���h�k��}J���/�}���0/}�X����>�r��i�CH*}�FΡVt�ۯJ�pҿ��պ�����ο�yp|�.������:=�T< �E�D}���D����L G�l�D]�]\�����ĮZ4[X��T	�?�������VC���j�a�ԫ&&�.�u9:K����.�����=�'h�x��E���Ofp�d����MP"�*�U^֭R�*��o�	�@�w�$�W��A�gj=�Hǰؑ3��@�ϫus�������3TnT���j�]��e�x��8��G��Y��i�[-h/ -Dn�h"�*%/��x�&lk7�c����c���Dپ(l#���6ɫ�#jbNưX:���/�������ř�G�I���n=t^�z*[[[�}ԙ�����&�Z���N+K�<��O� ���c��+��� ��?�q�����e�W�� ��zR2
�%'���&�~o���7d�{-�zn�uͦ��Z�H�c��.�Rr�RXqC��Aij�����ܦo�~[g�H-��/$������o���s[a���T�v�o���a	�V!B�ҍ>Jt����6�����2N�d>�Q�V�L����/O�Q�Ҋ�{W^�ArH| e'�gh]��������Бj���Lu�y������Rѧ�[I�?�#u�E/�\��G�wct\�x�;M���Mu�W[���&t?�#7�j�D�x����{��UΆ�ȹG2#��p���1�6��44u9c��"�@:��M�޻S���;�]��S�'�1m�06[M��G�	���ܜ����^#l�f���	%!�^J��_����gU&$l$�g@x~�{������}��J���0�
t�}�
��,tX{03�m����3[2�$�B?c]"�ݞa�m��/}�1?3z�2&Q������As�ץ+,�!���b�N��4y�����yRX$F��@�7�0�cq0�N����B?���( ���;T�j��Fj2�2���J�iŻc�HB�:J�1t����ك���yjDOY�?�ŧ5�p�������n��|Ζ����m�*�l�t4g)^l�"u�-o���0���=�Ь����%�^��C ��Q����벪(ln������m�D9@y��`v�*��z�'��t�S�X�)�f	��7� ���l� �Z�]cۑM7�r�#��CpL���%��vn6=�^awC_d����܅�P��%�x�5m�C#�'<�͝b����pq�]�����k%}��
O���`��1��o3�\\�Ț�TBR��^��|;l0��)��r>k�nlbe����$�# ^Q�
������u}1�^��7�`P��Ne��������5Lƃ��#m�b�-���IW"�a!O�nI�4������VW;Ķ���F�Xc����oo�˄����u��HHl�Ɉ�ͣڦH��o��m������HQ�#�UЙ��[�Jq�d%�]���i��b���T�
��c��O��3?՟���RPY�R"ڎ�=%��o���p�iJz:�X��_�v)%�\qnE��n���(N�^�.{���{�(z�z���m�_�U�7�/���k	���0�.�ɞ����ʂg�Gǿv"R���vk��nK�����FV�&wdtx������@��������N6���{f
���{)9eӄ�f� 
a&�E�~��-=f�Dj�7���;3������Y0S��؎�*�Д���4����5?2ч�y	�����s�l��8t��Y�+6+��V�K�'2���D>~r�j���1�%>qȆ����O��z�oX���E~"",�sA��~�Ad�߭b�����ճ&F���~����5#$���1Z����8�='��`��3���n�'��99l�a���[�(��ߚ�'s�[�.���f{z�yf*i�z޼�Da����X�[�^�)9�`g�j��}k���|-��	u�$�UI��Г�GN�9��f�w����C�E@����4�s#���;CN�QM0��A��'�ᵑ��/S������uĥ�4	�u䘻MtTo3|3��p�����O:�Ɛ��W�P�"�m���L�0��?��D֒��u&f����Q���E)4]o��x�Qo!���F��7+�Bn
�����:k��5�%�ӣ��vh	m�}�<�P��S ��|��(h���IM���%)��8��SC��� B�$f��Q���ҭ�ze��ū7lw�ޖ�����5�9ox���0���W��b��SZ�y�a��&�����$mg/jF�k��Dw[���j�^��m�\cTB�</�U�j��<���C�Q�V�*Y ��3ڗ�V��ϡ6t��\3�FZlv�_�h�BhGF#e��M^��%��QPaY�VfȤ����7v��p����^O��%�IH��-�������舀��,e�sˆ3fa'���r�[l�&��9�����;^ЎA�,	��xǩ��*���v:[�NVIfz�hz�y�bL&���-��^�3Ʊ�&��Gqj�V���tT%��5M����]�t[{�cSn�{�O��ꊙ�)�坐���$�4{�JL��dח�ݹf�IJ�Th�sR0�6Q�-0�ӕV	���&�� �|A��Eh�vL+]8����jJᚭ�0�Bp����Bo~��l�*�XJ�p�fORnC�\p�([d�}ܰ��Iͽ/~sˈ�z�I\�֖��洫H>�M�I��^�U<2�Q0�h�w�>��)Z��͖�y��E�8��|8����x�r���ų�*��`!��2
��f#�E��ac�陎-5�fc��[�&�1��:�.�	ڿ�:S��f�������Ghg�
9�Ё�b��u��C2�m�h���e��>�� 9��Ӫ��}&s�Ē�\(�k�nU}>�7�7)?�Xl�h�7@�Y���^��T]��_!v'k�퀄�ob���g:��I��r�)����j�GH���0�c���p����C�5��s?%�	Ǩ��` 묫#��'��_��27�@K�|�O�	��0�YT�H�k���}���M5��Ve�7F�۸;�g�%��o��0%_T�6/�JB?kkl���:������	���`��RU�!�����E?��D���.�F���Y�-���Drc������{��%繹pӅӷ�6�([��.�UA>����㍄$���7���}�>c��3J���[v��,`rߌQo��9�H�~�z���g�f�c0�H��ƽ�jֻCz�����ߢ��L�	�Ȭ�X�Zz��ـh*�sn��DS7$c���%F�6˳�A�r�o�B��5�	��Eǽ�[N�s�J^|逮d���lH��qQ���!M���%��Qڵ��cY/P9���sW�xk1h�Tf�U։��~f҂H�cX7}�q��T��FP�&� 5jp;qf���k�Kօ :����}�B�2+PU�0��6E��x;��Z	���{���e�;�f�vm{k�?����y�I�E� �e?6�g�����).7�u���F�w{�A���L�ȆA.�x�~P_���W#��nUw���s�i�6�MD���#���bbr�M�ˬrN����ZT�[$�Qv�H�;߆�ZC�pd-�q5U�FN���	9��G�l(��g����YbDa�޴x|=&�Q�,����x�9�[��3�W]"�M+��D�~�UJ.��&:���%���i6&p���Yp�P��$ཟ���L��5�A~/;m���_��]�I�#7	���bB�ϓO���~������CX��e�l���!�	@yP&d��r�����U/�Vl�82���q��,�;轉�����
pѻ�n���K����>P&y޲Z��������t�(�uVɨ��F:��r�a�^�u��4��Z�E(0Ja	��c]�[zĴa��A�0;��e�e�b��;KG�	��f�~��ዹz��m�M�ٳ�T�9���]=�'��#8�%OB#�O'��G������C��dpy��;<��&�4w��\��0͐5Av���r�jY�Ő�𨒰�O�?���-D�����$ˇ,!�5�1���Z=Wr��e�ĜQ�=��I��e
{�u�)��� �o4(h�u#���ج���H�\����T>�oh�*2��ʙ1BQ�����+�jɵv�v�P�w�,�P��4Oaw�;U�wq�[�e�]%r|r��ِRb�e����(���/**�����%�4򌒮<y���3�)k���uR��Z �v��3��59�h�,_x�%4z�ٌ+����o�,B$�� ���"��U�/Կ���ԥr��;�<�K��{��x���O�2?��gXK��MZ� o��
�M܄d���8q������/v�ˡ%�ܴ�@���~=��*(���e�/��1������˱O�(C:������.Wq'�DF���d�C�x�ň
J��͟���:,��(�o�
���ET�Fi��W�1��t��I���V��k/����D�t���= ��gGDØɺ/dv�9J(��۪h��'����C�r�켹t�����ܬ�a��� [�nД]?#�vڋ;�9E���2� ��{M`���6�Bnk���s���5�� c��0B���DO枿�H�%0�/e��1�p
5�~�����Ys��B��gK�.�0������^�k�i�K�[�yְVd�I����tCI�E�{*�oθ��e�k�7�
�Ծ��e�wʫ���,����v�d�FTL�3��2��L����U���}��h]+����<����Ґ���� ;t�@��[�U���M9�E/����>߲�?� ��i��ɰ�* n�d-]��]�~l�9��Ҫ�1ϔa-Xń�K�w�a Q	��F���1)ui��
[�c��C<}[Qx�&�T�,�
���Ҷ�BW�O(ؼ�a���H"Fs4�t���g^i�(�c�E��.�{�9�	@����xDZ�HL�Q�ݬ���.�z�0���p㐧�6�Z��T š�U���h��7�^b}(|%&(��u�9��e&z�+�G/��i�w�P��� j%�7�ZT��AN������l�U��I�4���v�M�R ��<�|;�<Y����HE�
�"UΣ,��K��W���Al�d�J}�^�v}�v'n����]$9�U�.���GS�p{ ���� �6�K�)�p��D%P���s��}�z=v�F�'��zP�X��6-�������p��A����׻޽E��i\��;>R�.!�əv�=�Š+Q�r��ө����Ǚ�].U;����/�֝��DB]�5�D�(�)�Q���?d��r���]2�̋��)v���1��Q�(U�@<RuG5p�� �F �s5�����u�=%$���SY	ʆ$�r^@1E�P�_�������bKH)7��~�X�E���y6r�����nM��3��T�M��\V�H��Y�Z���'P2s�?TU��ܳ��{
�e�ʼ�%
s��Z�Km�ȗm$���d���i�(5ϧ�s8�K5�u^9%��6�J�뫷?���wqh2�Z��d6o�h�Z���H�~��U/��r� ��挛��39�>4N\Ó����M���w�ѳq��j�K�ssj����,p�� mc���X���HB�����h�~�
��1��%�O����Wkv�0�� (_L� '��k���[Ó�v��o]�Հ\���R��p|tn��첬��WaG�iJ�E�W��� ������.�.5q(���,��]����������g�F_��Gf��\Z���-�`�e�I��%��;Y�Փ��i?�3�X�6�he��9�����X�o2$���XRC����}K�۔��|@�x����2��ť�j�{��˕Ҋ��H���!w&�U��AKԮ%�\�M�����������2]Ʊ��#��ڦx#Z�����3��6�R[x@�|��s����j��8G3��)�9���x:��|���=Z���6��=��m��)�Vo�Ǻ|������!E3�Y���wԲO���89+��}|��dw^��'b�v#_���)�aN8�!+�ܣ����L!����ǰ�;C�׌���[�Ϧ�?xVb�OM�@/*�P�����
l�C����
�,Sjp�t�����m4�]GnQ7n��DWk㜲{�:-��F����{a`����ן~5`f������č��I{��"\�qiIS~!�XI��(������kppY�2(�{p���ҁ��b��K�uk��|[��� {���y�7\&P��j�go�}� ���^`u�85A�4G������o��Y��'�e]ѩ�Q�(&�+e��V1[CTD==���LȒ?���|#��
AI?73�rfam2ԭ�ͧ�d_�N�F�l	5UMV��(S�L�0a��vmWo�g_\�����,�S�~�xȊP����K���Ȯ���a��ņO�c������n�-�_Bs���$�j���g��i�쿤��P��*�q���[�J���ܠU�CX::��[t����{{t�����۫:k��P�z���\�{(�¢II��ڢʈ��_R�0&�p`�����ԧ�4NX�jgWIz^��jy�^��Q���C����ג!Z��$0T�ٔ��-Wg�$N.�n��|U�"����A%C�"�<�s	w7u�����lE܂}<���M:nD�9�0��􀩂,g[Ο�V{!�,R>�i@O#|k����us�Xdb 5:��˧����C�%a�K�d'j��Ҟ���:?�ޱ9xAb�����N�˱L{�YUON����m��ܠ8�.�N*D�X@�)��s/<|�LD%�aA�t�j���%Ciٷ�i�Sj�՟�CQ���l��A\�uX�Qưp7ێ(:��E��ˉQ)ٹ��cH�I����G&g��V�{4�v��̥oh��wI�`���@r�6�ò�г���?
� T�Y���TE��ɻu�+�G��v �e2;��?EO<s�F���� _��';J;�RU�����:fS�T�tID���82b
:'D2^�s6�
���Y�(|x�T�&�h;6��o~h���õ�q�m2�Q����ܿ��'�yLWr@��=A?,_&��>�=��8+}]�z-�@�A��4��t�\{/J���y��j\R�i��>�U��E.�G�.���M����q��F�ly:^�z�_]�a��&�K��K�2l�,��ɿ�FGtP�G@�m����ՙ賍��kuN:Y!b;�j�7���(��˽k^�։P�WM����!H6�4'��_��4C�����Ա ���8����N{z��l���O�V��ǜ��D�YL6�T�w������l1�� �˱sZŒ��f��ħ�#H�鞎�_i��D�v��"�Z��X�hrUFa:tAt�N�L��o�>�+*`�C� ��0Fkb穚�?��[ɱ���Ȅ��?X��$_�v�Bsb�j�LA�g��^%ȵ�3j�:��d�̋����7VS�w�� �ה-���V�rG��`;��H��F/,5��^e�7\����fB��o�?)��-l�����%�	x�d+��E����`�5����X�+���7���t���2�����s��{8d*X�1Rq����� ���	�7=�	���
?��Up��I�����;��K"����{�����C#�\|�+�fN��p3n���K��eqk0�w� �:��c">w�G�y��Ps�C�[��/�
�8�?���� ބ)izϠ6����"�I��$����f=Gw��OIE�Y�,K��^*F0�ש�*��؈#��\K)�ݯbB�[��fx6</m2f��A�igT	|��3;؅�{��G���̍ΰ��
]��6Ч�Z=B譂�E#1��^K:�E����IZJ�,���+��Ɋ[$07l� X?�إ;.S#K(\kU�v��[Ks,�FQut��V��*/����jsP=f�7�K)���^�\��:��e��J��	ꃜ�k_���p�o�e8�WY��%��w���+4UY��M�k�|�0a��)�$�FmM93��{�p#��"Ug/�Cv��+�x�9U!��N����O�h�n��9�4ض� 'u�V4�p�,��樛+����1�P�[|G�~TF��+x"��U�D�2�*��Ɍ�%�`WV!�aߖْD�28����^�Z0���_�u׋�]�=��M"v4�q$���Nm
U<��,:��kV �����ܪ��+�2�/Łi���j�Ы.T����_��ֻ-�^�G8I=��Td'̪1�]�I�w�^�Y���-+��o�9)���P�H����Z��(쪛gf F����{��e���K<~ �A�����ȫ.$H�zS��.A·8O���|K�l;�l�f0g!Cz��n���}��JU��1N�j}��r�T�0-��9<-��/W��1�
�ަ�&��O��.��a����֟�U����+��s�fs�f>}_�*��?�5dd���_������b�w׆����YϱV���dnu��
��ڷ���TCD��b9�GY��K���J{����H֡�XE0hLΰ^�a�Ս�xj�]�B�EV���  wHd0�1��%&�JUd�T�7��"]@�!nE�	�cV��1\a�?m�'�P�9�f?&�� 5��z�-O��{a��Α�%ib���ğ�:{#�{Mf��-��»IϿ繐wW�2/�1����kţ��7�/��7�9���Lڔ=�fa�&L��6n�j��5��d.Ŀ-
5{��=?=A��c�'�5/
��yΘ�]�xp;���*#
B8���Tw�MIv���;�4E���f>��T�o�_�	�&��K��*GANM�U�� ��ѧ5��I�ɶjRh�j�}֒2��|-�c��_��W���!l�^Y6$z��s�~7s^�55B6�֠@g�\G���Dq,�{;�m{�F�\e��Er-�-�s���yԧ'�y=���h=��AʲH@��:����.������X��tH�o�,������^u�� 'rW��f�c(���4�QQo8�"�j�ڲ��"��+1���`���D�#����jj*�Bǵ��]�"~=?s�����J�x3�j���*Tt�"�q_�#���*B"5ɽm�`�&�����5ME��ӅM�������/Tb<B@��XQc�IĊm�{�?�w�t�,ߜź��y���a���A�C�QJDk�*�U���6e�mT�u�(�.����<r74���0�"��G��A��%:N=��|@�b-4�IF7'�O�R�	�+�= K���:uM]@�y�ü0zX=�Ƣ'�wz"G�H�1,��v5.�!��C�M�>�6�|oŤ$�j�ŘTֱ5m�S�B��:hi79aW��,fQ�(�tͥ���c���1�Qn��I���:���բ׃p<r� Ј�i%R?�O:��9��XjWG>�@���f�V���H�֧n���0@'�K��@�j��̔����x�78�V�+w��Bڣ�<����W�h�E4 ��}:�7?��N��r��)�N}۞h��IIL�`�w Fl�����V��;�p�\#|~�]�bG!Lуtzո�y�c^>���J��/�ӥT���4�WN�Bá*�i �ED�q"���+c�4�� r�a�����p��k1��`�a��{J5��R6o�.8tB9��ޱ?��F��c�)<��a{��	�-��)Zb�"�:�C�=7_���lx�&0�@�������*��n
���v#)!9�z�ր�F���%�d�#� ���"ѡ*T�WK�t�N��^R��?��XI2F0a<�g���kN�$�cO�@�����r��R��ӳ�z>�TW ����fS[����)S���رn}�~,�s
�3,5kuFb��9F� !�d�(��#�E�mhB��c8�f��
�F��l�)D\���9�6�G�8��+��]'T��WF�7��EWb�I}�G}���K$���J.��J�	\hxش]��k��}4�|�ӿ�= ����x`X�f�#)���<$�oT��zO���?�?��B��Ù�" wlA���8�jl0�`���E��=�=~  @-I����M�b5k�=�c9�ۿ��������&�9�V׬��n�j̍��]�[��g׆Ǜ�^B�6�0N�L�Ȭg��E�0AI8j���r�S��\�_C�;u�۳�㔅�	ƒ+	$�_�q|�.�$	
�풤ç���Dx&lS�^��h	�8��qOCk�R���g��A,+=�����[
¾O��)C�$�5�g�a* �=�=��|�(ƸV��q|C��BF3��,j"�*�%��V���g��m.ew�ˬ��I�l	Me[%ބ`�u���t�Z1�x'.c�%M���o_��y��h)<�@o��Ʌr����el�O��M#�viH��MΔ�~���%�^g:N"!	}Z�d�O&��N�lvK�S�7��,���'�o��yf���U�]�P�?�7�th ��)'>�I�@R�]�3�\}�I���ѳ:�)�@��7x����'�$�C�K+���>�4;�^�1��m�2]�4{w�����g����D�K8F���3���-A	z��1�kc�hefN�#�k}����!ؽ�Pp!��MU[�WY{���rc)�6���fe��?��Xs�Yڻ'��,=Ȟ��$6��2SX���}f�n��t�Q�ٜ$���&�>��Ww_�.�+�D��s.��@Z#K'���1�l:�D�lݒ����2�^Q�/b�\�����r���BZ���D �Ƞ�D0ND$��Օ��tש撠�)X���S3�1���%�H���+I^�N<���6G���������ߨA��"v���r�p�K��A_R)��uLQ�sμ_b��#�;˖r=�B����~c?*��mV��{���DШ�j�I����Z����J�f���V���R�o��~�K8�@����>��:������=��y;��x�~RG��t��	�W��������R�����]:��S(]��E|J�rgu!_�#�����pH�;ʸ��|�#&d�6G� }��(�=,�$���`�;�Y�̬�^� ��B/��Pi�I�i�Bk'1D��cHY��`-�lU�J���]XanH�߽��G�B���N:aIi�t�G9A]�+`2�Tr�yt�!��$C��:�I�v�6��ݮ`IOB�Ni�Q Ij!�r{rD�� �ۼ�&�VԨQO��<���v�O'�%Ͱ�4�� ���A�XN:���j|�0�pm6�v���Mh�"����4�`�e��j��-�#�`?�&nRÍe">yv���}���[�S�������h��e����$�{e���I�d��]܏%Ū�t0y�T�Re��Z�i�+�MqH2�w3��);:�Ԉ��5�P�JR�0�i�P������Q�>���bg�t�����4��~;��@��(�6�g`�����-E��ю긄�.�ﭲ�b��A��!��J��lVُ@����FÐZu��D�()�k��1�r�V��ɓӌӾ�_3&t�c��~V����JZ��Il�Zu]�R��6)��M7���ȍ>fe��"'�̺V@�x���") ���<�����!,w��p�%GL���k~�5\�f�I��"������Ш���@:���5�g洰!�V�蓧�>�t������ ����l3)�b��?fT1F�5����$�	S�l��#ֳ�?`1�,��<a��*��t�6�vR�v����`���$S��Z��~���0"��PFg�%���ɡ14HM�ڧR����K��O��\5ۤ��Kg�����y�d��X��dl"#s51��I��,ލ�*�n�������fg�6�� �[���i�b,i�)b�.�;�=d�D��g!F���M�1�{��@��G�a{y�J�F��h����l1�_���|p�l���?u|��R�N�ͻ�dt�0�` ���%i���ә��n)�'�S!LF���9��H&E��§o,��!F�z-.�6�;��AJ�9��	���'w���G�����E�P�T�qo���h�:!0R�YCAxP����~(����ӓeOj����7��َ��n����6_bY!!���USmf�i}�4G���*������hQ8��g�Hg11�u8@�UԕQQ��N�L��키�ZP��I�m�:����`��Q`\����?$�1;�C&��E��mZ��o�=��H���xų&3_�jJ2�^@�t�(��x2�g�{���i���j�I�.�|$�Q�U�CHy�{�ʻ�-< �_	�Ho��<�j�㣓'pݵ�"N��{� �_������_,�!Q�c"���qϧ�8D��7b������Z�gߎKIa~�7F��<����������x���8\|q��!m4e�N�y��U[��T=ύN�|����!� ��}���b�AK��-V2}�9��y�74�Z&��qc���mP��h�L� ���+z�"��0uY�x��dL�L/��n��y�J)�,�Zi����.����F�{��8C��A����������&�c�}�˖pZ��KD��/�;',��ј0�	��"� ��$�&�j�(����R\a�����(ߢ�{��p�˗�T�F�I�IVH*�A��Y�K�d�����vK�b�-epO$�]�$��8�Ct?kx4��LQо���ܘB�Y�sV�V��L�C40���qp���S�}��K�q|����Aqܲi!��B�
t�}����D[��K���!h����,J���T����^�ɨ^ײi��o~E�MeӞc��-��脶�MG�x׀+�G{G�%�~!Ւh���c\���qS�y���K;i��;;�T��,oɺ^����]|V�:B?Ӻ�
~��ݫ�&��N]�xz�^:JSL/�Q�hf�Ł�-e��1v�pxc������<.��j1����hH�j�����"��ТX�w��@�A��W�@%K�4�t-�]����RV�!C�����)�逮J���M���=�F�A�*��TI�xT��n����H�|%�.Qi�Ш	
ǄeABqB�3�oY>|�����ΐUu��'���
))谗Q	�0�-�����^���+ݧ�Ρ�HOne O�8f�<@����*ú�X�+)���������U�c�o�E�^�ƛd������������4 A|��X3�3��UE�s�����9��[�����jQC��${��y.���Q����h�3h��:6M0�����C��W�����F�����\�Z�G����~�v��Ů�%��nY`kL�u�6e]��J���ۜ�O�	�:H�U{�+;��G?�*Ӿ���׃W�Z^8����2�}���[:d�(S���ZB�:�YnΘ�v(��[mN1����Sl����g��u���IJjt"��Q�Ti���2�X?=�J��eA��&��_�E���I�Wf�e
�8�׈�E��3=9gR�6�P����EU�_ư���8��j�d�{s�/�܍(���;2�ޭ{��O_)�(��p��m�	c�>�V�*��3��tR@��h�����:|@'<o �t��Tت�Y�v|E�#ߥ��C3Ⱦ�X4x)E�E�R�e?g�q�6���ٗ�%�<eOi4��r��J|�Zw�B ��sO t��P^-믆�T������_B`l�4W�RuAC5�8).���� �6,;_��?���?e���b�ɀ���O~�����'�	'�A�m�3��!��5�,�G�G�ict1�t蹃�{-*Y��5�t�[F]/�+�?Wmw�j��~o�f|M�Ż�[�͖��`6�<�t��]>V/^d&���ڭ'��ρ��D��M&1���J�$�\Mm8�T���Z?R��s�
zĮ���k�lR@�t��;f��#���رՍ���tإ|k ��.�=D�#}2$0�3M�0�~�/��^�'(h-̰8jVs����R���G`��TsɊp�qc2�X��^���<����k�+��8��xo��_0����i�dH�&L����'�����JR��K{�!�ς|�FbC|η+e��pUi���'��\���{�X��M���`�$��Q�m[��EU��y饵�Cj��it�{�����J�#Q��l������tb��@h�v{l0t#ۭ]�Nk��h�0�3e����A��2�q�~��4����T����� ����o���8���ї�L�|��������}$WWr� 8/���B51�ؖ_A�&d��W�PxAL��+zwoZ����ovo��G�0�Nt/Q�� �5�����sPh���j�k wt2�i��X7wS�}�?�� YkI��b�~͜�o�r����,�J=��d�vj�P�H)�g&J�L�=�4�a�zIme�E�$#���

A$#���n��#�@;V���\�}EF��x3!�4`��J�YZ�����!Gb;W�,8/w��>NBE^	��<,�q�FV)w�a�R%��m��+�Ӫ�˽��M&��q�-P�{�+$R'|ʥ>}�Cs���T}��-?w~�4A�ϴ��.��,C"3ڮg��1Q��c��l���
-����~�x/������({�-�Y�>��~�d� q����@B�iv�N�4�vӸTbF+��D�n�u��7�(�ע�{r��*�9v���p��[!Q�N����Ftf�g|N*��f㝩�:S�q�L��_߱����Ԫ�	E���f#\G��\Hy=���xd�����n!
E�cM�7�׫���Bj���"��n����M�ce�����ݪ�Px� �oy���{Z�f��������d~�����i���9�vCr�W�QH7#����G� ء�T��c����7)���<L+�}����>��]O�'}����[��	�Zn����[��,�o2�'�M�$���oFmyp��J�n0\�3�`@�٭ʡa4�fX���^1.�ӏ���!�Ǧ	 �Ԥ.:�y�ƶAX�r4�:��iΰb`���05TBqzu�2X�2Dԥ�r穋����B2�>�7�{*�����!��ח5���K�3^GG� �X�5o@+�;f2Pf ��MM"Ɛ��E�t�
�KUh�Փ|�����-��[$y��1�C�9n�����`0ǽ��z�&K�g���6�J0V��x�L��>y���s/�
 ݦ��׹�C���e늓���9�Ёpv�G��Ǵ⸳����5B�����ur���-Z7�0�%��G��^1�	��em��ϗ|�������=cre���Fd�1\�\����m0~+"���#_1�Q����.�A������#�Zw�F��dWC��a��/2����E����mb#e�������\' �zT'��z�[�Sͬ>H�V�{y/϶�܋��*M�N��?��f���N�R���$^_l��P{�Sn��Õ�xnLvJ��a���M��uee�f���k�����v�CT���V�>=���o�zU��)E�g1,M�k��"b_�`:!�8�k�5u��9�k��0��� �\9���,���8#�=-��ͻ�����+!.rXdAL"i=s׬�2�=C6�-8'�w��yi���Hd�p��h���mȬC�,��e�H���ǧ��B|ZW����a5BGL��'�[Q_N��V����D��?Wqd�I]�/��y˅b"����49ۺ*�E&Kwꎐ�w�^�1u�oZ���d�����5�n0o�Uw�c��(?h�g�Rbv�dR���8�������ޛ�.�����)�Hw�bw~0�MBM�g*z�.T�)�8"Eɗ+�w	�;�ӿ�Ʀ�#F���r��:�ͷ�̽�ny��Tf7��n|�L���yT�[%���=FX2��2S�#t�*j!��w�39�C�sq�
�lXc��!�6�u�����6��)�@��1�6��F���xB�W$��l+���I��id��Y�b�Ɓ{�B`E�b��v�$�7�,�|Ӄ���0�P��F���nI���? ���o%~a�0K2��И�k�q���2���u�;$�~�j�Y<��T�7��=�C� �	�&�D?�*|�|<(�>sɁ+¥�U�����u���Z,��a�����9RDV-�rۖ��-s&�7�Nd�I��K���#�0˯:�̨X�����pX�To��O�v.3�|,��[GR�f�U}�,��*��8(��q�&��C�-�H8��:��ͩ@Ա�7uQw@h�ǵ�Qo��)��I>fI�_�*�Pf�5�s�x�vv���i��&������T�����|OD̙�����&"<����@�O�W�˸a�����XxQ�'������KO2C�wH��KŬ"P��1Ȧјg��"@�?��/3�h���5�m�FY�骽�(:+@owI|�I���a�a�(^#l�N)�1n�G����Z���&�S�MEz�.ؽ�U����_�3�*BE��m~�R}Z�rj��~n�δ'86O��<��m�a�^,�d�9]�JL�1o6��t����
6L,g�E���]+�ʨ����I���BcҌ�A:2����1uV��q;��8G�W���{厃ǟ` <ЗzCz<����^ʨb?���U���F�4�SJr�$��s�
������[�v�\��ez��GGF����Pao���Me��g�Bs���坟��U�>0_a��PՅ��뽒e.��H}�R*+N"(��]r}2U�);�Ak���{IVٓ�W�o�cv�ڎ�j�� ��m8�h����%����b*���)��X7	#�X�^+K;�����||y�
?KdB0n�I�Ns2(�	9��Ǫ��q&'{�=����x�Es�i��g���b�٬��
������}a�_
U����Ƕ�(�o>�$qib�MD��˕i{}��Ҭ�\��g��]��j�(0�nH�f���G��&����5����wt�C���P�9�L�roڑ%�����I�5Q���IJ-���:�0y�J讨sEs���0!~�\����|�5/�{y�
Q�Bӧ��B$�nѤ+���1�[��BK�����~]bi��a3�����f8�S��5��W��/�d=�=�g�4z�g�f�0u}�	��q�W�����*>��[������G5��b��6�Vȟ�́���) �X tl��n�o�E�ޓ�G	����9"�.I`�
Y0<s��U�$�e׍����"L�GӅ���5�4�}㒼�p �|W��\�7�w̨��a��Z#m����Hc�2����P�'[>��oC,[�	���|4�Ӯ�0kt���}5���}��p���y�u�K�|��h"��N2!_@v�X�փ��d����}h����-Q�*7{���<F��ȃMq«?^�n�6��͗����0޼�l}a�Chy��]�kHN_W���Y��3�&76W�(me�fEՎ�������.*� 7� $�����H�L斿�h�"T�٨hC�:����� D`���S
��G�&���
�j8	
x?,���#P���Q�[�*�hA'ۼ����BD�th3�Y%U�-;um\ 
qnV��N��Y����Thd��8R �A1�AKf>Mn`5g`��Uj��]@�sͤ��ܴpI^����Ϩ3��皜��'�����,�<3)W�kŧ���рD��e]�h�ʚL8�CD�e��xoh��,J��͓��SJz�7�YQ[�������.�\gduӘ�JFC���c	�Ey_2�0���ʔ�z}3�Km�Tz?\�bT5}��&j�m����#}H����U���ٞ:f�_ٖSa'E�v� ۭ/�X
%��X���j�d���5�Z?�!�<�D��ʃTgN���Ģ��r`�m����s]��KN�\�-U��^���r�y��:���0\"��~\a`�e�*���j�<���zUz�]�@�{���������"�d�<�@�*jq�&W�0^Y6O��I�O��S�lg�{-d���"*���54Q*�>�jT���u�n��x�zF.n(\���Iڗ�n�¿"y I��`�Q�Q�AXb�j��O�JS��@�ѝ%�+=�@��(��7��"�un6��V�d�s4�3��o�E���ş�U=�yP�
�z���.��yjp1���X�G�u��u��ϩb�o�h��GLi���٥�1:��I����A�V|�#�A6�^p��<4�a�L�7?f;6*�h�m)��b��8a�b)0u@k�|�f������%�=��(8����E��~���`ejvT�����u����N�4�������14@R}r"-�^(���EX����^g�n�/`��J�T��݃�	q�rZ6.�a��e�F)�mوѡL�J*
_��ZXg�iᩬ>�4v� `��|-����ېo�*�)�Nj�v�<���,�[^��Β�~�Ic��~qb�N�V��'?�U�:��$%�Wa@UR8	�&ڣ�;�v\���Գ���{b����S�A��C��+��*tIZ���DfN.	�xXaϰ](�/j�	��v������JR��l ��o��
�	�C��TK��Y�k�l�ۮ�����(�s���Ѐ�p?�D�>��AK�)�
�4���b3H���4��a���7';����?�&nv��߹����ϲ�q{-�Z���C��_
 <n�/1�vvG�`���V⌁i�]�����%�i�"�*S��=7�<�/�֩�u!��w�)��*�z/�K�Q<A��h����L	`q��]��dXj��)����ґ�-o�*֎���]Ny%�{��.U��
�ǂ����*�I/u8��������N虪�c�+�o�4Y�༣�3g��2��s�L��/�<�C��`"�j�m�T'�H��� �E;$�����sQ�v��ё���l��c\_;�r�\U�i��#�M��NV��/�}�N�
{�:�>/�^E�ee<k��iܩS�w}pu���C�2	S,�EK��n��%��7ZuiZf.�����u�����_tĈ��l��uٷ�e���	_�]q���_`8�p[>r�g$+S���" V۰Z�?
u�@/sn�H5��������6��3�g���'ӯp�>O�}k��P�/���Or�t�N��ƾ��-�y����K.)��_���ܖ�(���\.5�r��A-P���X�X+|�
����4�,�D�D����QV���:�5=5�T�)��Ql����T���Kn����i��3Yo�����ّ��w��
��5f�O�AĜ��m�V{%�G�mN@�#Q����RX�(��Eú�~�J%�����H5��nC��y��!\}���a~��� u��X\��_��_aʬH@6��p.����
�@�(�,�v$����a�E.��*�A��9L]t����%-(��� x����k�B(��.�a�P] {4m����îK��3�)"��aU�F��jN�&���V���.R��ϴ�`J�B�$/&�L�e~��:��z�QX��	��ElBL���� ����Ք!�UH� ����@O�N�|�ںvuF��c+f'V�;��@�3�>��@�ı�U!m�׵�lWIy���E�\�E/�՛�CJMC�ǁ::|.��v���L"-���)a@���)_���Y��
I?:x�v�{�e&��vyWQ<4�h1#)�zl��y�:���)��nI�PҾ����/B-t`�Yf)2Кe��.&�Ml����&m}����t��,�u1��.���QB�9�+�P�2�h�-��~�L�b����5h{b���`�n�#�(�C�[��p�)B������#̣����y�ߖ�+N�PJ#
��WY+���1��_��מ/xwc�=x_�1X �Q�:�b�=�\����F|���]ӭ�/s��H���wv�'W�NP�=�V��ݬ�p�
�R�3�JԲ$S�E
�P�2���C:���r�Gm��䛯ר@�_�{5��B@!e�r	Ģ}AZ�8�)��^���p�tF'��B*{��T�$q��PM9��N�u�0����puq`l;�ZF|F��Kr솴���
����	�6$f��:��\��&H��#�{#�x��Ҫ���%��-�KV�瑹S�3^�r���)�����%r�~�c��D�pj*b�|�p[-nk�MDr4�K���z���L���)���H+�_��
�ADq{�	]N�c�"'fX��a��D��%IY���蕧Q��˛7[K��հ������s�sp�;���K�DYs��I�l��=�N���Ck�����`/X%����θ��f�V���ڹl������;êEX!�
^�"�U�{Y�N�D�eS�6w�zҮ|)~���>�<m���/���f����,T:]�R��i�Ԋ���B�	A2e������tU�Yb�d��q3�\-�d���a�������Ӡ����<���o��]��2s=���8����j'��t��������-��?�ڛp��up� [l�U���p�������.�J�+_�hX�\�>��aˤ���=+J���2�KY�c���O��R��q$�m� ��zV�?y�`�N�U��M���n�<�c�Wb�vپ+]{�~+��P�;�r���Eܐƹ�{�'��C�:��Y��R���s�[�tҙ���sJx�̶��Pn�]��ۗ�R,�Q��)ˈ 1�r<�8S^�S�snC3��}X8%�!A���=l�T},%/�]���ٛ�z�:�A��	��"���[�m����<wy^�%�����{��5��t�Ѵ):�g����/���O�8l�|�C �w;0Aon�h�i!HM�=m�*/vl���:rK�q>G6T���K����q�e��nkm*A�}�=����W�0��sw�`�M� ���V����ŧ�n-o��w^X�R�k?��nڿ��Ar9if˱lUuKK��Rѷ����{P�Hį߾�nM�ub'�� �G��52���h�2z ����:S�������^�T(!�#ІG�[����2�TH-�|��]�5o^�g�y0f�4�&R��R��H���$�3<��i����0�~�#�yI�?ú�<v����F4�k>��2�����p����-�j/��SxnW����:�O۷��{�������"�͹nF��>%���[�aHUH1X/R��^u%� �t'���]5���-��g>d*t]&�����v�6��h��ME�� ꈉ��8���U��D%� �,�
\�"h��'��5[����
���`a��|#ɶ����F�簈���֛��B:�*���%L���7d}�wM����{������=�¦d�B@G�:�G�@�X:�,��l&{`���:�[8�E̒�`�Kw_�n�}�BH/s�/P|KqK)0G�9v����j�ܶ�	�am�>��SL����Q�-�41L�.��{�s�Ȟ3�)s�$��<��!��
���6�?+����4O#�&�Q�q�8Cz�{g)a@r���L�'��mRH)uM��(�]�X��
4��pZ�`�T}�#\�d6�1ɮn�Ǥ�k&��p5�Uj�QGnĿ �P���km��t��Q�*��݈��b!<d�������(Iu�J�'��].,��G��^���TǑy�����g[i����c^��AH�G�>��{�����L�屎W�N����B���@xu�-�K���J=��嫳j۶������@���k� jo�m�7NW&'\PMI�R�KA}�w��l�2�޿�!Y��k� �y�i��/�:���[�Á�'�5#w'7iC`��;	���n��Sૐ����#��������ڂ��z��zp��Qހw�~���� ��7��y���6!��c:��˙Z��8#\�k���?2��`���&�:�rS �}ׂ��*u�P�n\��M����/g���9������j�l".~C=Ҁ�ʢ����^u�h���[�� ������%y/�G�Ī
�%�Ͻ7��|������Gsy���dE!r���:�⥇��.��B税�-e�l8�L��`t W��4�r�]Cz��kf.