��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VYkM�#j>c߈Nw�&&R�u�c�@?5�X���ҧF�+��"|���������5`����U��o�x�x�`<�E���7E������kFC�a���$=��M���]؂�[a���hH�Q��K��IQ��]�uN��V՝�m�x�����ZFAZ��~���.��p&��f���ZT�u�����͕]U����}��n�n8����)��W<_�B()O��Z�N�Oc�*��췛b}�w�XM��"����'q�=�)]-��m��<?`�����WY��>,b�s=�q���KB���C���v�3k!P��N��~���z
��z��%����$��eK�ۉ^F)t��.4�$�ƈ�`x;��H��W��7���K|<������JOkR�M�S�g{��u������1��-�'2r[��f��[i��_Y���s;�����������z����/�*W���1U�7H�#�&�����P�w�,j���y��=H������6��=Q�s/=ǽ��SP��]��O��~����c�cq������!���(��dL�t�h5�����SD��N��$jm�r!�+'�Ŷ0{u�����zh:�c�['���Y�lc���[�$�w@ �+y"�G�;��p�v��(��RM��iב^��m��b$���}�f0��m��Y`Cȱn=��F��o^�s���6��W�Ғ\A��!߶�p�pI���>���	������e��,�6�A�����N����ţ[��}`�HZs��&�D$��S��UG?p�⋨J�VF�ݰb�(�-�"7���2�F�rxus�f>|�{&��T��nv�>ȷs��j��)J�����;�(�?�����:�'��O������)�J�v�7�YC�R�3��<K����f(���ſU1�h֌��X�{n2�#���S��6�ۓJ��=��*�3���*6�����s��A*� �z�>f�q9<�����t��M��O�E��U,���5�p�3NO|ߩa3�!�.���a�4��U��M����VA#l�0�� �{F��DK��OYC5jH"npM5 pg ���ݍ�����Y2O�$���MHڨ��Bq�wV����$�_��%(%r�N���K�JVܧ�ˬ0��!����ɿ�Y+9�>�FC�m �J�XD:�P�A�h�[0]$����RF� P���+"�"��[��v=�?r�'+Z�C�$�@Ҧ��e�قҶ�������t/��LH����|����42*n�VC�#�Dw��皆����Jh��r���iB�,dw�ܺ7*�F&B%��C#���Q�?q� ������W����|�/\M��L���;E�5L]�̕�o*��7q�A�/�ơ�0��P�dbB�&&���f��L��ρ��8K�>b창�c/-��B������J6.#�oE����V���0,�*U�1�!��S,��+��!����8���_��3�lY��7�	2��&���B�G��o5���A�B��2��]��J�P�O�U��7*T�޶��p�P����l�c�[s��Pö�q��j��Ȏ�R�hD)=�,�h�����Z��3vM�	J�?4$6��:Y8yZ#+o�>�k�:�r,�"s0��@'Ĉ��!
�k�;���-]�2���K��l��,�S`�v�$�Zp��A
�G���?;�R6F�5�k��4H�H�����a���* ��I7[�e����7�Ą��m,.gڢ�FC"`!�S��ӿ�ИvVJ��yi���9�N�*_7�a80�B�T��̟u��5�}�%� ���:)���������gOn�6<ߜ�f�m�wS����}�i;2�I/rp���4��)��@��t��U ���r��ԼI1͹f!CU{	�b�Ⱦ\��1(}�6��"� =�O�����V�"s��|���-���3�zWK�ر�ASG��m��_`��n��
Z�{Qu�6ԁˀ��ԁMru�9����/?��B�v��K �l����k�+�f����tA���}�t�+�.�V:�K�e!�o}��@���yQN{M�^���u�]��������m�#��&�Ո2φ��u.T߀{�����r�ȴ:

}�?a�䄤5������G�~�^�͗1[��YWW��[��k�v�8�^��"�����K���w7g�T��F8�~xp`=A ����v�E���}*�Y�Ep?��VZ%xo�� Z�2�#�s��q�w��X)�vk|K(��bR����2�}G�ho�?y���
T��i-��M����:,�ֵͭ�EVc��}��t'z4Jִ�UM��|��S8�v�V~�DB�伔�ĴPI��KT�_�̸�c���U��n�إ[�G���3'��?�)e�#se� L���$ �X�(nBEǯ\�rJ3K'�x�3��kVH�uZx�CX�뵅h_���{��gv=�5��:i�Y��견�S�m �ظU���@<`�{-N�U)J@:�pt�r�g��PUe �\+j�&~vݽ3�.�J񀡮/������eX�p�p�B���-�(��=y��y۽ݭ!38��Ua��HY�Jw��z΀:���lN�ϓ),HB
3TB>��
�B ����6 ?)�	�|d��7���n��f��Rj�u��W[����8nk��&R���~38.�F�6@�i~�~��/�k����B����!�K����u�d��L������T|I�!��0"xvfW�ͣ':u9m=Օ5,��@Q�M6�܋���ٺ �^`���9<5��%@ػ�t󗗔��M~b�U,�(�O��w��jRpA������R��>{��� ����
Ѣ��uۈQ�� �=$�r��p�SڡŖ�v|ˑ�'�a�Jy��rɮYkW��v���dJ(M���SGzI�ǈ��3v//LY�:��P� #���S5&v�p�!�"wybp
hs�()	ϖWi���*t��&�v�|.7S�``����E�>A��>2�̒�����.G�l=c3��Ᵽ�r�Ï�Ϫi?6��6_ܚ5|ڡI��eqÛ�f�w4�8�3��W��B&��tǱ��Z��+f_���>�꽏�}���b6���#Cwd��D� ?1�,,�I�����c`�K��H� h�P�<f��n��b�B�{�^�V�L�o �wŭ)�����z�h�YpR�5w���Z��bl�8�l����3n5�׎T��b[1�e{���Cٳ�oÒ�A�I�z�&^�ihc�"���	Ij'm�%w�aE4:r�\%S>���HJ�*xr_��J�%�"����GCѷ��]QY{\����ے�"i�v~�P��aj\�Z�-%�5)\Q��$�eewȦ�j%aO��>�v�Кŵ�!{VK���0���Pe{h8XQ|��3 �ut)�_-)�<��`��w|ٰ�>i�����*�᱂'YS�f���m�;��%�#������4���2���)����j"z��@�;�fe���5���!���ȷlo�B���cw+CK��E�羢Q�?��<���2fO�z�g�i�:�o�#GOQ!8��Dr�B������G�X孺��><s�:t%��0�}�>����1Ռ�����adlW�x�1t�3ߟ\����~!a 8	I�~���S�1��w�qK��@i��\�^ &A�>�]������%Ǘ�@�������B���E!7 �\�vG�%�E�a�����n(��]	���a	�[��mH��RC��PTQ���8�e�ר�V�4J��v8�:��/�-zo�ωw�7N��HKo����X�!�LX�T�z�D`�usv2���krR�Ym�J��p��]���9o��Հ��Q�_���V�Ƭձ�%�ɱ��6r�g�d��X�My(������ �ތα�h��<����|:?�%ɇ�|�ua� ����֘���( ��S�:!t�	Q������i<����H=L�P�V��zH/�׹�]k�v�?�S�	ǅL�n]l��x���㍋.Ga2
�&S��4A�Ҧ����WN�`�S���󴬗���1��m�}���"U���v��гE�}�^`A#Մ���e���Gርp��7�qf&���FXm���wSG��NX�k��S��C���EG4���O�X:�*чVF(.;�kV�Bq����i���g�E`y�|��2.~���y��"ԥ""��SF?��r�(�)�t����IϠ+��pm���4��Y3������K�~P�2��� P-��Wx�	��PO�: 6=�= b����z���yVV��2�.�
s�	C�K,�~�!��*�ȱzu_��҆/f/�����b�7|҃v�����!^j�LNY�e�wio4-V��������H��=x��C\�GV�O�A�PC�l�$󰖵7ڠ�l	SwD��mvm�߼p��Lw��dmj��ˈ��U�
[�d��\�~4c�֧�;LT�@>���?9A��fF��{�2|2@'�2�*�ε�l����.�ki����u����n�b��:���=���з@,�.&��ȩ��|��J׋@5��.K�Qd�Û	$_X�8��a� ӛʛ`]d���J�4�ٮ�c��]v����av�Nq�`'��^�iu��wl�D[~���-�� y�dˉj�?-ҴދX���^�Ӄ�,fթ̗�4��
ݭ�Q��*���	B����񜣩\Vw��2rGJfFUTlB|��\�&��v�ض�^��טLR^��>������3��t���0�ˌTp�ӻ�c�u@�����Ȝ�%�D�����%$��]	�,�7~�±�﬐���1����^���b����}X�B���  R����F��^���9}�M�������xq��TܙJ�'�����12�hn�X�+�W=�.(�~m;�N��Q]�$��ٚ��U��1O�2�w�}��C@�ή]^�CW�3hg��knt�:�!���~�hτ������#]�)�2Z��lpL,�0Ĥ�'p�0�>׬`-����4�cOd�v��ˁ�x�Ź�f��y<W:D�D�g1����G�jм�\���GQo5:�>C7���b��	Ѐ�#W�$$�Ս"�A��n���.����s�W:��-L��X��V�r/�@�(4	���$	�6{U� zg��z��"Zo4&�u�x:�W5������<����P���@û�`�����)g実j�F� ������/Q�mpX�� ��`��yx@�� �P!#T�G��Pב��qi³�r�L�s)|��'���7���J���}G�S-����w��'�\���#T���q_29э��k3��<�����(xX�7��z]2�;ܿ2��;6CQ�Av�C̖q�;M���"1sމ�
������:���8�Epq����u�d�2�V��Kl���!?�=}���]��J'����+l��\�c!�|L�4���8-�}����"������y��x��~ScCU���Y�х���|��K}u,)%Pb4�m�q��7p"�����j�D��Zj`!�,���U���W���D�	���X��䩎I�1{��8E���	�jB��F�]ٱVgó�lY
#P��2j	��fu�1Τ\�5�"ȟm�۠���F�Z�4;���j��_�)6	cL���cO�P��<W"�I��:��Ӎ��yD߹�@O�o+�o,F�����iG�{,�E�CɒW�9�E����?�06rz�4�>�e/*����lD��m��f�=B����DC�'�Ԕ'N3u����F�� ���~ߪS���[�����7t�m���C, ֤p�i+��i�k�$g,�
�b�f��`I�_t4\��������S�v1>�h*�z}nu�)U��-��m��������ɕ�e��BwY��!���W��w��1�9�z~�Gr�����ц���b�A��P=P�v�A%��q	�&��D�hæ9�22�DU��A��JVI��֡j�a��(L��^Yj�ov��WH��#z::�П�-J�L!]j9���%�t���{��-H���3ӻ�z�����
`g��A�Y��={�����4:�.e(���G���`�E�Y��a��V�݂���@����
8�����m�X`��/R/2����30%�3*��S���j�����@T�
r���&WC�D�@4Z-c!<O|P���AH��x6k��螦���/"g��k]1�@�Q�:~MB% �édw���dI��AN6bi��f�\2��1M-�3y��4L�d��*O���c�j̸��`�ˡd/2�=��/�D��\}�)�V���8���i�9�1IK��'*��c����f^���Q�Az�X���76ن=�;�n��:����;$��Sa�2��
9	��p�
L�>���<p��K��v�� �i2���xป[X`�E6�m���r����>�q`�� �q��|?@��۬�������!*ZNL���D��:��My1��Id��,��͝�7E6�N�5�>ҟCL��<J~F���<˶N���J�A(#ڑ�����jz�qT!E��=9 ��s.	��<��rC��w{�m��RR~K��q�3H�a�*v�W���ȳ5���=���T��j6$[�P�WC���{�i>�|=H5� !�w����:��u0eݤ�S��4�,zlּD�T($�?>4l��0o����<�6����\P[��V�����`�ؖK�Ri�N,�$�tmpLDL�]~k��^uS�V��Ȣ���ρ\^����@�_���-���5؂�c\.�M[{e�"|��~&&��찢����h2��ɲ�Ų��=�F��`��24�.��ڨ`�iz��2�]n��
��'��Eq��n&�\��k:�JN}^V(5(�m��S�V��y!|�_��K�՚R{;׮=L����K�H<\�L?��｝/�q�$�����b`F��:��?&V�A�9V-�������+o�޲���G�(@$5����⃸�z0+C߂�7Ic�r��_�~ד���rzC��|{�E?|�"o}���W�����^1G��NӐs@f������=�u�Z뷐�H�[����t;�+�(��tF6�nM�_�A2"T��0��B��B9rg��mo�B�&֎�lhҊF5��|�m1���ޮq���:���^ǡ3N2���S�h�)>���)�����}�ڷp�N�*��g��p焍9�����B6�O��X�Y������a��ԝ�������Ԗ�_��#ĥ�<�tu�7�+�A����j�=4ޡ�i�:�_��>*��@5K6=��7��G�Y@���Y�pi}�J�I�}�g�A��5���!sL=lQ���Nir1�~�_�rF�`4]�|��N?G{��t<=I�os��'�+g����O��]�(�]�tZO�50C�2��'#�KUhM2�� �W������'��w�ϳ@^�ݻ������H�Yԣ��� �3롵5h��|=!8����l����ҧ�8L#��2��&��W��F���.��5���8t�V�5���� 1f����A�"VMq�ll�W���>�2a��ǹpS��%W�a�	r�<�3S�h\�~���Eg��f�����J����t��w�^��#����g9w�6y�},Ҭ�� ���A%��u����77Mo�
�hnD�!���ՒR���Ҫd/�7^�6u�hu�+bNčj�DKP�!�2�̓��z���Z��g��%xa O�fF`��a�U�{�2���Hz!�(�ls�-�AVV�D�}�K��a �"TY���Ώ_>q��������8�ż��k�:2���j�+�s�`l'�LR�4C��x'T�qW)~�s�#w~*7�+M� g�ؽ�}�Svh��ֱ�B�=w��%�I�}W���:��)���+ѶeS�c��R���.�3�I�*`�����0��t��;/��n��o�Sx]/0����ki��*��K@	��&؞�14\�UOX���Xf�'��2_��ʿڇ$�S�I�i)�����syh:HWz�|?��0&a*�x���Vu}�x��cCu��;��ݨ�dO,%�����C"]�!�`�7���BJ�׊X�ƺ���g��n[�~�r���c�*���u	屠��s�]+;1ǌ髸��4��Fd�G\�����n���H�ʣEIA+i~���g��vH��ϐ��l�@�ÊA�
iK��(2/�K�kB=�������(�A��x��u/�X��O`'��++��|���Z�dS�
H&GE���J����<?q焰x3H�׬@ʩ��\@�N��ql�np�I�V�	AيR�F)3�y��(�#�,"a�5GaL���q��<w����v��2D��\��t� ��ќ�CD�Y����P�/�)q��_5)J����C���Ģy����n�f~�0��sm�
�L�v����y+�!�\3%"�F;�G���ud�*'<oL�?1ꋒ)��`��}�N�*ɢt;�ɩi�4	;�����j����M&D��[�2T#��-��D�"�D���I퓡�R�{ ��,65�i,�"�UQ~��,��%��^�*b
��Ԝ0!�
���$)j?�X��d����,/R�B턬v�M������	����}y2�>���u���*M~u�е�<#.?�m�g�?�)q���Ȩ+g�Sx��*mp�r�.���ޞ����0<TT[���K9'r�u
�k=��.�mO���˿�T�e�V4Aչ}n�0�����Yxnv��z0s�Zx@�;#��Ǐ�pY��#`�����GZQkÇ�g�h �H��W9�����y4�ʬ���Au55r2^!k+�Y�v����X=V��V��s��d�d,D0�����vS;�\ǈq�+��kG�Q��A,�c@{Nh8��M�� f6�e�i�A'����]~W��JG�L�$��F��� ��N�7�3�!�R�W��^��ke��3��PO���P�[����l�TȪj'/-K�����UBR68�%cl�\���<U4��F�5q�}�#����v��:Vـa�Qj7�񚿁�D����=�" �1�Y���KRvY
��+�$;�
4^E������불�b���|.XN^P�Z�{c0�:�k�)�������IL��+�R���P�&=����s��\�ă�!���}������d�&?�4V�X�� vf���}G��C\�L�Eql�Yb�M��dY�ND5���r\�Z�2��Ӿ*���Dg��~�&O�����ц��~� ��/aC9�Ҥ�C�h[�m�*�s|��=�v�=#J�Ab A�
�2�Nء�J᰸R?vԙ���=;��B�w�̿�L��~�M�ۡ��	�r���0S���K*[�4�����lˠKH�yO�F��Vb�J��0�����E�����8�O��	�ā�9z;$�)j�.�^Hu�k���(�^�Ly#S�L�Z�?��!��2N��ϘT-�,+��l��q�n�-`1�yNy棐��^Wq��>��I�A�oDꗟ�
�%,��-���2���`�8.?p�z�q�G3����yyYo's����H���ٮ���n]�9�,��f��h�N�<o%�4��XX��(��6��C�)����`��^�m��_r�X��̬EK��!V�n��K�7)�Ȯ���\�/z*3n�=/Q��(%�/I�]�y��3�3/6su�}<m�#?B �D�Y��3@�=ms|�e,���.HM�����L�v)�(i���){�Q���xw�|'�Ip��g9u-5�UU8��.%�t#ç�xa�te���7�؂	\-ɐ��ۊa�"d�&e���~�-�ߟC�l���4�P�����m�&x�έi����P!��D����@ƛ��Iߺ�+�%fY��l�$yT{�4���G쫇�ۡ��\�}���\��!n�LQ|O����L��^Xq�'�����9�]��l-�E��H�CnS�t��6DՅ��S�
r��9{4�9)�d���*������"V��}o吠,�����1�^��O ֍�h��ѭ�C��ӹ�~��m�OM�q#5��U�=:/t��!�>�^� �e)�Cܵ�E&���Rl!��W�k���k�H5VU���4_�,+/#��̹�cȐ�Bje�';�D;�8��!��s�
1�������t{���u�:�5�0n��-�qN��U|4�������2�ü~�M}$�(\��723��Mpwvu޶Aۜ3h&�EȺ��R��|�Uw:�ѽ`��O�j<��Tv?�1�^5��W#)/�i���v��O���[Q�I�.�[�'��?��6l>5�����KG�$z�2��	�6�J?�7�7�� ,�q=:@��@�%`��\G��A�$�<�Գإ�	�:0k�GE *��.�#��K�^�G�t����M�e���*>e\R)_A���b٦�ސﱨ7��O���?�4e,�ÅLEn,���$;�ߦ�kP���U31�}82,�&�܅�!56�f��R�	��r$�%�����X�gh�jg@�<pa�vWa>�z���h�s�(�ˢ����)���N�R�mnw'�@�GWt�SbY�o�k��Ç� ���R����<�/���MA�a2��4�U�K0,�mr����+CP�wX�t(Ҳ�#?!��~�O���e��t�=5��W���t3=��AxR�������Gf��/Rby����G�}�{X� �/cϺ��'_2C�xV�_ �Z(ق�ѽ/xs's�F�#����>�,0�oڂ�W:�j9؃(���ߟٷ�>VU��C�\:��p��PF)G�0+y�-ĎxK��U/��"�B�a��:Q$�>[�րR��<Sk�����w�{��VCӓ�^�7��k��5H@V������^�HH�f�#���C����]f���tW�"|=4N˖Y]f*���Oϱ�ߡ�ی�$�{��d�ܯ@���O7\�W�%G9J��+�Hz���ڰ���'et잂�L����j{���6VΤ��E̷7����[3$�
8���r����Pz�B�y�I���p�Z�LO����ѽ�%�������ge�#�	��_Z�c�����
�!��L�e�����\� ����_R��E�Z.�5�����`��]�����V�ׇ{$o�z�--Q�QuE�
���P!|j�J�{5���)2������0�Fa���!6��8quDHڳ�z:�'�Zf���q$[x�*�"4���hW�CB�"��FK��?e�]��D�Ȼ8Sߎ^�g�_����
Z���=_����ʰ.r��$�����3��f�%� P�4��ހ��D�:ˑ(@���ƕ���kj�"5)ft�#L�U?-��=�`b�L@�S���{pD�}C8Y4F�.��NCG�<�ۣB4p���i����@z��7���[Wv��'�u-<��7[U�%�W�"V�5��M�*��_{�^���N4n4lm�	p���
�E�������h�@�P�(u=���a<'v��It+�儼a��Ղ���\����W�19BN�0�h��cϬ�ŻO� Z�ʅ@�۱l���]CH ��4z�PEh�u��P�y8�G��C3����%ɹ�Li�:��3��jj�͂T���ˤyT��3 ��M�����N�"7�֯tN|���I�Vż�O�Uu-*[���ĿS�+��q��o޸�@��u�"
�e~��la��[|SBo9^$&��� qB�y	a1��&�0{=$���I�.�����U�������ؿ��qG�rs>1�T�3�Oh����#B�\6��������̐ᣦ�h_Lc��"�����jԭ�
�L�%(�x�i��0���ѩ����炪�`�e[˪q|�>���b�����&H�cB D���Օ	�@��AЗ�=��0�tU��c���Y ���Q��<l��H���u�t�2o�l
��JMov�X���]�1�T�����TX�sHx$���ˇ˗NN�ۇ܁&�M�1��-�ɸ�t�ۥ��}���x�p�:7�'��@�t<ȼ���>Ԓ��,]��S!��5������N?]Ĩ���Z{!�6zM�b�DH<�����T��Q���ȼ!�`§�5���Ⱦ��Qq�lwܗ#�ԗ(I�o$�k�{����;�����3VfiCm� ����VطԨ��zż�0�"���	e�3`�l�D5��<�2�m9�x0W��T����@|�P��0d�O��� �
�]�|	����� ���WT`u0�,�.�`�z=+�Pq�N���1�}iӅ��Q|F7�������T&��FA�XPp\�W��K�&\@�^5Q�ڐO�����[��M]	p/����r�%����nΆ�Ih�"����݊ Zlb�4EX��Kl'��"-L'.�s,S����zA��*#F�ر8&XP�1hŎy�TaD\�;i�&M���<$��
��/&*�6�G�P\�Q�޳��ɋd�����z�/ꨢC�|�[��&��b��J��R����>!���y�����xpu1�W��: ���t%P	�
�o*��N����6��r���*��sn���_h'5+��bHB�y"s��w��z��=�9T>X����'/DW�(�����g�k	@[�H]V ��ƒ���4���{�C�<��Whۑ����$��f{N��i�;��N��Cd����C�;@�2��O�5a~>Wj��荏t����	82䟗M��g����ҍ��gj��jb�����<�-��C?QMM�~:�����^�䍅�}D�d�iu���)i�{����\TQ��X�� �騈�>՘����+qk�M3�N�l�� ������%��TE $�MyjS��L�}�x8e&<<�N����qu'�fb�Nr��sa=G�ݹ�����q֯�b3�qs6R�#�Tw/��'0�C��Q/�c/�w�ǳ��`<ɗ9eEN)"}��jd��v�����V5�����ǁ���ړ��[�k�s��V�(u�vFh��flw��umN� ������467@i]�j�G5J�����x���[Ynb0z�|$eqn�X�(#v���s=u�ؓ�[���շO0bǨ���\����o��-�m�&�b���w���q~��T3���T�5���e���&RA&@jp�~`�����p���{�s�
�ߪ#y'B�SQ�0B���j���ݢ��L� ��Pc�@"�[#�F�b�	HN`����	h׵X���չ�,��o��N98ݎ,A(?D�H�6ͯ
5������,���Ȗ#<gGh�P%�
���* M�I<��ֽe�T�:�"[P5���q���Pv�ߣ<���٣����k�t&��9������wyk��_���8��o!>a)#s)��"x�bN��LQ�$"� /J��y�F]n�d�b!	�]�p��R�ށ2����
7�=-����1+�R_H[o擲z"�k�����ޣ��&���@��J�!`1AT��qBWfO9�$�3��vy]Î��>b�
�H�a�4#G0��L(�4���	�=��ֿ@��E�Gi9:�M��[;��VX��'��r�/S;��=L��<lG�4����aS�K�ܷc��1���p�̎jh{�X ���Be��ѥ��
�l�N�Ȅ�~�P��X┩򽟴��i�|'�g�EK`�ϫ}�E��m���[mߧ+;�㗤�6���7����n��%���Ƣ��A��
��A�[O�m�c�׮F/�b�܆�*�sx�`X�/�mg\6e�P�`�eOϢH�!5~�됪�tuV��~Љ�k�#�P�4�X���ӌ��e�1�Ӗ6SB9t	#:�/C��&��0D��Fu�;�ݖ=�C"1m;sCd)xw�������,h�˂Hp�~څ�i�>��A���y�gs��o%�k�o�k?�B��R����9OmKPB`�o��{EKD�+��D�P�zG�5����b�A��O�W��{��[�:�3�d��џe��̊��@�S�����UEs�u�:�i���7Z��Ed�ؕ�a��|�����;���W#���c�F0���m��L���,iԥ�E����9�|7dg�Qr����\7��.����&x	=�	/V6����{�Or�d�L��`av�yV�iLL��etY�c(���y>)�vc�7�s�v�%�v9�k��B�h'���l	�0��0�Gd�^g�-�h������;��F���g���9*M�nbkwO��"��N��=����E�7'Zv����1� �s �Z¨N�{�Lq��m�iT;�����n>�ՍR���KB�*�4�hP�b��6���k�qį/cMF�|^��7ɺ:y���u�G���ZiZ����ly�@:�*G_	o�O]*���W���:�Mt>�@�;�Q�RkCEul��Pv+�I56�nn�L=7o���̃��2H����� ��w���^_��$��\��F3�8<UҘk��NDBP�ؗ胐���ȭ�3�D(�y(z[�ҽ�.��K������é�On@�&�-���K66�Z��H��6��C0���rv��&���,Y�|f�q�q+����S4�EU�Z��L�?m�~>�]���u��ڟ�1���)ll�����J3����i� �X�T=�`����m��B5�Y�Ix�<#�e������2��<53�.�LܗgR,�}E�="��j�ܪ~Y
���ؤ	ڣ�a߼H�Xk�� U�i�#�t���T�dIs�t���/~3�E�O�:|�,�6ú��m<9m�3H���<Y./�8�1��i��C<��+��u��;6,�]Xհ\$��5}m�%��6�>E���\OoZ]�ʣ:j��b���rT孥}�0e��ދ��-�Nvp�9�p�A�抺�<��gE8�n���&��Bx�dܓ�l�c��L}w�?�^qrw\ŉ?�w}� ]-e�0�O3�5��Vn���"�35c�� \!?;ߒ�c��C[�
e��݄�'��r} [i���jlTsƉ@�|���zW>	X�\m&Ab�N���c��#�zҞ;�hO(ǽ0��d���O16R'�i���'%���¾�:���XP���G#νr�Ħl�'�D���%+8�u�(m�q���/��Y�� ��[|�r�W��٩c��x.A8�{38�[Z���q��Dkvs��*B٥op.�]��)ı�F�H)��`Z���:]��]O�#[ ����Y]=��2٥u��p�1P'�0�9�	��5qD�9�NY�O���V1s�l%��|�؟ƲG�Y�ٵ"g*���e��ەFK�(����u�k�� !L�E7S��a�Sǟ����{gkk���S�0.>A��U�<-|z��+�J~��柗f挡�h��_̂�5Tax ��Jx؞*�O3;��/f�D����$N���*Gb�&�Qyl�;�4�A-�då%�k�����~�U�%���밴掂×�+)�
��@gqC{Muv'���1�T�CK.##=@�/�JPlt�C�29��:��eݏ��0�6yd�|��J>w3�7᧭����4>��%�(-Iɔ��h��I���9��p$z�m�S���(4���r��Ӿ�>"�ۈ�u��������K������X��Nl�b�}�y"�����+NcQ� ��Nkm$����0����*԰���iVօ�0Nu��r� 9��@�k�]��(����܉wXwe��W؋5�al���C����TB?f������S�zI��K�κ�L�0�#,��N<N��*&�f���J��5��:�_=4�+?��A���<f�N~>�U'���`L�'�7�#�.�F)��"d�PH\'BF�T(����j���Վ�'b�{��fڋԲz~$��Ł�X��D���a p�*�@~;H
��[M��n�1R�1�h�u����:���*�f�(�A��,���
@US"�@Mjs[�w��*r�l�ub�&_+��ڕì�[�~��PǮ��}��y��M7�H=mO��nT7�ٿ{ֵz-�-ȥ.�ľ<:��$Wp���H	��j��n%,��荗߃F�Ħm�x�kv�1�<��O=7�̃jZ��K�W��?�WON��/�>�z��k�����·��X��2x����1�t��dv��O��(�W���i;x&�o-\���TD����:�>��[�y3H�Y��0o��8�73�ڣj�����H]���#��gXo*��u���G��
�N�h��ȾO��С0=��h���. ��)4I��w���>a�⥈��B,*�q���9s�0K�%��ó�L�d� �}|+�q�1lEGB�2�y7n��j�"��H�o�E\��@RT����=P�������S���*֞x/�h�K�1A�\!8��Q�:�l/� �//VE��30G��7�����(�U�Qq�zKv(8��r��(�J[L隓26�=-���C�ô�oȀ��\�ȨD|�Հ6#���Ёr�=!�)s�y>��`ᓙa@q�q�S�,3 �x�4���9/zn4co�
��k����M5L����f-�I�Z�����$g���>���b�5��*���a�ʉ4��	?Q9��f�B|���S#��hH�\8��W�k�|SX�c<���%������K��r��nY��i��ʇ����z�J7�P���}�=�G��&���h��l̮X��"�?cT��%L�H,.a�b�T�,�G����2�����.-4��r�-��+�DF�%7+�gOR;j.�El(�q�"�7����w6�-�GA��\�Ѝ�u�b�!�	��p����ۃX�#����������eٕ�{��^n� K�V�T�&�%"=K]v <-��'IG:~��>�� :��Z�������^{������~�{c8�ؙ��s���2�(R��h����Ab�]���#�2D�oȢY޼��@� /
�=��**0�{��d�Q�����k����*�!p���8�˷kd@����=է% h0�_5͋�g�ɽq��t���IP#hϫ%<�_�o\8��P%X�e�4p�W&��/c�Gج��a�N7t�X/���T����(O)�a��#`������S�x�,���u:6�=���I�q��O5�z.�a��#�����.�?���/ǅ��ð��Ż�S+~�i�<-+�oS�=��!r)�O3�s�ExS��n���?��j�	���3g��q�f8��j�Hѡ��'w��]�r��b$�T;'"��:8�}����|v\N>��u%�����l~�$�"�v�E}��<�N���c��Qx�*��enQ&�}մ�XK�x��X�_��)Q�IF���T�xJ�G<moX�~�F�3қ�q��t�� ��c��=Hlw��i-���'�|�r1��fՔA ��͌��[��:��<P�c�̕7>�<1Ԓ#��t�&顛������-J$)?9V��}�\��1� ȣ�Q5���
�e>.�­&�R����ߵ3��ݑ��d�vD�>�dĮ?�A�x{N%V��FΒPĠ��'�[�^$��%�l:;h],3��f�0����2�
���>�E��M�S�j�l��ﺭ�yA~��ݖn�}Ai�f��u�2[�>R��۬�����#1���.���Z��@+_;��b�	[B���e>H+��V�{���pt�k9�k�3(^��)�����Dk?;�E�еAuX��m�wWm䳤�#髍:�5�R0)
���{a�;�2B?{=?�?YC�j��Җ/�Jz%�����o��Ds���:
�C��Z�V �x�?̺��WpR�� ������������m�I��8��t�쵈�]���It�l�Y*w�B۬?P1�)bS�u&ՂLw�o��XZCB��aӴًC���#c���_�����P��Z�F9�^�a������(��@T%���gG�VMZOn�{�NlHP�;���Q���Tı0�����ʳ�m�!�O��Ö4��[�3��8�yXRnVȈd�WFjK-_j����m�$J|�m��ɹ����&��Vt�Dq�G��m&m%�a9o舍ȻBZ�G�.:���WGL�/ޅF�;0�R��Bm����T1�=��s�ɠ�7\�̨���p�24 �ԭ�o�Rh���\�'�QrJ��%h��7,�Y}=Dvwt�q���J(~��d`�r^ 7+J���gY�X�#��-� �6�{��:*�2!Ǖ�<>V$K�޹��7<�<ݛFk��@^�-�Ym(PTm�b��Z��M��*L����g� �w��