��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY� �T�Q.GE�@�N�\ T���@'� ��+��7L�#a�݃oX�dk-����qiѢE6q�A� ��]@���1��jx����jjP=�^�r_i���r!d���|m}�<�>2�:	}���/�Lմf[wnhq1v��-jp�?n(�)�\���X�G���hȱ�"GV��Yٷ�{2��g�������c��)���%	87�/��%�� �?��.�ƅ��oW���lH�l��.���s2^Z�ߍ�yHh˧N�ܐ��D��&r��6@+A�C�#jY&R��:d��=�����]��iR�˷a��.U	���@=�4Ow�R�׳��u�f!#�̓���1��J5��)?�QI�w��{x�ok�H�z^���%Mn�0���N�<����K~`^��A���m^h����_#_��OJk�ҵv[~|c_�.|L�f?�.s�����Գ�37M�t+���k�ɭ�ݦU1�!����2R��X�n���3~ޏ�$���6�'k~8���z�o�s��yxm����Jo�#ח������M�?�\6f~LU-�Y?�_(䡻�|2��˺d�u�_�l�>��LO���r_p)ǼV�j�\o"�{��H#�k-ǥo�Y���.�T��?U �k��Q@dbk�:Zg�^�z[t�(�6���pFD�mJ�����u�� �N�R���SH�����RwT=��V򥁢���w�ͲR��U#(���%�V�[$2��~#�5!���UNN�]`�ǷȊ���ƐC�p�������{���K�D��ı�^���E��ȋ�6�n
8b�!��/&O=Ym���9H���	������-G�ư�)7�$N�$�j�j�h��bvCGg�
�ؾFX���ډ�M�6|���b�K��Ӫ	���G<���8+Ϧ���l��gC7h���mz#ua�gc�#�Q����L$y�1Yq\���Y�hͷ;��a`�����YR=�?�̮�����%�_k�&��ج�L^��a�Q ���ci�C��d��x?�f�#�ht|���e�5����1��1��]�lb����ҵl_�񎱝v�75!ц'�ʩ��U����b��rHd�D�F<����$vo���mD��w�=}�	!A�����K�>��5�"�'��z��S�����+g��ܛ���k�����G'ErN$�6H����:U��OR�19����7o�_)�
�_��G��`�b�X�Qrl#HHh+�S=���*@1N�U���׌��.�ڞ���K�O���ɕ�2[��f�[ri�����iߦ�_�p��熵r�~N�5*�fX�8ti�Č�+��lk�j�&�t]���Cq�z�a��w�����l;|���3v�];����F�	K�
�&@�=#klE}�
rn�0�s�yې�o������'�q2�O��-g�V姱lS�P���å��p}����L
d�Z Z��[ꮾ�!R׽���V{����] B#�_�[BP�nO`�!`� \��#�ۈ�03�`6�wƺV�Y�B�����-"�{U��Ƅ���"��z����ad�������_n�c�8
O���m�e���>�Ŝ �5�Y��@����e����y�V	�^�&�D�?�	�L6K/�I�D����brc�_�T@#��g攱C��P�����K��_��t��G;�f��y��qL��1�,mΚ�2|��(���(�P����yp��`��
F#t'.D��!5K��ֻw$će<�È�K�uL�������dRW���Q����jh�͠I�. ��XN}X����a��h����_�-~�.L�-�>�9ʘ�>�
&vj�򉉝�ɱime�Vvi�r*�\�Ȍ=֊3�@��)�c����� ͗Z�0i ��`��:��MYW�ES-����7g{)2Wr>ܑK�=��ֳ��ιv��O��V���jk����T�5�S؁�8?��K��#�N���n��>��wkm�DBU@J"W7/�0�i��u���.����/���!`���h.����!����s�횓�\����Kam@��HMk�)�$�+阞`Y�@��ƣ��9]P�.��QЂ���t�� A��^��UM�MI���.t�1	`��a��N#���u��$����o}Ky��;�|γ%���>ݘ��	���a�7��c�#�!h�g�h��;���4{�>����6U"���y��Ո��F����BíњF��K�:�aSNoj��������������Wz|uʔ�3��PA����OΝF�Ż�K�O?U ,FDd���E"�Ѕ�4�V�lm�؈Tc�r�8ר��m�W�+�`�3�
�2$j�.��day�5�k{�N��2��Q`�xQ�^��4�8��j��3�8��Z��Ef̚�qk��D����Q��A���m(���(�<�ޕ�7 ��d�	����%w�\�iQ ����\�s THi�N�l0L��g��(ɐ��rs܁���#fĄ�����^ɯt6!vp<8p{���,^���V��v�Q��T���(�B19����n(���q�&N�ڮDC�cR۴_l@�.]dw�F�\>Nl���}OP�\�R/ȯ�=�Z@�����H�(��M.��́8ߠ�	#��^�ڤ��΢���-�fO���F7m��rw�
V(�^�u�v�G�A�;sGM���c�2�Y�Nf�W��)]����2�:�S�e���M�e	�{���h4�a��ԡ�߬��خ�����y��c�V�x���>��pP��ȴ���OHyZ��pt>���Ǣ�ʿ���_K�Q0��+q��HƄ��"AWo�3��q?_�>�	�R���'����(/_� [�qWo?�1�#�;�ǧ���T�(=���y�k��T���	��J��A�?��|�TClW��܇FE��=%o|됛�Nqy�"S2�FsA���;�Tq��T��Ō �#��<���@�#�K�Bk��kp��;�Z���:�#	�\<f�"�}�T�E4�E3��ɭد8Z��o'G����p��-B��3�RB�9�6�)e�N+��j�_�B*�c7���:��l�Y[��{����k���//�^)��W�$�~��ZZ=�]7��Mo�J>�bK���KPM��̗4�JP�����51���+6��#_���r|~s%y`g=;�C�$�m���Bl����R�#�gVF(<��s|~� �goF�]����3N��2>Ĵ*�7��)�A'��#��a��˙5v)ȃ����!ҳ��w�يV�p�Xg�J%�'K��jP��qp����l*�(d�u��J&!K+V��6L ����W�o��r��xy�V�?+\V���	Q[=���d����u�w&DNԟ�ξ���Q%9��j����4<�9+`�������2�񘢇Hs���5���,��ϔ�����F!���tQ'���6�TV�M���ѕvD)]�˹{$�`�H~MU�dE�B��H�D���$ay��~M�J'*�lU�Yv�ݶ��l|��K�a�f*�N���yQ��3*W��o̹�}uK�!|̯��L�nF������N�w��[��� O��W��^��r~E�0�Z��:��շ�D�&����D1u�tq��8�|��I�[eG�S���˥�X������Z�u�n'Ȅ�W��o��>iYH�ޙ0,�YuE�-�Xg�`����n_P3` �P�@��W2�{%w�	����8��[�'�ȴ���~DWK��d��ƯK[�vqL�3��}D�+���>}�;�=_$�E0
�0�uo;�؟��G�'�A�-�#�qy��Q(�" Ɉ(�eeAj�@ZBQh�^�8Lh�b�\pL�����r}��AoO�J
���S�Ǌ��a"?�ra������g��2��$,>|ˣm����KC�����1�!Pi~Z1f�͚V�i��N(;��,a`�����.�Hj�\�T(�]��>	%h1/��ȐP����m��$L\�B-��,����=v��)��ͯ��bhbZE�ۓo�Q܈-
��#��^^�.Xgc�|Cқk� �q��;2r��pE��H+0��:�؀<��2��uE(������t�Ǭ��Ō��pBf����Cr�(/� k˒��EO����([u�e)�a���?�����_N)�V)��ݭ1�=�
1�50f��w��Vj�:�[���u0&����pcU�P��Fg^ͿuݢR����nXe8rUn}M&z!��\����gg�����9��2A,~!0e�F�$�[�xߍy�F*V��IF� ��B������ni�)�������'r�.����r6��u���S߉�d2�=������XncL:-��s�m�0���:��DK��YuT�)�3�o�y�M��rD�HBz���L��7����j��A��p���;q�`���:�3��|�O~�Z�����L����fkm2T�P0���*����h{����5� �e-+���3���i=����fKv�]ҧV�)X�>ޟaT4���}� ;��s��Xʭsi$� <�ޝo�@I��&�����V��!h흳��!��0@^ID_H�崈�,z��9�aK�b[��I!�q��<�H��T�Vl���F}�n8;$ c��c�wPk��T�k_���%Q-�{Kx��6ֺ1*��O���|�8��ڢ ��0�#�0Û֊�,k�8�� 5M�S�q����._F����I��ǔ@�Z���8��?~�E�Ԩ��96$�h�q.oIUn���÷��Q�:	�o=�!��tz��̉��[s�P{�߯���A�>�&��ɽ�m�bN<��a��@)�? ��#Ko�x���i6���D�h����|n���D7$|�S�������������d����뚅XgA]H�̎��"_z�d��ߘ`��M��S���:��@C{��.�8��ՐT�"kͬ���Zt�'�<r�y�5D�;�=���Ab��I �<g�t��V������غ�����w+���*_RX]����e:	����l�@���[�ʎ_�X���ܥ�iG�C��)f���/0r��mg�ǰ����5j����؏]��:���ٜ��/A��g��^/� pJ،𦆦��睺�.�GF-/�p�q� ���D+�����&�8�?��}~�s$ь��%Ӕ��A::�l:��&'��G.����eC]���#T�+<hu�|�w&�$�����GU�<_�?=-�}���Y�wh%�U1�dR�=����"/z�	�u���*��hB���-"bSo%��Ь�vc��@��.�]	����%O���k{�|#�F�Lm���%�t�����I��z̅�$a׺vy��'�)�OA��E��q�@D������+!6�3j��)�s�^R]����[}���:�Z-�A���'��^mKZ )ӹ�#����f�%(4H��Q\&.|�w������q�r��%m��I��� 7Ӯy��T�0�$��}��-6��Uk�c���Aި9�����H3��~ӿ�(��V! "��;��T]�G�����ϲX'}��"rR(HP "u����Y����:b�j �\����ؤ���J�/��A~#FρU�i>ND���e["�لl�H�f՜����W+�Y��u��(Mq���@ƣ���L�،�NŔ.�ɌR������N�I���������;��k�o8���x=\N��MaؑL!^-���o��Dj '<,���jsR��o�A��R}ӎ�Vp�Ve����n�)֚���+a���ވ����C���� ��J)���T
�0��$xt��tV�QD�ˏ�S��#��[���v%��S�6�ʶ`�=�nu�Y��Ei��P��|qB�D/}�őVE@���i,.�\���ܬ�/b-�Z~��ë�R��E�x��=MU>���]�: �i�a�\��x���a�� ��D���#R���zE\�g�8��і��Dz�#���ㄈ�R�m�Fg�c�R���Ћ���L�\H�CD}U~1N!%����%ҧ81\&V捓a|Q�^�W"����@+� ����;d�c�K"AG��?�D�*i�*��8����w�0|�n�
{��ܑ� =��p���be�A��q?��A�k�y��;u�G~�;+��k�-rɀ���%���-L��&J�8�5����A4Rʠ��S���OR�p���ǿ��d���]<?ԓ�,��6I+�	��v2�b��\ÃA}�|��~�c^�+ V0|w]X�D4������z:�/��I��-���������SX�e��/;�Ϟ�fI�~��n�����%z�\�+)K�l���/Q����K�Ͱ*�	��5$�t�m��R�brO�
ฟ	$ܳ���ܜE�9G�n��R��;��[fT��Y����g�e�����J�n@�0��Z�K�R[��S`�M�L��e�[e�N[�sE	�dQ(����.���B��Эp9u�$3c���ź���P��K�I�<b�#Em�$?�-u%���P|z��z�??'B��F����ƺ*�yN�5��;~I�a
JN��� ��X�1���uH_y8n2����#���6�Y�,Q���eO�a 僷�^A�����S.6LLi����Y�aQq"�:����}�Յ
ǻG�8���#��OH:챧�A����F�ua�x�y��2D��8���Nma�R[�3zˌ�|�W����]"�A�~�)��Vp��E�w`��_���%S�H|I!�M�忥%=7�Y�������{���yw_��Hً�W��U�/�*���ܹ	٪���ģ��|�3�%��,���m��R@�@�2r?j�����H��k���z����e塷|Rkró¬a�<��=Ʌ�W)��5�B�1&Ő��<����'	x���M9�I.l�.���,m�U�BV��6�����*ͳ Y�4��_����Vz�^� � =|����Gs�
ۗ<2��5ʖN����{T��ؑ��ק�0�
����c̔;7��"�.� ���|i��E��'�^}��`�2;�8���a�3{�te�J�ITۢ2�8@|=�)�	qR�� }�'x�������`ظs66���ؚy��KF�N�����ըq[��#Z�QW�j�sw�Y���e&�`6l�3��t���4;&4�9=�:�ǰk�׼=�q2G�0�8
��հ�U�L��� �`���>�!X�7Y����v��8$E��c,�a�G6�P1�1�-T���:O�����w��t�N��,	 6��wY��A��J�= A��c^�'�ޖ6Z8])����D����(�sc$�m�.��w�f@�� ׳�]��Ӽ"#��[3"�z�E�(����y�*����;�� ��w��Y�?���dƊ���*U��ٺ0Y7���?�5���s��?� �L�z���v ד!�O���*tJ��X�ƕ�\A����o��E�@)��M#8z�T�@�0��:�?
��I��\j���H�c�HEG���4�㘎�r_���0Ϡ�ɷ�Ҕ���jT��%���&E
c[��H���K��JCMf�� ��!��B���T�e�GX��-��o�j����`�L��WY:*L`¯���N:��coԘ��o��7@R�����ˠ7�
č�]�w�{A^�th�j+���O5/��F����u�O��@f��9�*�6�&h�����,�GNՅڲ�_�t��{��#PQ@,k��&K�����*�i��݉���r]2�����w��`����P�oz<�4X�/�}$� /�崨�l�,���׽���7��m0ڧ���n������}�&D�y��:�n�ħ7�pz2҅���eCkߵ&����v\噜0�;	���Z~E��ۼU+����q�bQ��`u���^��x�$�)��|
��\E��b�p��A���B��� ̈��V�4f�������Q�۞*�ZA��OJ���g�8!e�`�0�<n���VP��tm��к��..�.�zM4�mN�/f���{UϷ�� E��F�nB�)i;�V͜^�Wh�E�p>�v'#=A� �/�@2Ζ��L�2�1gc��l<U�U���lʑ���F��Bl�&?�>�����:Ց����#UH���Ә@ȔT'�C����}��5K(�Q���Ь����@��Egl�-��N���TҮ
��p�5�TeV��ח�Ue�"RZC��ʥO�	�5,�a�d��=�M���u.w�\��9��,V�k��4P�̈́B �i� ��< ��Rw1��7�b5`S���โ���j�ե�Sʑ��/Wx�Wxđ�����P���w
�	h��S������<�VW	�����MQ,�d�2��.��fD.{�ud���n0e��=TG�>��~<�d��,W09�?�T����qKq$��������!��1�/)�j-'ģBAS�Iq娞���)�J��dp:�{d�����^_�ʧ-$˟�&���Ӿ��k+)={kّt� A�+i���]{=�ɐ?�^!sɷ�$ߺ��,!0��C}P�^�v饁3���r] ��Pj|���!����c�H�;ط��	�x��y�c�r \o��p!��FAP�̪���R�EJ�~�uxɽ�]<^GH���}�C�׬^�D�mM9!QN�ڷ���;��#0����vu�I%
[���B�A�)i�!��P�:\���vE%f]A�*iaa<�1>��/p�b@*�� ��tGk�=�B���e"gG�S(T.���,�f��/�Cy�15>tĻ}�n��"Em�e2��ŻJ�'����Q�
����K� �B�(ccی�1�����%-��n  Ʀ���k�%"P��zs{��� �V���<�gh���}�9j=-u�!u_�#�pǯ"ֽH���57�2~�Jo]*�3;o��QcC�<��B1���k=��C��1�=�kK	�N~b���*�;I:�6)�#��MB��U,���U6�Є?� >h���T�ώ]l��Rj@"��^]�g��^8k,�G�@�LӬ���O���,2�e��rG����Oz%Wr+v�8�u�Q���n5��/%���%��˃��
o:�
���@��=�Z]M �:���=f�-��|��1l��҆&� ���L��e4� ����?�:�X���e��U1�n���6+�m�v���&�*Y��Գ��-&�����;�4�m���jI�p�l3��p\|6�s�����0�ȟ��� ��X���4M+9�l�k��js�Jy4}e�j�����b3b�{�<S���ןV
�����Q��M'�t��ƍ��"�H�O{[���F��:\��_HM��u��$�80Dl�۹�u��@��[������قq�T�uy46����0ŤW)Z�)�#�~h��i�ox�n�feRo�=!������y��aS�0tk�*]@Ԁ��j�ܜ��6�X����zz�@�7~�QQ����t�6l�6��כ|^ӂ�NF��y��G@q*�r�r�a��:i��
���U<�N���1�ȆՎ�a��L\��X3����t8�F{��~L�/��9�-p����v]�����w��w>���ʟ���kPJ�3k�7)D^$�}ָ��T**���c�ě�u�'< �)�B�Ց�cd��ʵ���kZA�2�s��9p3��6�=�1�9uSM��̃>�PD:�U=lcx���&tDę�ŗ�w3@Mf����?Y�7uf`_�檖�� �LOѬպ�IF:�r��I�H�f,��<��M�C�1��|�~1� �/i�uZ�!:U�)7��A+�Ǯ�A�q��ue�!G���:3[�n%6��=�����^��l�[i���ѐ�T{��	�Ӷ]���a�+ʰ��L*h.�ų�5zᓽ�s�����E�A��rhRcsY����oDtO�ɖ���piu����)i��i�\"ƈ�t�d���96�΂���<v�������gV
�O�/��`P9�5���4��ұq�?����H&��ےP��s{����<%Itu�����CvF�vԝ�dib�n�yP�hnoّ� X��^I���ig1	a#�[�oP�^��p�������X�i��N�j�����DO�������d�5�v�7Guu��Ѫk��G���}��C�j��MqE9�Y۪Nŭ*�r��`-9�0��x�4�(��L��d�>KS�j�����0�CLg�����8L��'������_��w��g&�4+E����e��tV��>�ߐ]��(�G�5���T�BY_��:%>������/�w�	
�K��t֪��_jX��5RrO(OT���ԯOok�g����a>�8A+���_bUi�oo�D��r��% ��]1�s�Ԕ��\7,�k�����6�'��N_jPw!���|��z4������޻\�0LKm��M� ٗs��[�א��ޞ�	#��q�Pz�Qn����[bx���)2����� i�mE!�0��.�_$�"��&&��DZd��U8 �{*Mj����Ͼ��r����O�����|a��`FJG]$\r�ˢ
=Yw��d��3ǫȜ���$�EN����zE�m����5_�Zn� �N��N]�ʼ]z��Jf�+\�� >��r�j6���	]u 
&u��������j�[W�9Ψ6�З�h��]��q��ך˸��^{�H�Fm(ZΫ7Ғ�G��W��v��Q[��W�xH�K��<ÇK��v0����QylMw��}�0����X��L�@���M�~F�ո�S�ϟ��x��ń�k)廼0�%�H�4'��ҖJ~���Z07��[���%V<q���XN�����AqzP0�\y������G��(�@�*��