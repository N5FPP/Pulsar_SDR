��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|۶��-�Eݒ�s.P���ޢ';���SS@;t@��֗��Fp>��6�{������(|�#�����jҜ.W�DA���><ugLb:�	�bG��7���S|GA��]` ^�G'$ƪ}?KT�.�<�<)�rX��}�]X�a��dp��	j�@��΀L�Q�$�M-3�I�7�,��l����O'�떴���P���[���b���?�yxWN��GRzбOb0Y���i!K�H���P�.WwH\��nO@�~�Q�?���a��)z�oE�ؠp��?ff��j�0������;�lĉ��+��Qs�U�f��f<g�ɿw��$l�D���řmY/yCw#�ӎ����+�,i���`�R�L�����"��>zc���>���Of��>����X��ټH|[��1�Bu�!#*;�A�����Z�.f�,�+� ��T�#��b���w��|���̑�z]����N&$�X�i�'{�E�=y�KV���;��"�4Gz{�elw���:�_�EY��zrd��mV6�͐�^ +3)拋=tB��O����s��E��!��(��y���~(i䐥b<�pqjWd��["/��}��� !�Tw&�����6��s1��g��Ț��#0�ȋF��~�9+ʯ�d-��	��l�Ԅ]�pP���^9�qD�#W+'�@�O�/*��o�
bŎL:/��1,EZ0�~�Q�:hoS���lS�Ӯ�����^9?uD���p����������ba�f��:��
X���I�P;�]b%�L_'��7\F��@�;#����qy�+��J!�M��P�T]��V�-,8yā�#��܆Z^��h�-��/I?�qQRS�M�ޥ�����.p�� ���L��z�8X�V* �Gu>:��Rz��v)˲���vEaz����=㮡ʨͺ��mb����7)�$J܃��N:ߪ���#�H2SP���M>��Z	�z�\��碟I!��,��F���{�5�(��,.A�N��>������qO6 2�w"Eh����g�=��j� �A/�J�*f�1�i�a+�Ǵ��0!�<�����1.R�)O;*w�Y
6	a'�7�:�;�cz�3�?����)`�_��u�XqIE�����DH&��>8���R<+�G�����z��6T_�l���c���B�޻x��{ҿp�1@�a�H9������]t�: ���p|����ߓ������'�?��^��#p1��&aD���~#�P�s,%������Б��!d~~�������e��jS����F�^��/�xb��ݧ#_��BS�Z
� ��cQw������+Pk~j��K�>����&dT(��Nc}�Ԑ$� �fgn�v丮����0H������s��Gfģ�����1�n��ɰ��������OR,^�}I�-������h!Ν��G��Q�6/er�����P���`nH��Z�d�|P�{G����cӃ��J�W*}=����b����� '�?��Gkרg��o�@;܈����2Y����^��з��E�sub&��թ�a\�Xu�%v�M������^yC��̄ԅ�	ٸ�M�3Q�F�N��c��
Qg"�@�Lc�H%�@�;�^A]96������ϾR���E�0ΊϠ�4h��.L��a�3�����M2��1�WB0��A�q�*�_�?�%���h���6�
���^��ǀ�@L�N@�_6HW�J&J9gS<�/@古�<�������A{����L:qNh]pl� �	�t�T8�[���m�
~���{WN4=3}c�L=����)�KP󓻇��4xLҌ����VhF���xP��o�J��#:�uc�bc�������Y^�J �1������R�	ʔHZ'ڕ�~�5!���l�{q=��m�p+�~\�M��FU�̗QϠ�2�XgP�u���W2�
RH��F�ח���1X8&�&[�r+�ﳳ���P�u������s(��
��o�m�:��0�_
|�)ų]_��BMO�D��P3I;v��h2���m�u4��'K��>��X�:^oc����G8�j�G�<	vVS�c�٤ˎ�p��Ƅ�3���r9i��]��f��s�}�Ew}O�|�蟜q��e�ve��9"z�%�k��x]>�$�`<dў�Ś��P!lM�]���-8Ѽ[Wa�ޜU��ʣU�ҷ��u��,SR��{%�&+����+�\��S8u��U�2����.�JX>���"C!6'�,ި�hxN�o?#���V4O��Ŭ�;P+>�M."�WZ �輮�A$-+ɔ��������Y<p����X���&����j@�T�Wٻ�@2�jS�и����+D¡��%H:ɪI��&��ď�f�G�8�v"�:DF����� ;�.V��3Ѧ�u��%��V���_g��͛NJ����	������vD��Ps^���m�%������X#��RM	6*�̃3Ed_��a�}��ÔGr��\;H�/����rn�e��7���=r�"�rO"��\���1�a;;����R�,h��l��� I����z��`�h#�F����`��Id���Wm�ӓL,�7U����k1b��;2�!�`M,�[�ߚ�˺B�j�A���� 0<�j9�����m���n�N�^����ٍ/;�QƐ�!j�6kj����ޮ�p-�jǓ���O�3��w���?\�r])I�a�>S�񭨤�7\��P�����A�/�"���g�^�i7p$�b��c4ZX��߁l,�0��?0Z?����̔g]��-�UCQЬA��}V�a�4��8�hT�;�|�D�*��8]`� 8�8\IG;�C�ȥm6e�x%ymt@���+IB��z|J��̇C̉6$X�LCN=~���p)����)���\,)3��/,�X���-�ԟg"9� S	��!xQ ��~`:^<]��1�mIJ�q�觩��u��s[O�H5�@�"[-�g6r6z�T����]vJo�7㋘V���C>��f�h�Ӣ��%���S��g�E"I���m��4\�L��1.�l�Bj> ���u��DS=�դ���>�F!�?�]�Mk���H��FUU�.�����*����������qO�~sⲦ�a*��&x����N�q���ē��|�c����l�XD�dāc���5kY��ac�dv�-[�af%�xJ�k�Y>+^.VM�������b�Z�d���/��ؐ5(
�����</�r��\LȒ�v���}������w8#֣�V����[�PB� ��`z3�<U@�5}n׉5f渆S��:�o?�k壓4��Q$���@����!���[7��#Nb�5���]Խb�⻃��pJ�ݷ"(�k05+����3e��e��z>�/3+VPo���?g��9��D�䢘��q
w��@��s:�0���ӤJ���j	�c�H�Z��,al�T���J׌����{�5�x����k��\��Muψ%��A����<NROa�b����U�̽,Z����a}���/&�SEl���D���}���,x�����QuG\�����.u�{%�P��HtN�C�O����$��'i��g���[&&�Zi���e�jؤ�Y��G���ٶ�s�����f�j��ᖷ&CJ�J��Rقfkiv����'�7~��I+.",o��&�8�=�gdǭg�{���|袞d$=G���a*���<�=�E��y��>���?5Jͳ_T��F�\j�K�hh��b��_�o��or���#�\��i§�pYL��3�U�s  �6��'7���|RLR����)�T<J5딩��B!���=�!�iF�l�Đ��}MC��ʔg�Q�7ð��I������e{����,CV���;I���S�
.�*��=�Nd����q+�~��U�]?���p�>�&oZ�k��ѕcͮV�Eg�X�¬,�1��n`9�Z XP��Ƶ�[�������M�*�W'�M8걈��N��NH+��t�(}�dnrk̥
��iYE��h\
�����ćs(�@��%J�>���8O����bƀ��OWU�}��ξN(�O����#}����>Z^�@�u���9�7c�\�!"s�4��ηNQ�S��m0����R�Q#i�iX����nI���߉?��L�R��P�����M=���1�-|��	�r��^�Qp�FN���\��U,���u�";m՞ٰ�O�~�*	w$�*�E�ؔ������3�z�f�V!D�_Y�>dj�1�(��u��h�ߗ�d#&��p�C6F��ǟ=����})��CR|�Ф?�}3*P�.F�:�H���f彲��w�R��v��xpw�X��<��H"�k�$�y<��7}|6��u8$ 9Q���ԓ�{F�"jl�؊��%��\���� 8:!�_�b�<;�Ec�u�=��hP��w��ހ�܉y��q��,Ӱ9�Ł�-�P�e���0�'˘^�w�@*�q����������Ԯ���*��\˗�aɬ�E	�Ӈ!u��Ӆ���ۊ��>wy�Q�ӒHH�55X�U���6�&���C���dW����a��;�D�-�[��@P�NU��K��O��N��H�ұ�ns�{"V;��ցJk�t�]o!t���5e>�l?�s����MY� J�yϕ��u\2|!����(�pM�Q��]�&R�
hc��/5+*�ܞ�D�AW	�Ʀ��>)��r,���/J�V?9Ҿ��\�IqT�����I~J%�O/�ҍ�_��6��E�t䡺Gf�K>
@*��[L��ۯ̼q>����K�:e�ǅڨ[Ê _�ݻ��tsm��%&2��9"@��������.��(*�F%�2={��n��$��6��z틒�Ħ�+:�|�~�Ң���W M�gn���y��K�4X�Ǿ����j`v��A=�R���i>�`͝ -�1{�5�6j��Ě�V��߭�&��MP!����!��%� �!oe�)wcR����H~��=-ho�o�7�M�� ��SnK�N����O��Z�^k�oG��P��H�c�l�F�&��wN����L�\m��6�.XB��w���>���&lϘ�b��6��T�(�h�P�Q�/R�}��u����f��ŷ��G��UZǤ��t-|N���aM�9ƃC�n�V7��U�������h0gF��$m�e��V�>�-�M�tO$�v���C׾X�~1a����|5g`�~�q�oá�4��7��v��Lq.a��cJ/���etȉޕ@��o*8}�)�g���,ɼb\�]k�౽���1_Hg�?C�}��zm[YeYr,*���V������1_T��e�PV��"cZ���\� �6�����f�0���5|A^����w�bY�G��"���q�ORy�
>�^j���,Ae��>�i�f	A��5���K�����t䷙�u�T�[r�i��`l�\ѳGG%[s$�<��٪�l�q��0Ғ�CO�A�)prb�r��F<Ս��� p�J��|M'3v�h��}����y��QNA��� S��I��S����*��,Y�[��4���u������d��!�����5�}��Pp�=,��rve�T�� ������i�Y�X�[@�y�M��&I+�'�}_)���ѫ`v<�:��A�씒%b:�5�����ĉ��Z�`�~�Ej�2���L��	GG�A�T��fHY���Y��d1���%�9?�q���	��0���sng%/uE�$�6c���O���/���:t���5�&�	��z�`[��<����y�d�w�&3�6/#|�_��aR����X�,���g�v	�[I��1l�<�-��
� ?[��sQ �I[d����J�F��!l���K�`���
�Õ�ۏ$5�Ղ�H?�n��|�3_+�}�A	�lml<k�bu���%ٔP�I�j���<���	br��!���Ҹ�D���BH���*dl��ƀÒé&	J��_�x0( �KI�VY�:�W��U���<�C\�Y��4�>U�-��I	9��+�L�Φd\	[d�Tb�
����6�c�˴)��K��8'1��k���gЛ'u��Q��O�i�b*3����|9�h�嫲�x<�7d��_y7>*������d�f�6���X�&����>ōf���ȓ�X��&��lA׬��g��������s����
i�Q���H��Z�7��4+
����-,�#c�]a��.
�;��M�c��dЭ��h�S��~#���~B�
N�5P�q�e��/M���"��ܻ:��k�CYT�r�bC�!(�hz{*�@&�չԬ��
'B��p�ü��!䮊�L�5<_
¤�)��Ơ�T|^4��W���I_JF�K4�$�>�`e#�z⣙�v�3��#h�y*��'���Սuq�\S�;f.�Wu/�c����!�lYv�HQ+j��v����i�����w�B� ��;�1�(/��K#��E�N��0�V�M��c�u.c��H�	j���Ub	�Ī��L�ݴR��=x0-6���w����gq��{�b�&�}_`I�fWd�TN���j��b�	A
�(ӓL���h�򬭕��OK���bd	�j#S�!oy@�K�*�<���|tb	] q3�=��kd�������8���X���0	��c�	! ���4��_��P���n��\�9��`�GC¢?�D֙����&���>wW�b0�D�44���Y(d��|U��'� ���C���*�D9��'~C��k����G<d���BP�HW�wM?����|�G����&<-򞃡`��/�:��VNg����+�K6�G+�}�K
6��A#ۍyڏ��ΏP�b���#+Yk���F�~f$I�	�o3�!`�_@�E�\ε��������
.��֏s���Η��}��*2� �>�ۓVJeo{!��z/��\5U�LUX�m��u��o����[���6�/���~���{5�\��f�#��i��'������2�����;�-bVH�E!����y�}e�9�+��6�X�'Q+5r�t��S�,m��ݚךu:�1e�q�����)�R��R���j�SA�I}�Wӆ^��1ѥ9~� �* ��";P1��L�?�m��S���c��Ц`X;XU�RS�/�w�2�(�L�<��\�W{ߎih���%�T/�
J�N�p��7e�	2���}�)��W5�E �66L7�B&d�!
jeI�Ϣ:JE��pc;���%8�Գ�!��܆�	�J�(�۝���� ��ν3Ú����>�&<q���������Q���xq+��8��=����y����2��/�\�~���<q��k��o��%%�XYͬ�6\��E`��R�ھ��"��A�Y�d��F�u��]�or"%1�F�C�MKF=7��e�h0&�W���EZMLJ�{��"��ArW�B��P���~��������:,_��S��;���`���Ȉ1-[�l> ����6�
q �QU��_ȏ|�����c��!��[�
~n"� Z�<b�b	�IO��`��Q��f�r����mk�$�Gz��,j��5!2��A�`c�Y�V�����U��<��wVu6�Q�-蝽qAM{�o3�ހ���F,m�`Vӓ��k K��-�a�w�	��.��]�!�x'�4�â�"`-�]���bZF�uv����l+�L����7'~#��w�������$�� ��Q�Q���h$���
�f�qO�x�N񔲬�im�b�':Y���%�;���*~�����K)��Q�D��i���<)�I�	 ȷw^`����,�mEJGR>ՂY&S� <'6��AF`�'	;.��6��U���bk�/9��$(쟸aT���8�x��-����=��L���xt��'=��(*�~$����z$Z����nKe�BSK�#]�q/��e�Oܒ���ʉ�#�YB�:�w0ӯ�UG��tM2��~�g����|g�tV�)�6���������)��xw�������}�R�֮���H����ϑ��E�9a0侇�U����A�/y�јn�3���4+Ł��Ї�n���_�$�1
r�v�G�d=�� �g��:�A��m�gc�!���Wy�I�!��X0�t!k����� ��ɞ�������Uvy�7M�h�w#����s6@��mx��Dg|�cal�>Z1_�|3m8�N�Yt��g�{��f�8c���S9&|ܩ�v�DeȦ��(�ŃQ&a�%{���sd�B�t�R���ojvUWk"�R�U�xbt��X�j�/k�N޳@l�̉쨟EW7�~@m(3sI����!J岽�! t��w|����>��Xֺ���F�l#�*J�0�g"�9��0N���_���D�;�P'h3-;C�]e��1�ڮ=�.+ʒ��v{'�Њ
�:�@eW�.Z�����G`o���Rb��!�3�D��O7�ї;��j�ϲ�I��*(Q>;_w��U����r@E�Cl��koR��������Rjp�w�4)�eq�<wgH��,��K��b	4/�TN�\�W;�E��2�Ӧxtsi�Hv�a�r]�z^����C��.g�J�bR�V�&��I��E
)����&/����XNE13V����bE�2}c{\.Z
=�9E�(ä����
��@+�-�_�,}��c��#�r{�ZyG��j��Ybx��u^�#z�x읅+A���ӣ���s.�&�I�h�zeC��O�B�u��EpU�?�}�Q�ZЕؠ�ͷ�2h/�Ep��w�؆&�)�*�U���D)F���'x��r����s��FM>$Ǣ5l�H�1-�u��ٲ�,@�
k/��^��{��N�?RV�dK�rp �J��+��Zؤ��%I��8�YrWvq���@_T'����B��� �뾘�1�R����P~�a\k��1�)Bօ½Z�3f�*kh�%��{�b^��U���zA�@&c�#��4~��M!�B?��{Y�KF�s�'�pA+,!�u)"ȍk���:6qf:�y�CAU��/��n�^~螁���H�0��ԣ5#Sx�_��N7t_��Ή}f��eeh��rբ{S�o�r ���V��I>�F$h3rk���8ʿ�CEs3_��ՀK����)E��cNV�&V���\z�7�RyL�5ƟÞ�[a��P`�f~if���z|���*h1
	bxgڨ�{DaԬ�N���h"Nzw�	����1��� '�Lze�(���6ΛZ�At�*.<:�<\Uz&y�b�#��˩�;9���ܹN����cz+�?5�����_�j͟$�^�9�����c*��^�;l;�F�ӊ�A�]�X!�Q���=�Ǘ���?�U����b�`�`-'C�1�SŴ���qɁ�=uD�~�cȡ���SI��[͇����}���H-�[9'��t��A�l���u�ڦQ0{�M�=�T��A�P"��M)���S����{dv65$l#��f��{���C�V !����
���C�W�r���u��c^�6��STx���)i�Jy����nI�?D��h��Ы�9�s���%v8()�n��AT,T6��cp�-PؕdIү�^�*����>Q9hm#y���D���K���_P¹#��?"���A_�j��6�S���X$|L,���y��_�ȝ�m3ث��#m���B�$p���,��C��zKt@���)�"�M��J�,r��+[ჭ�����D�����w�,�������k7,9�7�3���������T��`Q����Q�%"��.�~��b����0N��~g8\��0��wrT4���a$-|[�����Ή�wu[:�|�U�A�gK)Zu.���Z�ɤd� �춓�VF���EvY:v�3%ys��u��sb�j�oq�,�#��X-�e���Iٷ�O�Y2��� :�~��?Q'=c�+ `�u^d�5N�5��Y��A2h@^}T/d���<��n4Q�����Õ���g�L��q���ԥ��p�ޖ�֌�8��?�.�S����k6��[�"����������x�c�ۑ�]R�T�d	���S݄�]����Uf<ՕY��V���AN�S��IҼ��>�V.3o�,���d���j��Y�tnQ�	��]I�p-�Ӡ�	�u���#���4T3A]葹-s����"Rh%�rT�Yy+8����V�Y���峓�
�&vgw��� �k���;q�<=T�+Ͻ	i�>n�Ȝ5n���e��%����O �q����a��dU�� 5`�66���Y
Y�=��WF�t�י�+�%'�.>�2�#-W$�{�^1�{��0�j���!������o�;���LKLj�%̧�1<�%Y��C6#�롛;T���]�ƱL�/d߽a��}�*0߳�R�xK�~^���Ί����U���S3ҫ�9�֙�g}]l�#E��3���-t��R[���eNJ0n��8h1ѐ���zz�8��kT`��?VI�a�e�u�n�.cW�E�B
�
� ��a���,����M����*�uPc�[�����?�T%�w��&�E{�S��iC�K�����j$8t�j�?1�4���DЕ>U4��Ԃ[�l�� ������5�%׻
�� �"��*^�B����s�A-��?��1��!y3>�-�Y�'A�NR�����_&�S۰�)	�.<t��l޹.z���(r3����1���=e�.Ԇ���>IB����o�3~��[���#�yDp��1�nX���ݫ_��kI�y���G\9��g����@VB��̔hL���*��\_k�Ӧ3�f�Tu�������"fT^�oE[�`,���^�#N���.���0-�RP+���u��'�O��a��,�����T�����q-��Sy�C�ǾR$��+>���f*�e���q�����a��g��0��M/�ct�6�Ki�<����=��-�ٹ�筏5̦!��y;�G�ƼC��YW�O 2�>��
��	n>	��)�-FW��>�l.�DBb����Z�>��U�#�������W(�҆~�?R%^���#���\���7��,d�V�Y����ն�y�ɪ���}vDa>'�<�*�f9���)(9��<�y"�#��&U�ه�).�݇˛C����:�=��5��Gh�XW%;���YEQq0/��hg V����w��O��"�;���%H/�7�qE��V���Y�`� λYS���0wt��$��L��F�^{��>G�2�MD.�)(l�VE��$q\�����Z�������
_�'��7x��1�Ynҩ���w��#�����
�*�J�cc�[��]{���hD�[U{T���)�}P�5j�H���,�@�[��h�k�)=��:��v�#4����,]?h]c���⴮Z��U�^����9���e��є��t��a�د�"�(HMYz�����a$�LbEՆ	��/Bt|���q��޺��w-�D.6;{��;5|���q�̱$Իs\�b�愉�"e�%`I>G$�N"�����(}(�^���O�m��Z�:3�b�i�v:Y��[�w�f_|gb>��R����C�Qʏ�����H�\vy���S�
t5$��*�iN�_s�xX4�r����릍��ɕ��������C����mH�٬�v4d�lC�웫�'�[��V��.�%����T �ȯ���@*B^r�BltF��1o�����Z_��q�����0��lb���,K����Nbk�����"6C@����-6�+8�:�/*n �TRy���x� ���}z����	��R)%��H9��8���Eib�<֔<%i��7�^�A��sv`�΃;����o�U�!�J�൥��~1p��4�	������T�ƿX�b��fH�t����I��/MJmDߑh�'�������bi�b=E��ޙ�k���G^�딇������v)��͚.h�V�`���VE(H*�;1`Yy}�L�e�8Y�e9/��2�V���#C��H�6K���;1��}��p��2�� ����Izw� �����P�w;=b*���U{|ܧC\
�N�rը�5���gdW��O�9I�'��=/@ʗ���)�`����N
%�ݳ��ێ���Dn�ʢ���ȃ%p)>f'�����h˭��ȟ	&+�|�+Z]f��||e�B�J�ŪH@u�����g�F��0����\yFKOlh�-ٻW���4	"hnS�7�Io{�JĿ�l�m��ז����t20�~)�C��,Я���zݷ�O��h�ˈkD�Q��s�U�y�h���I1D�E�t�xq�2Q��B]��E�aVU�U]ׅ�,hV:4p�Vf1`�-.).�oN%&"��!#����k�h3�`�o�q����}�f�iR
zTZC��<^�2�A�e+��+B�ֻ#���::7@�S��7:V����z���n�
w�6�VHx��G�����
^��g�-�b1��v1����J���y}J�-���W�;�uK��P=��3&k���^JG�2�˟���y��	�QI�,���*���_���:���H���IG��=�����*5���-d��S���u�mA����Y��!S��O_.U1 �#�E%h߄leW-ln�YR���d{˩�"�3\T`M[��"�	ո��L��%XtSqdT�n�EroT��Q�&=��P����`�jС<[��"C�濢�&\� _����N��pRF���T�ȁ[�'��b����<�C�&F���c7]Az�wFns��b%��p[~e���v>8jVzhLi�~L`�זPƃ���j�W�M��c�`T�'epɶ�N<����\�2��IX�A�h-{�w�6V/�5U��\���U�Jo���?�B�Kew�����ܚ�c6�e�ӐJ�;f�ݣv�i�)�#J�X�%\�I��+J����b��X�K�g�T�J8���%w��`O��\ͅ�h��V#����'�O����� B�X�u`H�Μ���jhIEk�����"�P�E���</�l�mݵxa�Åm0�v�}��J(]�rn����R��ۛ%Fs����r�H��s�����ZγQKA:@���ΣAu	w?.t��zS>����������F?��e��/��*�
w�7;��z�S?����(�X1^W��9M�?S�����v�ޔ�}��<�q�)XN���d�KA��iw��0���(�;��B�J���5�t9O�.��B�<F��4��"_�_6o�����p�Re��|\�?���e"�Ɋ��!o'�o�5��m�h�'l������~��:��"R��̭~��c�z�]�?��USDy
�O����?��r/��o�2 &?���\�bs5�N�F��=%�0�V8_wޥ��~Z�]���6H/�k�h�CZ*�����42\��L/j/�]W	g�_W�엀3�R�_)���Rg��������͓5g�yh}4����\E�~�{�&Y���9G������#���M����ly�D��>I%_]l&�������E����=�L��o����׸�9�Rzg��ܴ0�Lm���W�@�
C�����/x["��Hsg�|�۲�46�
Pћ�Xd���KͩP�.ݜ	Y2{Y�b?0��J�����<��z]X̔���&�d�5�`��·�#����68&�A�;�����ixLգ���I��7߹F���s��R�*y
�Zu�}v� � �!j��eu=t5��[�B �R�� }p� �=<iK�W(?ك�Ru�{���U��o�N�D��s����c?z�6\5[��Pd[H��]j��uч�cV!�g�#l_���񽞘�`���$��^�(�����`��ebAU�����ިb�WwAqY�*�TL@ؓ��"�?���%���)���$*���J�uf��|���xb���_+ 	IR���i���t���@�Bgf&����f'f�=���Wm&m��=��
�EJ�Xc�C3oT���w��n$;�����H���*�������r漎����a�qk}A{�'v�4�F� ��('0*Bͻ�� ���/�,�F"�8�t�]J�J$��_}���C���/bZ�!Sۍ������Iv	H��өDo`BT����>I8f�5�� I�Lg=�gt`
�� q�|ޜtR�����5��n��؝Gy�?yav���w���\��V�O��	��x������띄n��7�K�ԕY�6�*�(��u7[<٭�x�J�~�eVԲ��L���y�uPd��GJ���>��y��������0"�*�=}�苐Q��O�N�j�:6�*ڸPµ�� �W=R�X��|6������MM�+��7s�^����/&Z��)(��3-F�	�/{}&�⭷~Lx˾����6>�9r�~S��>	���o��#��L:ȷ[	I_G���0��j�NA���-�	������]�������P�ܘ
�������V:au1ﰭ�\����"���n��A$���5@�룯��������oD�ٜ�-���G<��(	���xtL&pϮ�l>�x$�Z"��8�a��u��rboJ���?W�B���xԒybП{���m�Kb�^Z9|�Ü�c����^�їC���wn1��h�M~.>�EzK�P����49א�^b��L[h$��qQ^b�K_y�0���\�_g�G���uϩ2��4�=z����Svk^��Ut�Z]Y����K��?����Ϫ�`]���m�	�W1u�$*V�`]��jgS�N��i��/�'�)�~��=8\�#�q�H ~٦?�H���D�;��q�@դ�a&:Z��:~���f�N^�e�H!���������-ŷ��¸�g)K_`]%'USJ*+��mN;2�cp�����"�.>k"�nG���}���R���=�Zj'W `�� ri�j�E������f�p8&92����F`���j#��t���γ��7/���|˴����|b�cv	*-��,�y:z�РU�5��xb5]m�B�^�b�|u����dUя�����o)O�H�
I�e�u>�~~ۺ�+`�VI���C�`�����J�x�jYʰ��?~�!���}���!W�ꄿE�~�'L����^r�,b�k��O�J��኿I�&����`0�W�s�w-j��Sk��冪�e�c[;�7�{�\�����4�WV4��
ma���p����npZ�趃�Ъz�����"-���B�$o�2�B�%�@o��Q�^U`�`���̀OKz�uz!45��;�=~��Ɠ2�Y��_ȍ��%zpf��4�(��A�Ys;����h^��@����� ��f)
~a��p��t���=�tQ���j��k{5��j�b�oY2x�Ԇ'�n�����*OJ{�!m�i������7�*�S�
��i��2�ƣ���1_���j����uV���KQ���2h��&[�fw�-��)���]�����
&���>1�ONv��EZ $	����3"$�]a��:�XH�����@+$��\{���Y�_Md���B�K�M����3K�料�#=�˯��\��g�.���h�����R[�7
�G��ZxqR׵��R`;|W7�B��t��bAu�ߛ���y_�%��,�T�#K.�^��!�#�X��
�m�H�g�VW@�a櫐{�q<P\�*�}9�W�����2�=h����a'�NdM���.|�ӻ�ćZ�>=WR�eP�(ŧ�N���@�u�O:������$l�袤}%�|!tgw�����w1�-Ǐx׫=+i�]_,����sI5:�G�k���A�ⲵ����{�>�eBAm�4�#�L�֖yT�z�����dK��y� ������3���kf�q m�
HL˭��"@ �-YTy"��~c��!1�ȵ�e��4,^e������K G����Õ#¡#O�!�c�ډ�X�62
�(0��IWhѝJ��SQ���զ-n.�,���5�d��\��ط�a��B��9cs�I;1�?����_]��YtHs�Bmq+K��iF�l�����2�~��Ɲx�����@h PI�]korus�q�V!O�'�rp�LxH	��ש�����URF9����X�L�C��Y�Og�c�&V�FXŔTеǻn]����Z_�\�ZD��az�lJ7�϶��G���_��4ab����Jq��6?-�9���ִ��1�)�&��h6���qN'�q,����rCL����:sJ���ce��%x����M�&,咾(�7kG#-07[
�"�m�v��
�f��&S`�qW������SUkuC�nl?-�{ɰ��86���z�f�y'����0��袗�M�b�z�C|���,��T���J�L�z��):a��1e���_�
.��*��I�;M�DGæ��S�����``3��7ƕ�)��s�<)D���O�ٓ.\������~�.'P�Hb��M���5qnD���k,}#V\�z���F���^`hzW6#Wt�ը�_��c�5�T$h	��GmN㜊Qr)Ds����x��M����b-�C$�Օ�]3�>1+�XE�q3d>����%*}��+��G$�m�-�K����'I���Ӣ�L&���<��a�|��/^�^^��{ͼ ~���&  B�ͦ<��e*-qI��Y�3�u\{AE�3�'e[����Kr�\-�� w9�ݮe�6�[���b���IRn�������jp*�=2"3»D;�"���1kjv`f��x��R�WD���u[P٨���O��7rÈѰ���u��UP#���y��G7�%KK�H�_k��lፚ���]ٳ�E����KF̙Aʲ����6�Lՙ���E�jWkG�m7�gR��w��K��&+Z����އ呯y��\N~_���u����gs��C{�h�@�O������Q����k�_b�,��-�)����ӂf۔)����ͷ�:�O2�bHp�)���+2N$u2��>΄dg�=���Żݒ��u�߹�e[��#���ɖ�2�BBXYe�����n�Fs���>��2�.\`Ȯ�Y$�U�݀m���b1MM���c���/�,�8�Ol�c6*I�l��f�>��Qj��ڤI�8Z�pz���y�{���e�o�C.�D���&Ҝ�H��q�	�_ݱ����6�wC��S⥅��	'�
a�i�.���;_n|Dn��<�D�J�̨{9��,�43
��+ޟ�/���!bI��"vE�0�Q����%��� ��qt���޷ $eN�Z3���!�|:��Mlld��N��I�-lԴ11hri�B��̸J�b��i��(�Fa��y���TM�f\q����A��Ύz�[�9���=1ġ�{IR,���.Ү�q��;�l!!�_�Ǯv�*�p�!j���WT��2��,w�\�B��N������g�/&�d_9�S�\(�W��RVu����>B�e��H
��^��_=yj��]�[�>��v�f�W��x� [-B�L���c�2p�w��l��d���*Ĵ ?W)�i��f��ܤ��SBZ[Bi�j����m��J�D���_h�>����O5Z-G�:�<!�A ��"�"G�o?�e��M6�ȅ�����Ě���	����ͰN74���d�/g�fy�ˬ��;�xBU�"I��;b��X��Fq�>�%(D�	���A�D���wI��� ���ə�\���<����faR�Ǆ[�6������j%�g	�M�V\�G����m��A{�͞~��5@��Y��A��:[g8�0z�7�yb��%���P4^�iO�p�!x��7�'��ifb���ܺy����*���Ԏ?IpQ�a�����e��G.����hk��Q9�QcR˞*�.^Q�����;��D�.��a$���S\aqE���N�%�67V�z44u�=h,�Y�3,��6�4�/��@�3�[$��1�D����
��e!-#��y9�ޅ�n�ʅ礧
���V>��6�'N|�A��I�k�� ��C����ЎN���&�J�f�n�K����DW���I�ouh��p�,������i/&�;�
.Z��Ij��r�8h��1c�YR8W�QHP����W %�,�DZ�߈��i%O�v>Ȧ$���li��gN�C�����_hUP�ߔ{>�u D��6 �=��{�E҄LFו+�*��d}/c
���	E�ZG���}��\�r�|x0��ٓf�$�86Ȇ���|�h8LF��`�c��S��� �Z꼴�3����1]*�B���'�d7����q�&����Z����z��Gx�ŋO�����u�<y�!]E^�ؼl+3U�J#,��c�I����{7��oJ�=j{AM�(b��xk �x]��׺+��%_AÛ��h��bM�_�!��v�C�'n2��"��e�'w�u���� ڋ�8�M�vKo1I�;��^qU&$���d}�PnX(?4'f�LP]Z�����@貦��*J1l��T�����S�Ieae���	�?+�X�)���w�����\��@B�O:?.��ӈ�6ϡ&���<�r���IT?�r���eh��j�"�^lvY��*1uuV��]�i"��xGa��g�B*�����|�:�^����5���S4�i˂i����H��i>�E..��h��OP@�5�(�W���9s��w��� 4C;8��F��࢑�b�S�*7�\��@I@dL]8���\j-_�p���f>�ntA�@3��t\��J�����oE D�������6�)͓�Y�{��C�H�Q6'pv#������B��T�E�vj�Cd'\i#`-�m���B���z.�޸�:~Nj��QB^4�D�\�;��t���D��K���76���t
ʸ�Ė��B���	�a�I���҆��>�aQ���]5 	�3���<�O0��n��  ڕX���֘�&�>:Q�+�DM��.=�[�D;�t?��or��Y�{�4���%ǝg(�%!59��Lc����OQ+����c�κ��'"E�'��<N�[d���T$@[�RO����.�f�F�d��sk��CV���@�v#��q��ُ(�ho�ÿ�=�2��!�\eOȵ�i:�O;���w���;���W�޼}7:r
�{ >�6�Ԍ�tҧ7\���@Ω�Ř�du�U�����V��J7[�IԾ��*@��J�k�z�� ��=J�������\r�/嬘lDp��ڴX����+O(��g� �Wh�� �W��]��J���f�ѺHЋ�Zݣ�rSھ��?�ָ�c�Ue&�Le	II�L�^4�WA��IPlr��z�-�C1��a ������yg���F�k��o��h��恸|�#�?�e|�������<�=��[��b���`�+j���vu-�,��:��8�C��l��_��\|�����\ࢁl��J�ӕ�B�&���z���D�ۏQ]S�+h��TWt�&��Jv�����A�z�V�o�hF>7��_�e��t	򣥇�Iڸm R��AT�d���d�s��O�*V_���
�&�fOʰ�;*ļ��G'9YXwCf�*����dĻN'@@f���͞�%����ȩ�����;U���������s�Pj<�G���c�W�#����JIO�i�[E��N��w�&I|-Ex�x�~[>��u��%�&aBˋ�"�4�M�5���cſہ�A9�}��H2~�w?�C禖nfOX�q\��pR�Z��?��!{_���$�]d��Jt
Α����UG��S������0����#�H��(��o��F��tEny��e�b�kQ���ܖ�K�X�\I��I�<�f��-�-D�k��d�)w�/���4y���v|�A�E+��e{���J�T�^����4�� 3c�h;���S�� �)�ق7�͈h] ����n=�&{�s2�X��X2�~��ժ�}�K}�F�+�S�̏�r�4��E�,D/�z��`7��,�@b�:D�G��Z�ȋ~jg
���k�/�9WbE��s������Ѥ�xF�.S�����2XN׫̧@W/����T���%l>�����n>{W	Cנb�w��<�xc�0ʜ�����r��ݸ<gw�S$���I::I�]�*��7s�Y�1M���gi�H+a5��F���h��&�i���t���">�W9��$M_�i��f���|x�G��n���3)�E����t���{:�?}��B�O���dl����ߏ�9�hG^yӹ��Z�nj���N"�����oO��V�r�|�9/GQ�n�����u�rl.������1�;��}�}Ҍ�o:*Zh�e��x�2R,���0/�/��!��#�-c��_�QUF5��޹_��?����ьq��E�A1� _�r� ��yd�p�����1m��fq��Ρ�A1���P�b�:�ڔb߰��w�D�T��
��")Zŗ"S
�ۢ�p�-�SIL��_&��LV^�ѭ��Y��6y��a}��5P��;�)aY��Z�̠s19�҈�U��g
v8Yi�t{o���0ֳ<+XR��c<�\]���lF	m��?jUa\�
��(�qNDX�v���%!����6oL�jG�ȷ)�PF�b���J��S+q��7nY����6؝�M��(�;I���R0R�;��xL�?����25x�/����|�ܴ�U')�#e]n/�� f� u�Y�x��zƍ].��jb#x��'iC��g�����wd��c���F�׸�GD�Q0�x��q��{�U4��006�Gr�u�������	�5	_>3ĩ��/���BG5F�E���tͮĀ{P���+"�ʓ4���2��.���r� ����[�@G�����g���)J[�3�I�(�d �NR� G�������O��d��.<�{���?�mbZ������)9���E]U�_ai�Yi���Z�������y$BPP ��Ɵ9��u��L1�K	��Z�Xk�{졹��ΔbR���������1�+���LcJ+�#�y2��]:Y1���`MwG�=�&���nZ���(�s&^�r��QZ͋�+<|%�}�2k+�;nG��CG�W<�P�M(n�u!U�7��y���1�L�ؿ����3v�e��˙%w�չ���9�s�C�VɃaLH�P�-�RY���5�o���������.�:?�8����r煇�-ؠ�ب�Fڇw:Q��H���)(0=a��F;/�!�j/��k�J�v�i���R}�	���]���:׏�GZ�SP)����<�S�c {0�����A��1�Wlڧ�PV�z��.	���ǂ��"�<��ϕ��eF�l/�����]��Nsuܱ�l8�wOWGX�@�>�-��Z6�%�P��b��J�
z$�����#_ιQ�eZN������>����/��#�+�:���Q\q�}}�I31��eR�ХR�i�TX�Y�����k�c�Bv;E�[f��'rFb��hEH���m�A#� �E- b�;��%h���v	%-l�߼H�ڐ䳪aEl`YbBQ������h�v2�!��j���-'GRZ@DyW�?�����z &��D��'7l*�_�7��|��ݕ&*_��A���	I�A������tg���;y5J{������iX�X.�S/$�� R�gNnt-�J(`� �ԲL���f�D~U�K�z)�T������+���
5�&��������K������6#�dK�;��a���}+��7&"�r���w{�T�� ����{&�[�m�������W�o�bb��W.rQҤ�O���o>��Eë;V��������Iy��
��H�!�dﻑ,��E2i��@�%p��N
�!G���~@��_�[&��1B`��]�6'��Q��#�_���<`5.+W�_J�k������]@%)�8�Us(j?Xv�,�(��ɾ��-Ek<�:%����p!��y+7C��̧��Y�P�ё�uJ�(�@��5��L���Ү�k�bu�Iu-tr�X�\jP�S���m�ڀ'�c�]�7��C�}��a`�6��6���`.������E��#�-έ�v����MjL�:5C1�Oa�o="�N�z�����
���f�{u\�(��4������'��2f��O�"X�>e�X7�N�{q�_��?T�G��SF�uTh@��6���@J�@u�ݒ�I�Ԣ�t�a��g��D
r��f>�\��"+aLj�����3�\x�P�;`R��"�˲�l���ğ/Ѯ�0�V@Ṷ���^��H�6�Fq�.��V�1&X*��'S�g�Z��B�SC2�|��/h���?���BrJ��
�}�v�g�F58ֆ[^�WȾJ���r(���,.��l:&���:s����i�ĭP;`ȯ�-��ԟ����T�v$���5IB�M���X�S����L���mn��U�c�Z����� �f��x2�g-,��=6=S� ����d��u���<܍U*�X0�[]�;?�!3��a6������ÀQ�y���9�}��d�lt#]����RP��>���1
�����$(u0��J%Qt��SJ*�S G��*�d�A#G�	].�i-����b�CRx��D�hM�l�t=)\��)��҅�N��}jA��)}i�����.�ߊ2���yD�}BQr#r���Z����Pz�6YS��j�l��;B
T�c<mY/Tf��YG'�8q>�α�W���#""�e��"�Im1�q���"i�xS�G ���"x��J3�>�A��a���EJ����å��cSB�����'�jh��[Xp$2$�8^��Z2c<T��A��+6��dC�4R��Jua�P��n	%�V�h�S^��_ƻce���&�,��_M��!�b�"��"zN>�X�HO�J����Z�qq�8e")�-�ג=UY��o��[���Y�wp�B�-�7<��P�T0U:��=��
"��"(��f񇮞�j(9�rTzx$�N��0A�l';ש_�4=\=��@:�(�\�+�Z����Ѹ��(�7FR���1�#�߆�V^fǉ2S�(��䮺"E�z뗠��4-Q��ћ`����$H��Щh�E�{�L�p�x�0�����ãM�	&���F���N��(���-�o/�$�}�s�=�����ٵXO��ٱG�`���}���������S��	��w��7_[�BB��Ѕ��!������n��B��x�����2�=R+^�'���߈�^?���i���4ٜ�x��S�I�]�̛��#����~A�
0���%��e/��s�-��$���o��7adiQ���vs�$߫A�E�j8�&of7��NI}3�5+����}X����'��Y*�<�lɻCtOB�a����63�5�i�������k�S��TL\��]���V��x�IϷh��c<����{�*�(��]���}��}��)�G�ߠD�y���92�a���SJ���!u����+l&%�bā�0����@��#J�OѾP"�N�ΰ�D���݋т9�JQ X
��	����,��6F�?�Dlw�:��x�:[�`�-K�F�~~��B�L{�_W�n����j�$���`�F���?q�x8���bO��ʜ���Ŵ��*"���V6F`�<����$�\���U�m�?��m��6�U2�U���`�PK����XX$?)������!���v�^ZV/�g�)*ZL����B��܎�1R�u��st���~�eJ�j�%p��|:�U���AvX���r�"��Ct�b��ysW#0�d�sFg���Ӊf�`��'�ĕIFi��AC��xx�m�	.G���m>���[y�D�hoU-���:]As�|�N؄��{�De�Y�gnH�=�|��ȠN2� $Dߡ��~�o/_:w-nY�g�����,m�O�����'N+?���g{�6-��Dc[5��n���
����~Ջ<�R��{:ckA�Ǣ���S1�'�	S6�=����>��o���{&���e�3���<�����&��cŏ�G��:��� W��_]|�֘�+d�M1m��}^x���)�˚%=��gusvZ~�Vm�r�d����é�%#�M���i�W����A���=� �/3���[�5t�XZ� �KRh�d�S+0������EW�43�e��q�I������B�Q��]b(<��i��ZTJ^n��U~�����g�3P��7��ϭ��.� s����1�6P(&*� ��oE�H���\x���ț�ڰc�5d%��Ψ��N��JŜ�ވ���^���$]��e��NDXcQ-��[Z��i��\��t��M������dO��=��ȢQ��s�����WnfKi蠧����ǝ��[����y9�P~�=�����k
�� �{� u�BX2��LC�Ow�~d��J�b�	�;�pF�::Z ���B���'v5�z���<I�������7q��c�NI'�[U���%��'Buq����SD�ݓ�!�=�2U|a0�)�ofDf��C����i���E�m�L��o�h�A#��G����c0\xw?��K��BKfJ�/y������d�_HC�J~���_���$b��O���ã(�yLt�Alć�+�&�7%=�,�i�D��6	���$4�*F&��7�*L(ۅ�s*
��t���2¬� D�S!c2ت�^�����>�����s��ٳ�A�$�����x�y+����&�$�y��~{��&�4�=�� �z��BoŘ�����Z*�|.�z1�Wjބ���Cըi������������:<�z%��0�r�DSB�s��n�������7����ɹ�t��;�r=�mg���{�%���9k���w���]9ϳ�A��k9��(���m�C�C�'�F�o�dG����u�Ÿ���?}U`ຸ�E��K=��9-_&���=�lT�� ���'��,�L�k|�|.T6�lk�F�P�Y5��@�ԧ�e'h^�2}�|b��On�|��WU�%�eIw� �~eK~��Ʉd���ӺB�gʩQ*�JAD�֒_`� ���{�$��w�l�iEθ.v�����g��#
%/�}��2b�����p��������Q�>߲]媡+�m,1���I=���"u�dK� �ޤ���3�	|��L����?.�����5��}�;Ⱥ������{���T���鈟�
"��(���6���.�a���a�Ϝ^��W:�2����ɥ&����9�ۻ�4��B��8����0��� ��ܯO��� �C��ol%� ���p�b��o�Pe��Ô���"[wg�'�Ue)8�%�;?����DO똋����fG�_L/
�C�by�XgQ1�� Ÿ�ڠ�&?9���Nh`jbl�8�P:��l�R���W�!q��G�Q�2���,��T���؀����{�VM@Q�G����@%7��v���Z��D�z?2=�Y�dJP�&��ڊ�Ca�,���yl��M�7X�J���g`K��v�~+�c�<j`ɏ�y�����Y�tӜ�)]�)�L�gɣ�����-�qH��"�7�||hډ�z�\��9xJ�VLg��1���DH�$���O�����m��0	��źd�W��Xnv�'�2�40ޡ�E*hW�~�d�������W��ٌ�BY�����#X��[�mr5�e?'��]�M���W�hZӄ� ��є%d!¦�;K"��9A�峝#�{�	��[(��3��a],r�E���<����<����i?B��JCk��B�A;Vgq&�D̥�G�����FM��B2}��f�p+
h�떺�2�����@��c��}������Pb�m5��)](���ʫ3��z[s�k�T�8jfٿ�����V������r�!@=ǳ�	�ZJ0��y�޶�Z�|������)d�}a�����$��<|� ˖�I�b�cl�Q2��{�79�]���I%��%N�ۈ�	�#O�s����&r���E<y�oo#ك29�w��p�Zqx�%����&��*Ȧ5j�j�W(/�P�nB�iF�mU7p�:8��%�H��l-]wZ�'3e B��o����R�V�"I��9���_]K&�VFb���Rt�]%MS���f5;����8�q(Ve�rTRI��^ W�g���/[��g�:E�G7�'�Z�iY9��xf߭�>��{�\���|�J��''�{
��״�1��]قv�ۿgdH[T�4ȓ���#�u�T�ǞR��,����\!ݭ����9�=pȾ����W���3U�/Z)��[����K?C��a^)�j�S"U��F�N�k͌����ڠHHŁ�E�vnn��aCo�T�"t4�xPd���j��+g_[8��jI@����l�NԂ������xdO�����L��d]���%������������;AC�f|�-*)�(�� ;m�� l<SImk�=1�uq�򺉀+=s�< ��wlFer�~�#�;Ӗ�H^���U!�=x�8���dL�)����a���.VB�v�FH�6��R"�<�=?1�*�G��O�i��M�	����ɋ�jz�(�jKg����|5��jd�� Zm ������&ʢ�����6Z߳���a�����)��� �z�XG�*N�kE�ǆw�ԋu��n�I��r�'pSR�� ����˷�M������KM~�W0Dyl���|}#Ú@�8?�04VNXq����U��>ɂ�MzG��6�Љv8j�_�Ȋ�F���}߅��u�d��*d����h��,O%�H�g�NHpW��m�9?K��h_@��h��./��&<�h��R|0@���{٭�����|!}�c�Ţ9U�傯!��|�jd
�����|�omP�\�%7�p��ٷ��モ|����DQW{������ֆ|ݶ'Y`̀*~ڢ�cC������V���]���R�O�n�˛����#!R������\��Xٶu�����u'M!WH�<�L�s��JB�m�,��ep�Bd��jh�|#*���sOϰKd������͈MV�dL�0��ڭ�~�����4���3�f��5�^����U�����8%���l��$�-�^�a6���5�I�����QJ�zW��G ?
!Q'xcgɱEl'�����g؈aG��OF6g�a��Y��녆�E356Xd�g��9��o{g�!�␊�_���Z� ^ E��<���̪EJ��H
��ӹj$Ѽ��^��&�I�z��f�\uM����y&�7�8�t�=s�g���<uh9H[�KG��q��F��3L3�bE�B��Il�"D���2Ҡ����B�	F�zf� �4���_k�'! �p�0u�z*7H�hb�̽��I�u���U�F�/��?I��2��BE���FsV�';P���@�s}���)�z��E��� � ���2:-ن�^=ae=�1䗽�VK�YH��4��&.�Ek�T��v�6dM��ZZ;���ϲ��N�@>H�\u�n�`�戟ŵȌI�G�|�gk��rq"�N�P���/�kp����� �[&=	G���w���Cz��'���O���1��&4�%��,����F��6�m���(�!��98X�Kavn�(WW'2�Wv�mb�ݨ6w�Ѥ��Ln7�B*1"b��W�V��w��su���c��x	(�q����$7\��B�X'+o��,���Z
Z��`d�Z�"�/EU9&s�f��Oh�Q<w�R�/��D���҃&"�7 �ԊK9��)������� /^a-}"D���2-|�iS��x7�<�HŖ�x���t쯳���@�Se��]$q�hw�>��A��DF��ד_$�x �Ļ�"���#�WB��^&��/h�f��=�-c���$��[$�9�;�k����n|</e/u]�ǭt�ﱗ��"I���F�?7���a��v�?T<�V8�����ʄ��`[(*>o�O�2����H�zبC��^�_�7i����5XI���nu����"�P�� ݓHU�,�j2[�cڽl��w`x�ߐ����Rke{#��\����8i��tSGҧ�@�O68�sZ;:����"�GC��hgu񏮖�YP	�#�
�C����u(Ul����=4h�OQ��벜��ϧv�]IkW�� �8�� kM�uA�7YD�j|lg��V8w�Ae�;k�)h*E�tf�l���I�m=����K/KUT�T�2�&��_'o�݀G�f)��1Nr�l��~V��UGa�˃yG�����qж.��D��ih���Q��������v�9X6��!�ǩ�$��u���r|�#7�����/0�Yf}V��PC������z�NǮ���/x��&H��>�
��&�ylR|�׉�k�p�<�j��
̌I�|���]<�PV��ox �qVc�O���g��<���4Ԗ�M_�,x����,,��?J�-�&��b��[℆6ˈ6nCN��Q�m��MD3k�j����
��l̽1$
�'�"��!�aN���yZ媶�V47��O����Cy��&s�Mu��s��T|
!���AѰ��8�S���I�����GJ5i�ԋ��U'�"kIJJQ[�n����o3��`�K�H�����)��\���,��P��B�x@J*$7�ǻ+�������(8D�������r��u7�̖R:cR�:~�~�hN�k�2��9��( �$2�c>� AG<��:���a'�L�g�B��鄑�-�v��DYPT~�|�T}����G�����;���"T��L����./@�^�c���.��.s�*Y�.��[elu�����s7��zUt��A� ��4��cc7�YYr/�ݩ>lv��=}r���{7u��i�Ԝ�'}
h͂�EK
��oV`I#���L?������$T��C�͡��+rt4�e�U��������J�6��P���04�s�����`>��}�/�2̵C��O'�lA� ��#�T��2�2�no�c.��޹5;��*�P�Y�t�\�U������D1�-����V�<㪤T�!�/��Q���v�9��U�*K{��S�1&�
G����u\��q�3;)����u&�0y��Җ���UܹB��� (�N�O�9�p�q�A�QhD��3is�K�)ɇ�N�t��tܶ���;h��L��d�q�J�K~K�=0!9�LG���C!���D��\:DBa�����QXITb�
��²Cx$�1�@U�0Y었�������\��OL�1��.�w�ȌMS���k���ֺ,/O�m*`���f?���f�����]x�F�@)�8"od�t�~Ϡ߂�Uj�`�<K���i��L�Y��H�֨8_ ���p�܇�k��<�Y�j!:���y�2�� :�a���	����J��L��Z���,?
�C��=;�y,��ͱp�� ��b}��R�&�W�Y,���oѡ�,h�U�FN@X��26~��c~y����f/����L�����z0dF���|��R�g�or�e*wouQ��#�[J�Um�b6��j4]+����>j ���.H�����=���U;e��bt����s3O�6��fT<��64���T��2�~� �I\!Z�-� 3�(�� ~�$�A��#�8S9~!;2�����0B�f���o`����G(ӥ��`|������u��6QЌ�=�ƀ��qok�w�.w��	������%˘(G���laUm`q���PPR>�����y�-֎���S�$���%���cc�$%�	��vy�g�����x=@@�Q�����]�ӫ���U��Woe]��b�̷
��p��`����ca�����M��x���'e�x�m�����<^奒-J�e���Z5?4l��Uk/�O3����J �9y�^���m��v����׮�AK&�g�\v>��C`�3���t����6��	�3�ɚ�u�%\��3'����ib��*�շ2�[��,��'��a��=˷1�`�|�N�W����
�8p���	-�Y�����vhu+^�I�Pd+�۠�J��S�����e��-F�y�TY��6���/�!��A�h��#���c���8kMGN��,9m�B:�P��8�q�#�4�%(��}z��t?���g0͡e����&���!�LMr�Oq��4/G�-�H�i�}=[��5FJ�+�<�@tYt\S����@���j�'t	����:f��s��
��d�,������q��ۺ�#�C�Y�;wr�.�����	�!)�Z��s�?Ŧ�RPU44��7����Q�ͤYÙ���=CFG3�~�b���H�V�%Z.@�r�dE}"���"����D�:�_��LД��u�)�y4��OP<Gs#:�\6�QA2V:'��xR(�ݑ`�;�ґ$�|�f(��ʣ��[V�� 4����<pf���+^�7_A~��~ G[�m������s^!%��sE�V*O��V��]���ӛfKX7���jEO��#�N�f':,�o�A�="U�6K!��'V�^�� ��M�MT*�ơ+̓�������;p�`�X�ۯ'K0>6MCEg����[�a�,w��ķ���}a=�/F�q��;9��4}�!�\��F�]�a���揩�k�}�6y���IiQ�{�0)�Zɝ@3�ϻK�jv-x*�ܔ�O�mZ+z���2�<���:���0V�<��E���&�e_5�6ۘ�Sq�Bkm:E�S��qO��`��o����<��(.I��9��&A�t-
�mp��%K�Aq�ün��a�͔�>ӄ;w�~���*�Sg��0,���`� �T���:��<�R����M����K=8���l�9ǐ��x$C͖��3;����1��'`�Q{��b����"gv{��ߡ�#R�� �[�t�<���('�y.�����zpr� {�6�f��䩫�C�6�������f5����,��(l��-��j�h���p��b��
�p[2|#z��DO��[ۓ���5;�\�d���.xOVPQ�P�`2J;�� /w�86����7�s���O����J�~�(�u-���G�"y�-���sF&0���{(/n*��n��!����̮��+��5�&�����n�z+U4E��4�!h [��̬nF��.�<7�6���Z�C�V�mb��t�%� �Q�����h*!��	�����g�鲌~���Pzd��|+�c�v�TF� n@�����!gd�x-j�us���$h�VǭT���K<�+;�e"f�I!k �P��~0$���������x�+�!�M�b�N��&$CVe��;��zl�+ʂ�Ә�3�\[��X8�VU��X�	�I��a��	yp�6�-奚K� ��ԔNWԳ��C!q�"�����K����~�Sù`��[����+SۑA\6Q���q��_u
c�
(7p�\��@k�J����X�]��j�Άi�Q�	�7�c-[�H+�J�
H�2�[ԗV�g�4S���h�2l]�;P���8����:��FNo��#s���*��ao�ڎ<e�N����D�9�}]7�N�N�X�mlp{'�cȽ�2�����D�9DA�챕��n�q�N&�6�,��8�����yQ�E�����Љ�{?�6�6:� ��͎�YomC�L��ֳ��g�#�q�\6�R ��DQ	QC��������� ��dh4�jT��i���+1[�S?c�q��F�x����l�.� j/�}��V�����/D�Ʉ�������f_K�fjǛ�O7H�-dpq0��>�ЅhZ5�?�w�N�{O��l�J�m�M��渉���Y�xlO�1 ��zc��o�D��?.���D����'i���=܏09��unʺF)�l$�'�e��Iiߝ�)6�u��RCIw������u9���/<��\�8�|�CpEPU�`�J1>0S���%H�0v$�}��"~���9H�'-�BP����BQ�ﹷ�[
��+L�F�����b��U�{�	PU������Q/�ٍ���XO:��;L3�/�ׁ{���`�Z.'�)n!d�Ɯ��eF0�O�n�V��I�X'���ȿ�z�2T"��~�V����Aɺ�٪�w����]��@W.,e�k0�`{QQ�b��r�[F����τ��,�>W��?��#���
Λ�hZ�%�<{q�H^y9!��>{B����(�cT���&Y�`,��s�*��k+ �C,���3��GÓ��k����?��g�x�x,��,�d>V	��]����C��[��m�i��3��N�:�TR��u�r�R��4y"X��Z铉�>�����5[,����L�Z�E�l��֖��)�t���M�f/'��<���AS��]mK����Ȫ�ieÞ16���ޘmC����fǠ���L����Ċ�ۘ������@��(�z��P�n԰�h;��-?�Bv	�>Ʀ��v�*HK��m����J�?��3��l��_aށ,׾k��84xޕ%�� HϞF裸��9�&E�I�^����n�de%�Ƭ��U�W�bF�*��pcH��K��Ģ��d���M��0c�����d���Vgs�z� 4��>JjB#� f$U��*�S�i�M�����=��N�d�݉�7>�b�y��==%���F�cP�a���Hh�`&;�b��?�Ѕ*��X�O�E=�Dg���د7�d�(\;�s��s���9d��>Z�
��*�S ]��k�T�.�g�E-�+��Ba��e�
�#��cYo&0��#����͓�/�m
OW�i7��3�ĺ����]�x8/lHI	L�!�7�ڟs��2���M���w19��`S�ԣbf|q%���ޭZ��10�È���c�7)]Q�e�wm
iOhO�������J� \�.��}֔�WS��'�λ}`s�������!�Ύ
#����^NTl�u߇q�1�.�3�!��H���w;KGĝ�'
iH��
���Y�Ik\֝���J�s��y
İn����~R��������M�p�oƍ��AM�P<E�j=i��M!nX��;c����޾�~]U����y!K��sSzܿ�v�U�L��v��Z啧�V��*f�긹�Q�^B�r��|I�k�b	��$�5���2�٬��g�e�{�ʼԄ�y��mPNM�\�L?����D���
�q�Ғ��گ�\ ��g�����_��(e{�_w��rWU��TI�&j���;�(z�
��ai��m�qN�(��������(�љ�Xa�����
³�?pP�u4�x��e�����)��Y,F����w�sG�[.��,�1(k�.�"��1�1c���T���x�㈹��@6�c01���U�Պp��v�zwk��}��V�N$|>K8��,5�[XZ4~Z3���h���QN>(NG��,cù��7��'�C�,�tX�&~#y;so@�Q�G�Ca���8 � *HXz)ʳ�)�}��I��}�:�Ijg�^{ �!w��L�;���^�\r����/`	J&7y�)Qi`��� +����.���Z�)xKڱ[����ÉP�	�e��s��z����M�7�`�0V�l��H�M�s���<��yL!"gu��i�J�6Bfs8��	h�Ig����(�1����i�)�M�B�|�VǑ��`hF�"y��y&�(��>��H�]bb��Qk�9"]}��ٟ~��8�����k�.�Ŋ��������q������x��5�� ��pZ�t�	 dU.���@z(;ΰ6k/�d���_}b��ZHbD3<
g�opNV[(�ْ페��'�Y��w��%���1�\�c��+i�WaRАD��<�L�#8B/�* �ݑO�H/��/ിn&6�s-94�T]�e���,��(����R����M�����_IOD��S�hYJ�ˍm�N�r�q|����*�w�]o(O�o���{á��Y���X�fA_]�Q��(����}�p�ԈG÷�z��H�z����Bޜ�v�e�$4�bC�U��Ͼ]��E��PA��A5/����V��Oy�ש�̝�j=�����'�j"Z43���#%�Y�_��J��ʺ"���^�K�F�`�d�z���ފ4������ �WR!$b~��U���A�b+K�u�-��kԠ�t�^�?�01��d�F���4��*+Aʜ���{z���;�FKF8���*��{	:1�wH�f�₻�J(�=$�ps�-�~t�t��;�u�ӎF�I�ƥ��M�L�@�+���K-�y�.I�d�|7����Wd�F�0˹�Dx�U��L��2��ZY<!�F��~��7	I�t���H�U����$J-$�M���r��枭?�y��sc=$r�تL�
�������jM��{V�m��G�:��rl@�
�`�%P��.Vl�Q ,��4��~�*���ņG ��X���f&r�(ҪMJib���o�W�^>�k�-�p3YOH	q0u���(�x[��W�Jd\>C���ʼd���|���i2�U��^��rc�������I |����ֿ��' g����ۿ(�<epp�>s�:�����uaK�s������Iۏp���Մ8o���\�We���`�eǭ���ړ���x�X�zΠ����6��e)���!��9EI�Y�)�>�6im��"_K��A��c���'+�"�&N��L�.L��}V���B��Lw`0g�����{���M7���t�����Y�LXe�k  赎�ʗ����J<v��Sa���n������e9kK����z{�ꓽ����t�?�����;-��������AG����Z�>!�]�K��um��`�/�?+G)�G�U���[�Y�F��EYK��g�E=��񐡰~���QR$>�� ,���°Y�����D30Q� ����A?�!'P�Z�ٵ�a�o��t	y�8��W�^����2s�J"%�t���S���h���L,'e���ݸ��=jgl��uLfM+@fh���d<��A-Eb��p�̄A��}�4�b�s���[�(�� ��d��\8lz&�ԵxFܪQJ-	�(�T� ��RZ��
T��oI%/ mȮ�'�x�9Id|��¦)���m��#_����@��ăe��Ա�5� N�&���),�A�<F&L`��|1��fm�T���f�2�R
���!����p�L���K"4X�珸��t���߮EKWF}��ҟE&��T`��B �E<���X��22�=��"?9�-3�T�W��o���&8ɒ*���|�S�����"-�!҉TY'7W�A����?�0����8 ��I��V�c>\{\f���q��^d������I;b����P<]Sj���b��\��;�TO��6~~��d�ts$g2���:&(��h����7�u�{��J��	Y^�>0������[^Ԅ�I��+�3[�+��J�'4����J���.
�\�����{6�]�L��(<��;D8�Ab:��ƿ�d�V�: ��pW��o�HG����w�+�,G�f*��m�DBl?�_��X��w�[_���=��|�*��A�
�|��
q�n�Í5����?Z-MzHѐ�@Bc��)�+3����+R���oV0��
'�Ĥ���D��`�h̟�0(A�!o���P��=�[X�!�;�np���;k�/�~�e����@��_Vi��7n�x���97�f�s���p��	��1�����,�+HWg�·y
&�$'���Zބ�|����00���M��]Z��C�;���b�3E ��f�w/췷�6GHg��ԘChq�@]�!�·M�q��r���G���ܥfb�Y� J٤h��3&^�̍�	�K#�C�ڈ��`��J�̞C!n���:����\�󜮕�Vte�]��]�X�����g�h�#C�td��@����ϟTXȭ���`4��"��e�>V�G��@ 2]I��ַ�f��*G`�wl�%t��nT}��;���c�Ծ��$�k�}��.@�S�q��=��s�Y�ft��'�>r���-{������ͯ�+��O5������>�H�q���|�TI�Hm���cvz��"R��鉶���Z��y+_9����!� �_�/3ԎJ�� K�H��޴bN��k�R�#�e�!�9)�g5�	&&�����+�V���vt�3���ܙR[8abp��6k�A� �Q�y,�g�	T�1F�`�� �Q�GEQ���U��l�v�
��Y�t;l�	1\�/�"��8&\Ւ��$�������T�Z22���[w"±��K���t��8s	��w5R=�qRE�#G�6�]����a��,T������0�p!c�P���d<U���V���E�eB�jrB$�w~�G��>�vn���9i4Ne���'����Kd!t/ĵ�>��_?R`~;�e��3!�Pe2�hb�b���1;����;��!k2�+(Q.��j������?��@\sґ���S�zg��U8+�JW۽wa*J�k��z�7Ƅ����,�� <�l����;�sf�:p	iej�{�<��I�\Rͯ�C��qûF`�DJp��#��&�>3��P�s��+f��:��_]Qr��g{]������!���h��t����$�ٛ$��f��lpeV��E�*��|+;�uoz����O-�����h�J�ܓ���W�Z"Z9��K���8n<x�OX�c�3�ϒϵ<�/��U'��ؤp7�p�Ai����*S�L#z�J �1ZU���o˃R��EJD�1�K��y�he�&�ȭ��~m��Q�d�W��9ÿ[�Ǎ%v��ڈ/����Z�:--i�/1���mM���
L���v���FY�t��A1����1�X�QX�]�\�<��X�,���7J�'�����y��P�Q����ZB��p	���A�:;��ь8���P5#om|�ʇl�p��R���ϲ�}�'"BD뜭ḽ�x�A&S�n��v�0M�b�Q�0kz�k*�zW��P���*���������L;y�U-��Y����?�����G��Nh)@�]:R쒎��;�V�E֗�X���U�-�^�hɞ��eM�ʞ	(D��x��^�����{���� �K)���<3�WPa%o��ۍ��>MP@�1Z�;Sv<����w[��}���}z�MQ����l�
��D���N�PL�X��R��',w�b*����.�8��1,�T}t{ۺ�>B~��C�>K닓腯G�`2]�U�a��P˃J������<m)4�Bu\�M>e����E�-*Ӓ����^�Wo��0��D6 �����()ؑR~)k'��d�	y���
ŷ�G�b��J7���?S/�v�'�4� ���q?�<����?v=0��F��xG�����S��ĵ;(����K�rw�N��!��Z��aed�����=���Um�Y{׀dtJ�Q�{�\�J��s<��~mX:�G,�ݓǂ�m7 *swN�ge~¾�[�Ahlc��kŀ�xA���[� 3a�Eh���y���m�n�G!�!%�A����{k6"��L`���l�#��:xل����1�\m%�����+�K3t�.��f�]Z�TG�o���=��@T�˧T��m����U�S7�#�<��@�WhT3��po�	r
�P;"�P1�lQK(`ߧ &��f!����.�	��p��>.�9���ڕ�����9�~�����zu�a���O�����jc�7����;%�ď.e�6�^�)5̩��ne$����=�(E􄰐�dq�T�j�0�k&8�+�� Ӈ~we�����Y��b�p$�p9D��ƫ{���;��0#����1(�����O>�r7�j�+qUccs����_��Ln�u�ɣ�I�\X�D1��x[�V��w��y��:�p)toN��dw���9�fb��T=����J��iۺF���(h3T9�Og�L8�бz���q��}�\[?����E��K�ze?1r���K�ʾ�ܕl1��l�5��T�`�z��Q[��%�n����+X@�C�L.$��`㧪�]9����][Ѿ}h�Hs�D6!���
�?"�ɯ�{N;-����/�*�B����f�+��"U�ƃ���l/0�L�Ǥf+9�)�࣯�?��7����+ ��Th��ztյKD����7<���K����o	g}��"{���O{,���#D�ͽ�rQ�m��*!�zQ�yb���ku¹\q�X$��[�ik%������f/�r�Rl.�²�"�8|KS�.���'��_Bm���5e���~N��X�q�;�x�4�)R�VX�����ꥈ�$�mɼr�[Q�cw�fwoMؑ�2�L�G����s�q�&@\��=+�G��8lj��e�D.��w;J[���z�ȱ4���05�+ߺ��l-��CȀ�	u<`�9Y�Z�/��jXm�Z�u�T�����|��V�u��O^��:<��Ob��E(�07op�:�
�}�W}��4���ef�ES,�R>�s_K�S@	E�����E�p찻��D�Q���.��K��L�EB��oM~�N��d-�2���k����7n�qWՁ��y��QM�&O���F�d������aN4�g>L�x�O(�n0e-�%g�]�}���˦�i�r�����1��e5\:�\yδ�	����h���HG ��A�	A�D�㖅��LG�s��P`��{��辒�Ӿӊ2j!��
.�0�YA�3�j�0m��\p����Hu\i9���b����ݑ���Iu�H�,�b��טG@p�oVzͽigj㘤�;(��l�C3�K�f_�l.E��4T�� o��o�8R��"�>�� K��)�@6B��V�B'/��$."y�&+��lX���5�&'_�5�	Q��u{ƒ-qMt�?N^*zQ�����B�>*�V&����謬t�q�O_W�N�k�ث����Rl��8�ƥ�?�irK�\��)��Q���������5&A,I1���*\�� Yģ=��dR�B�LV��+�D�>|���Ş�6��r�HA��YF���l��Z���&}@�Y�wEt�Ԉ�+#��-������2)�[�_��9������C���R�J���2ݠ e�Dl�6� Y���J�Z ����I��Y��q�B�/+rƲjI�S-3w�~�R{��+A?�C�)j�ř�(��\c2tX�@65�(U���F ��2�U�;��U%�o��)����5����(�Y�FP1;����_���@I�2Ȅ��x�kV��$c#}�H��x��7{3j��38���;�(��V��v�]�GGצ3�8�����X�lًɝ*+$��4.�f�R-��p�5���E��j����YG6#��<`�C3v̷�NtU�#�th�.��cO����}��\�����LB��������d�F#;���Y�S��9bE�c�QB��Q�C"ŕS�o8X{
-�K0֠w\5�5�֭�\`8�+��s�aqH�o�D���Ճ�1V�Y��$	�V;6hܘT?�DH�呕�6]�k+���W�H(]�Z��]<�
 �7��*�(b{�6� �ى	"��2�>2�k�*�.o�b���o�^"�