��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��e�ik3�������w$����g|��J^]�e������	P-}2XyI�F���rZl�;���ј+؆u�8� �΋��G����%	��m�.G���b�$"§k������k�>��}3"�B/^�A#�x�k�Z���AD��O��#n1�y]��I@�� Ŧ�1-@?S<D�#.e�� ��ׁ��@��R?���� k�^���a�{�r/W_~�����2���`�I��x�s�?��|��OZ���?��ᩑ֥0�-�	�Q���a�P��d������zVJ�>� �E�t�>ϼM2�d��S���R��k�p&�VX^v����%c@q'�\�
��ʁ�r( 8Wu/Q}�.����ʅ����G�IHܶW���b�W��Z!~쮔[g
T�1������p{��I�1�䖀Qe�1���*R�-���SB�w�|d�7�{��g��0��� �[/��L�+6�Φ7?���i���z@��{��8�w�#����=��g��*o��O� �p22���^ދ%'(|g��uޖ�*��Z��B��D���.ถ\ad�6=N9P)n�� <��5kwj�}D�ePpDa���6WI؋�G��7�]���R���"��� _,�&@dQE��4�;63(v��Y�`�V2��,)q�C���#b~��HR�d ��瀋��!�+�v�m��y�tMR@U5�#�gp��2{�2�D�K@
�˜� ��|ٯ*���#�}j�UU�y�ʠ:�R����/��O�j�L LՐDQ�h%���׏�;�����Na�8�lf���AD�ZՂ?�E��)1���ߊ��K�/U1|&hH��ϻ����pO���V�|n�o:~5���^���s�+���T#X{%�N��,���S�˧��Tnb;#�����B�e�������u*7�Ķ>0����eκ*q��N�_�������y%`�����-����N|��OجÙ'��]7���M�w9�;I�U�F�%p�h(�Vؤ�2H�#��H�R����K��	�T4��m��Y��~4�1O�>T��qL�Ϗl��BAd�Ҍ	��A�,�=�������3C0�S��N8)F�N��H={�Ol��T�����Q�޻'_}�����co�AV�Խ
�y���ؑ���?�w�~��7�Z���%A�`/ˉ2a΃�	�Ks#����yDc�>Ѿ�VՓ9�t.�X.�|C�����Q��Y�#��lVq�`W���GOM[k˿[̨�����pz�C������Waw1���7�;VRh���E�n�A����<+.���zp"^��L~	�X,=���ıj�m�ߐ����
�����b3gI�&:IǊ3�K���x�h:�+��d��_ ��X3aH�K��a�.8�Dn+����6�5�ďy�|���^�$���ͅ5��Q~
7��a�7n>���Q�JR���q�s�����	���Ė����"��,�P}�ICڲ�X;xaδ�KU�`"4d��F�	�(97�ݣ.2u�z,`��)3��\��o�q���	����w��Ġ�q�{{{Q�Ϡ�p���<��0�$_�sO��*��]6���)��c�r3搾���R��E׳��'p����g�%�qX8h�)�{��h��H�ۥ��U���R�@�k����:�B3L���u� �[�";����]�eK�3$ޙg:X �;��%G���^t�F���њײ��(oM�z�gN��`���FR�JG^�P��	��5`^T�YDk'"ɓ���q����Te2�'Vl�y���L��%]A�Zz�.>B��꿟V�m�
�Am��E��"j��1!0�-/���T?%M���%�� llX�G d���3��I7[�X���Q�;L|�@���sq�8������oU�Un�GS��j����)�SKE�����+��C�Øh���������&�چ;��f��Z�HӴX���� �E~�eU'�M�`����xI7Da%EwI�k޷�GD�p��2�U�����r�ge�I�Z���(��A�T&� ��H����TM�������ǲ��(g*mQ��4PIG�#v��U[ɤ c����e�U�	r��\=�>���(�q���0 �h��d)v��W�t"s��#m .�ep�a��&���y1�'yYiၿ-#z�D�Ϲr>ޡA!�yeܛ�x?��I�xئV�D]>=�(['�	0>~��C���L���>�O�;����ТZk� ��@�
q��;��O� Q�ۯį����\��د"�/m���#p{b�K�.85Q#U�G�śQ�2���GY��*���:҆w���m��,-��ӏ�9`�����ؓ�A�;�w	{B!�����ڱ~���P���n��WN���&
���� �QF�"��#V_85',�Ѻ�I��b%��?����@ %��_�;�4n�q~EZz��s晴=R�qQ�΀Pd��Cް9s�IU '�!oD*,���	�~7W$D��=����;,��-�E��gG'��j������bܶc�8�'=_l��A��L&T���m6�\��־�Pݓ|��^Z�䭺�=G��v�i��ۨ~�Ĥ����]�����v�Z��)��Y�*��2���.!,�E�kc��P���Y|5����}?��gM��D�ЊGl7��� �vZ���<JN=+5����/��&����D�O7ѐK:pnJQ��, bl~R�xP.��z����j�l,�(��y��� iL�ik'�� �7��UT^\�g�m�mt�v\�+}gX�8��lK�����<�}6�d%�{�GY[�M�Z��dȠ����/,�"ac��֔b���n�j��Zu������k\0�s
c(�bCJ����v�)RQjV_E�-�YM����R�����V�E9��3g���^mF^�JSC��i���`�����`�49�� n�p�H���_������~H��ψl�������wz;g�դ�`�D�WYRK����]��I��c�J퍩?�Ш�4�F��R�(�o��r[�5۠�kU��fY�u�A�N��I9u�N��Qo5w✑��� �7��~�A�!5L���%�@N�[�O���q�Z� PXo;D�+5V��2r��U���7@X�P�8�,�5~�_}sa�dگ��f�p���Zd�}�Wu��X��<M^l��g�!U�����O{��_Q�YH��4�"B�+ù�dh{�	Rm�d�F��:K#z\
U���c���F�x/:J�+��405e鬴h��O-��ΰ9����J�wd��R&����<�P���$�^��\�%��yp����3��� ��gA t�P�ړ&:a��K���Ƨ/3���]��k��\r�����*�!gr=�k�1P�������z-+j¦�����A��Xܱ:�w[����;u�[$��cb:Ze�V��CG�J�qS]B�F�凞��r�64X���Pg��Pvod[�Ni��v�㼻�Z�T9Lm��2a�v���
A�����q.,?@`hW�{�CE�#g�$=r'>*,��4�eHS.bY�X�4�a��mMӯ~"����?ڳ���XK/1�)R<�b��
nh�GM���ĵ�.��3T�7=�N3_ H��/R�O�2uJn�3I�!&�n�`�R�u/T�Q��Y�:?�,�&���:���v�e�����M��G����p
�/�W^����Tv�퍼0q��_��W�X�uF��E���� ��u��#��V�/4�FB���0Q��Q�a���2zh���	�";D�����	a;�ye�5��V��2��3��Qp��X���7$e�p���OY�B���q��Oυ���2��V�_ʻF�D<]1cǫ�C������lom�*��$S�޽�<@D6%�R9�e��ʶ�
`���XG�΄�j�U�Y��&��Ҧ|O���-#8ժ�tpT����u��8rH :hg�����f�ۭ���r�[e��߮^�C٨ ���̌kl%[�=�����hҖe��8\Ƿ��J%$������B�}����zG�����)o'��s��m��L�e%�� �ɋp�h��,�����m��[�������������Qr�(�D�{�y������V��d�3��&bq��yk�y�Q��z��UN�4l�����AR���rz����6�1�F����^psV����U!B�3L�E���5�Y�����:����4A���9� 9	s���߭���N:����Ar��j�]�:�Oh�jq����*' [w�ȒH����ւ��|���K�z<پ��zO]'S_>���C��%<t��6��OƵN�v��>h8��S-c%���~J} �$r���&4�>�]H *����&�%��M�ş�~�cX�TX�k��uP;�T����\�����h�E^2�Mn����(��j�4Yp�ݗi.�ǐs<9��}���"��=/p�a�7��!��"x���J��#<�_;O�^�j�d�Z3�<�p�"�<� �=!J��Z��B�V7�vsz	�w�/�*���b�ւ�K�`qՃ������+zZ��*�/�&��U#�E��\,�{�
��M4]d��+<��c�PO��T������ʆ�%�j�V��3@h׈ō�&�Z��#&-e�/cC�6�Ys�d\4N	�__�:�p�99��g7GD����!�@>9P���j���L��(vR�8��Oo��m+���g����z1����BM$�f뛎�� �ވ(1��b�<4�pRo���G�X�V(�(1��O���7� �),W�H�Y�h�_��V�$�@6�/:fе��Vs?S^�oL������.�#SKKrM�7"t�uq��־�]@��[˯��I�BoGvϛ��u����h�ܐ��|�Wb5�N��5�-K[jKϻS�����������oi����u��g��
p�?���vr�0�^���ܽշ�;��� ࢝v�٢�rH���QRb�L�ꞓNS�3�+ձex����_va����aq�w��և�^�G��F��d��{����]]�)�Aڦb'͊��r��%��};��� t����Ep��0�����_��1��Wm� Iل�]�g�f����^C�*�Ķ{as��{�X��hv{qXE�CH@0��A�؈��8sc
k�,v��ꢇO`�P�	��cU�p��u:�ώ�/�n�
E����G��c��&�(��C6��8�ё.��~ZĊX�g��ɀ���@�ġ�YT�(�PP_�Z����kM���� *�dS|�2���2J�g��<p�E{�T#_��](ѽ:xY�r�Đ%>����'�[�2���L�aB�,� Y5��OQ`u���a�Ǳ��Y���d�E
�O��v���L����x��h���<U_��{u����u����m1�ɝ�$�l3\R���ŉ�*��� Q�K`����O�^��CK�����QM��.ͣ.�7ownU�K?(Y�=�;S�ty��j��CEKh�/^RL3kc ��#-���z �^�f]���Š9��T�A7vgd�tV��ܜ�rkQf�JC��&GR�<r����"��|���,~\�����%��Ҵ�Qv��|h��g�P~9�nx��Z��� }�����{����Yڞy��:h��b��
��4: ���rWi����G�k�������>�r����Y?�>ZL�Ҟz��PJS�B��h��.Sb5��t�\k�URv�c�W���,���m�S�~g���0?����'#��הOk_�Qϭ�k �R������b=�b3���#
��g�>QQ ���"� p���<HE%�6�8��G�5�9[�o�%�/�YJJ����m"��SdOf�;�i���v��۸���"����!�t3��3�3�hk����M�R�8�����I$��b��F�*5��b���At����QJ��}Nf�U^�W�}����\t��;'PVg����+N�}W�������a�w�g��3�v"�̤�î/�yf���ER)�˥��6 ,zv5f������Du��oIj�4g�;š����@c#Z�����a��r!�Lɒ���Hn?.]�d�<G���Ù���J9^�p1zN�Xvț��-xO�q�����`ƭ�M趟UQ���K�(@f� �J���4����ʹ�/W���V]�`�o�`U�ҫ�hM������
}(�E�=H����灹t�c��;�_���A52|��{!�!���r�tl��Am��F�&_ܺ>���%��͏��G˒��G�PlH��q��u�2|�O}j����d��J'j����fR:6<��t�'���Ewo������4��>\|�g�w�?v(6�1Mv�bI�U����B��@HbZ���d+�k�kS����5��Ӳi�?8�&�Z�8�9�[U��"v^�	�%U�h��Zt�����z� ���3�8���Q��W����o\�U &�!�X*�,Ǉ��������Y�oz�W��R|몜�c?@��b	r�������k����9�"VB��yn?�+^pĹ-jl����9x���5�c��r(�)��BZђz8�64 �W�|ce�RUeFH�z-��"&�S+��57��9�7��-����`�6�f*�Ub�$1��3q�Y�Y9{���<�Q�l+)��/�L��2piMZ%~�.  n���j1w(��;tY��/f�ZF'!J��!�0�"��^SA���NQ��T2DWy+Rc/
�B�epj�G����G�?H0�����|�2���Y�k��l�+�w�����"*[�m�d�'�� /�2��z�JjIC�L1<�$œ�.sAI���m_�Y�Z�n��
���H0Hv~;�բE� ec^x
¬t�K>UaD�j�8�v�>u�XQ�r��ͪb��Ŏ�����ǋ���+�x©��5��+�ɔcLVIl�f>Fy2�z��D鞴�+�52oA��|]�/d�3T�9N_�H��Rz{�@Up*��r��5��ɢ��=�	Jh)&����I��uu�r�߾b�>�p�Yj�?T�Ei|���'�^�8o�B��4���Lki5�N�����7��n[� Uq=6}�����Ė�w{=��7�ayhf)����&6�ny��%-oe/��}*���8/��H�� z�)�oOc�rT��l?�&���O�7�N���!(��f4�y�L���l:_�k�'�<��+���s.٥j�^-�W?=��8�E���U٘�V�˶�q��ʃxm���I,�l�����?ۑ����ǔ�K6	qg�ugU6^C�Ҽn�q+ֱ�~E�۴�_=������IAT�b�&�h��D�!�6�6��A�~r�"N�_��%Q��s=�gЧ��L���Tl�a�����HU�S!�&�ظ��;�����q"���ˠ�t�5�#�ϙ. ����Z6�55kt)�`���SW�lD��h˩��֚=���?��K�	��bny{�>;� ��U���8�`:���r��N�c���?����ĸ�{x�����~D0�w�O���/�\ϐ�|�v�P����l]�I��Q�SE<���D�I����Y*>�]1R�^����a	ß���d=��`rS,�U��Ds#I�E��Q�g�9Z�I)��-,�΁�)��i��,򝌙D��Ba�8�)y�6]���;���h��\i��!�e:�zUR&N.�`%p�7��3��/���ރ�AO*aMIoT�WT="��r�w������f��������J4�hs�I�,ˢ�gQ2�v=��c>��Q=��_YH�Z�L�%�Y�5�nQ�`��k෦)¦�=c��#N)��C��=�),��;����f�<gȢ�D��D����TŊ��簸9a	��&]�yt2�w�خ+K>��B��Ï��8�׾.��-qi�&Y�Z)a��b+�sI���sƢ̦6�ey|�K
Ac+�>���C1�\��u$�s��g��]��r)�'�~/�4s���n�����]T|d�VOΩ��F�����I�lD�-$�Q����9V�����,�=���e��SC��J�I�2V���)SVlރ�G	kw��'D�ι�ߨ���J�J�d��f��w�M��P�O�#//V�q�/S��?����1	���k���$��/Q9�t?w����X'��ie�Xt"��'�����Ò�������.^`��EP;U����=M5���Lpʆ]��gn(��N�f���/�3l���D�*�	�ԗ��Q\U��~`�kᐯJ�)��Vֿ.=t��hP^���اE�*'%�tw7D{�؆�L"İ�F����R�6aZ"�3�`}�*zD��a�@^�0s��9�7����@���0W7 ��>7=В�0��sgطf�7��Cv���>��B�*�����,���J�P�(�B}��v�^��m�JI�ˀ��(�k�g��f@�Z%L54�n��F^��z��;�^��͙_4����"xf��H"�mk�D�2��V��i,����c#�h(57������ަ�y�9�I{b���h���>XT�ݻs��en=��ۡD�xp��+�5��V5�����T8�z"�+�f|kO=��Ȱ3��ph��$���㍈�v��pk�p�#ֈ�� 1�k�~v�f&(PyC1����~��_ң��'��'Ot`2�Ih C9)�[��TF���ތ�������hϭ��ضk��3y�{q����m\���f̌�V~�C>5��D�S쟹 G���ҙje�E �����tpn$uy�`Y�3'ec�0��m"�����F�4��!�+�m�e<*��Z#��M���Rv|����Ǎ"��iy�RY ��u�p�A1ں�0�UDe���Z4	%�&>	�b����V"�'�y=i/�@=����B�9�Nf��� ����w�d�^Y�c���6�h���I��X�F�a٢K����jʉ�ߨa��(��M^�m7u�+���j_V'=�����)-��G�J|#x�FW.����V��j^%��p�hB�F�Ԁ�Oך� l��kD́�/~3k�� D�rg�H�"&�z�r�nj���&��H>]<����'M/bv��1p�)֒v�(5�_n���w�� ��4$A��4�()�SZȚ�Smڹ�h�t�vo����Rz�]c3m�'���_?���Ť��?(JX��o%�o�u��._�$�,+M��!l����`R"�.і�܅:wIP��˗�B!)F�v�.˝V���/�O*���×s:����k��Wxk��%)�0 ��	I��?5����Px"-,hݿ���VM�=�d�w.}���h���4�*35$�G�T/�	��:7Q5-[���X:�'�{��e�� �m���lū��Mj3�s��Qڄ�l��Y�}f��`o �������4�}���66r�!� ����dM%a�E���g�%��4J�~��h��������_�u�����d��M������6|F8����BAvPJľ4~G����B��&p��N������/�-����zL;��0�{����r;_;�;��f�̀�5qߝ�	u7A�~V����댶"/)�].���0L���zQ�֣��9��;���XB��i0$�1!��K)��h��FDtU{�I"��N�9&x�R��#좶	�o�ь�kP%�dR> (��$g�8�;q �6Z�����L�7�ٝb��h&e��[dF�F2�W�n�]���S��S*({��\�Ǹ�bB^�֪�7�4m
�<��:e�i�4(���EJ�͝w+ݑ���^�|�W�$�<|�-�h)ܣ0�9��FU�����EҎf�#�&TpQƶ���U��|��W���ɵe���e����,��&Qj�F�7���R �`fr@W�q2�ӏ�̭�(D�@u��i�f�a��d%����*�I�R��Z4�ջX�ѱ�����i��l�~E`O�.���R~�=!J�P	�ӧ��g�n�E�Sd���c�9����J}0�d�F��[xȮ�h����8.CY�8�/N<f��s\��ݴҤ��m����JE��(c���rE~�~n�|�L�5�x'	Z7FQ�j����v����]��>��,�
�ez8T�i���MƂ���\���o�I�{��=���!�mV��\�`�]]�+'鍚��y)�s���)N�!y�U��.h�p_���L����:�4V�T$
o�s+ٿ玞M����q
0d
j��+^d��AM�Y>��yʞ0��c�|%������>�I�}V���A��]^�/3Iݴ�:M���>&�o�T�J탌ٝ�)��;�	a-5-I�ڠL��Hf/Z(G+*��hV'p����,�ɛ�,��	�E�E-��_Z�IA�N�0jN�>��d��%RIXb��R��S �������\�˜�;'��l
�	Kh�7��Gf��^�΄_��\�O�ّ�h�#і;d��a�ׯ��F\}��ۊ�5D����n�ozo���Ƅ~r�c���/�B׬�^�Uz������s���!
�&�IY2��0j��K�#�^�?��?nQ/�-����oh8x�Q-{����p��N�e�
�'�	&���z�K��!A�3j�dq�T�f�!�-�<O@<?�t��s\���+��=V7�o��9@�л�� wV����*��py+4*pIeH���͎�v�,{��f^U䠡���nq�Yx`�y> >�O?y'Is�7A0)	�B	��MJ���|	��斨��PW�*��/%4?���]ԫ�p�� ��qR���Ԍ�g��י�[��ʔz8}gl���z��?m��
;~�r��
I5�E.����\f�)9���Qd؛�K��%� ��T��@,z��M}$00�ު!;m���X�y���M���O�ph������(�ԪKc�������и�A��ņ����*�B��K�_���AT�=�7+1�8|)N�)�شm;a��&���T���-[NN��/�r�7�C�����5��P��%:�F�]�"|��o�͏O������*rؘP�P=	zl2�C�\^޷���3���0g� cV����႓��Y���7�'EZ���8\��*��1�cEv�	�Wq�y��H��u��}&�?��8۾h�XσxG�.a��i�/���d}�j�IJ:���1������L�k�?$)���p�X|cVt�f���F�?qRLB�p��"�5�uL��
Y��!���<��WS�O��56"�c��qg��h�K��(�����v�%������Y8�n�U����7�O-��#���/@�pe����x@���ìV�+�/��ѳLf����qt���W76e�k�K�K��TCA�-�/R�Q��~'�w�T�.�~ց%~S���;��]�Ԛ�T��7���O����=,H����^�5�,�(�uh���C�����}T/k�+�t��=!.�[̒�ȣ(����{Q\l����h̻:��Q���j�}:к%�b��L{�o���6�6����3�K�&	�E/�qw��X�PS����f�W��m�) �q������DI�$��f:*�EnY�m+��<:Ь��*(?"$�'5�Ҍ(e��g �t@��:��	�~gHo5>x�ԟW�A8�+){����v�n��I���0��8��&���z�R���)Ϣ��9����.t|���<}���؈:7jm��»�	�/#c5�	�nm�h�(���f
}:_=IH���L{����$u�X����C-�z?�̉�򂾷���s&b/��=ql�/&�����Be�M/�"�����
#��x%TZ0)%�6�M� c�2�B#�5mx[��Ԝ���B�:� %zNXD��o�2뱇�N��W�?����eɾC�W� ��	�%�����������]喔�e	�h��H ����C�gU�ø��pwru�u{�AҲ�������L�kt3�.��K���{x�֣�"C�tQ�����x-���s�F]�O�@6�ϙ�$�/���;��T��{�+6�%P�C=HS}Q����K��G��U��\���`���[4�7V��������
}hVD�.�@c�d}�m�d���C�Ñ�1����8�;�p��HV���}IbU�έ5�= \y,Z'� a9.���y��=���4C#=<ܹ��Ae�f�_���z2�0S�jax�4�O�JE����&�����1/������"Vܙ;M�[��>#A ´�]��mW�S�M�J�]9/����2���y�8���Z�3�l6���j��ւ4�#;"�l'H�Q�T"�$6�^5x~	b��X1:�N���y����g��ߨ��uh\F���U�g3��gg]�q���!ž��g��û([J�R/��!�}���vM$ �����s���,��?&0^UO��!f��i(��8L�snWV��h�B#uz6����X�`����m��015G�B�&X:�qO$�7F�8�i���`�l��%�{z�[�c?�Ά�񥼭9�'�d�4Vݟ�8��`W��e�d5a�m��M���O ���G�m$vȱG^px�2�xj��|]�Xo '��7Mݽ'�:�Wk��@����z���x�s�$/ ����qV�J��Τ�D��+��iL�T�y���/т �