��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0]��?l
�4�!�ߦ����"�p8"	~��kB�J)��NbM�L��\jO��#y��r�3wA�y�}�S�{�����X�.m�lM(��R�g������B�*�NV�X-?����$��$�3�s�`;��y�@�u�ߗA�R�|�Ԝ�+�)]f��������҅i[^�"[��t��00��6�ĔR�*[�]�V�t���9�c%kz�Q��*N�| ea�z ��@������mU���h�$}���~�k��'C ��� Z���>J����ׯ,�'��3@akCc�U�U��?��a	6S��K󊀧uh���Z��&���9�+�)�b�В���ɀ�t�]z[��z�/`� !g�!*��P�����I�<V�� /o"�����@�g柅˳���.���5����9�i��)�!Ҏ���f8�vh�3�Z��ZC�:3Ϲ@�+��&�Ư���	��������Ϋ< �����"�����!b�'G����Z�!�R�l��Ã���3�����y���H�>����/{���?R%|��n6���gJ�2!b/ΧW�}�/FM��%����� ǜBk{�.�-�ّWz�*J`����'29�05�J�NYŪԚ��N�F2���������q��y�-Y�	����D�0���7��%��,�-.�O,P�y�w	�	�JT6'�Z�Ҟ���4��\��י����Ə��g��y��E��q�"�ӊ��N���H��`����=l�r�Ed�tP\��� �c�G�����/�('�'˷5����+��3]ʸ�:xõ|D,"���V�d�@��^Nm�D�dK�+l����E�ȟ��_��O�՟	����ȢM�6��������U�²��;偐&r�+����q���_j/�/3Ew�?'�Y���7ϓ,4���W�X�`]���eop�B����nIN�_K�����+�-�J��^��8��c�.)��+eR\_�-�/��?���}��@�|�VBp�zq�4���tsT������wPφ�(�,/��3�3~����]4�_x}����M��t,�Wv,�,�t����#���ιXz�^U��#|n���q��LlW�'_�@aQ�Ѽ��Սu�7�q��"�u$��NɌ�mL�d�"���e�%4� (
k_}6�T�\KMW�(1(�&6�w�rPX���.Y�u��cY�dI2������fۻ��Y r��s2��y����X?�S���2Pt�(gp�o�/�`��:9�2�ύ�
��A0�;��������j
1���P�o6{Q���!���K1Y���j���?��"'����)�I���G��𿫢����K�q4�ަ&m�i��N��ko�����h��]��`f�0��k��Bx���ë)JV瑜--�'�q�
�h�Yjj���O�t��w��S�v���Xt=X}�JˇF�L��qɔ>�#Q8�T �;��ԅ�>��6tph~�nJk�a�ayN!����P��U
{M��.��C&�-����b2�%~J; )WA9�$���AXY����L��L�Tt�u��wh�W�p�A�������F�j�1/U�Vy�h���Y���Ĭ�����+g��Hں���<@+fP{W�8��`��+��B����Oj��D]�՟j�Ԕ/8qL�nزC������X)z��8p��0��ZԨ?�z��X�U*9��Z����iTH���UU~;Q�	i���Tb�Kė�i��S�8�Į��b|h�,�9~������.�g� ��u5F��	��V�$Y��Q ��*Dw��r}{'����!W�,)(��T��U�رm��Ӵgc�T檟�d�\���pO�o���xz�}9W�Y�mq�x]v�"��v|�ux1��=Yn[�%]�5M��{j�Z6:����"|�ۘ�}��qǴ|A�"Uʑ�Z���(�ʌT�0֖W��w�!��-m9��.�)&�"<���ʉ}�B"#l:�}+k�d,9C06��u�j^���
���b��Ǖe|� ��2�<��s�����:ł�L��-n���א�B/�秄�B���T�A@��+A�l�Yz3�U�T��v��E�-VU�Qk�+�w�8��_��ۭ\,��5Q,/@`����A
g:��2����!!��ðUI��cD}ʿ#�i�6��§UO9�H�
�{	�Hj�VXG#�}���FX\���W��$���7�܊�7�'�m{|�=�G�8gJ�f��U��Ϻ��[�H���4�	�v1.W1.����s��[_&�N�K�g�(=��Z��1_�R$�Ƭ���ĺ!��=#����8�I���D�B06^/��@��!�Ֆ��8H�ͯ�<�ex�J���e�O�P�ł�L��3u� �`x5,R��H�J��4��Z��N�
 ��F�;e;餼4B��PݞdlMt�__x�!H