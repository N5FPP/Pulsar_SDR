��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^0�"��l8���ƙX/�H�#H>��X[��M�w����ҽ��P�鶡�þ�I��mVݷM�Y��j��im��+�|B��YR9���}�$��9J�z=���r�4b���t���`M�u��Y}�*Ɯa��|���6\��1�}KE���)1��ˡ�(�OZ���\�F^��xm�?�##y�h�Mc>���Y�P�Sik���",���c<B���&hLH��������)���Q�(O9ZTP�1��
�yM��x�2�1�vw_�T)'n���݊�'KtN���1EPJ�����վ�\����K���}�<�!�ϤV"�����4�I��N.��s��R�qZR��t�kF�]�����H��vZa(��*`�� xn�(��L�G�+Y�u-��6�=i��\�_���`��|��s�"=ȢO���qi�����vK�=k{�_�"aB�1�%R+��<C;�mXՆ�!�Y��p���qj�h�85�A�������gz�ו�݅�K��8��7�a�"�%��/�]�'j�v־;�qig���)~�+��P ��pW���S��I��x�q6+b�?V��+U�8��(� �ׇﲕ�~۔�׃�W�3���[�*�ڗ��>��C��Ab�i�Nlb����5�w�T>/��B�@,Б{���gH���ލ�@���2"4]y�+��@�8�����qS���H�<���Y\�i��>h��RE�%xURb� ggF�_��p���:�|��T	���W^�.�c��� ��m q����YZ\�.�;�gBt�GVݡ*�z��£�~+�Ac�����?m3����ᑮ�$�2��=����ۓ���s�#����v�n,��u;V��q
!�����k��PL%Hꗝc�_-�6��oq(KH�E;Z��#=����V&^I�8ªGS-d�&�ˁ������I#�#��͉K�������K|�[`��ON�ߢ���@�ֻ/����B�+�t�|�մY��`���#�:�b.c�R�7��_I�8S���T�g��>��D�h�m���0���^�騆�g����6��NY��?���4+�s��"��Ե�e~��{��T6~�od���Ty���"��Lu�SaW ϰB��c��bY�8%�h~�>�Og'$���Z��B�|s�22���v��f_4�@LX9	�4�O�i�����=�y�jJV`/n(��2���jG��*83�A��;A瓦�k�Ss����>�n�U��5�7��N��� ��,]�����g�~���*����،�i��c��r�A�(T43�o��%]�TD�{@6M�dڰro0[M���#��!�MB�m�BbF�S��|�Bh%u׼����-��$T�\/�g���1�w�r3Ү�3� ��X �P�Uq���$e�0V�@)�hҷWeg�
Xc�-��<����CtK��I\�Ÿw�)]�E$s�E-����z�b��{��;E]	�����E$����f�G�^tf��ҍ���vJГ�1h��G�?�^��̓��Sa�{">���Tv�ʖ01<�����	؍U�m) P����QM/��&s=�����aS���"n.{�����i)�x�K"^`k3	��{�k�.���]MI��SMI����*��R�3Z��{��t���9�QH
J�K'�!_�vGa`��i��b��#�y�X5��z�f ��*W�*��v�22�E+����C����'�*�8 0$��%��:�1�R�b����P��߽V�(l�v	Ѥ�sm�:[�9=��>���6��I�����M�AJ~�����������O��ሶ�G����Ƽ-� ��2d�r�O%˸�G�����|l�#�E��s[��0n{�����
����mJ��n��z+@��d���j[��������T
iE�p�/&0�l�6�rհN���{xHL�<��0�>̟�xɀ&ͦ�Fȹq�=��޸��4�:q5����K�'[P�Æ�2C���-�"ad�Ic8ߕiT%E���iʩ�3��p������a_��|�0?i�_S�$�\l�=t�P���
5?b�}�G_�Ƴ��5wT.��å��j`���h�\�
�2���+:7e�s�et�4�g�5�W.tÅ�Q��g�%6�����מ�{����'�	���a�2zs��5�X�R7+�Nl^e��6(L֦��j���(%�MS���
�F�ЭR=µt��+���w��-��
N?.��?a��2{�?`���Fw�}���!b���1�K'Q8|�r�O�9��J��]�kv ���p#J���g@�A}g�x��GV`��?��BM�mҠ�>�Y�G���w�g%f<�lv�p'%|Zz������zVI��)�^	F���a�oV
n4EΚ0�=�A�ִ1f��{7#�*t6�:45	Q=���e8����B^8/;����pdL$��=g~�pq�&��@'���wE|#GC��R�L+T|�0L�0�����o��A]�p')Z�A��j�1��/�����FEn,�}�G��.��TI|=���ky�����PY�8�Y؅{"�~ͯ �z��&���x���������e�h�����2�t�(5���Eث^���8�$V?�A�m=v)�?x&Q�v�*�K�o'im�b$<��������ZA�o!UY�=K6��hyɌ�u� ��V�j�y�X���͘�A�|_�,���u�4��.�>�\���"# k^�w D��@b�@�65�|�"`��k��R�����tJ���p<��OQl�r�:��t�����"a�	�Y�����),H'�|��Rm���/|:��|w��O����ۯ�3s�n@���׮�@��y�A��� ��FФyW�i���^���ͭ���-���%q��
-1c�~��])m� �-�V����0���1�ܻ�k����t�M��K�p{����w~z_~������|�� �1V�\Wv��퓤�O5���ߺÜxM���x����p`��d� ��i�{T���L�\	��}n�g:��� �z�$Ͼ=��4�`��:<�lf�ǎ<.I�q��5�p�)sn�=��d��^s�9�]�w��Z�����[ձl��-�@���� XC�oބ����ᚎ
.��߄0��%w�j�!'�p2=�*���Q8�i��ͮx���!�����}D�:V���w��2T��o�[�5��8�O���c����3o���K�����A��ȶ���j=��1�9���D3'lH2,�m���<�k�u�}��1�eTL.��jЋy��V}��V�^��fܳ���ثYM�#rk��Q~��i�ﴋ�a|��#ن���ŀo,>d�e!.��\�.MQ��ʳ�E�s����Oe�yA�N?fU�^����}�u}>���r����GO8�O�4/�c�pN/ڈ�P0&
�r�kr����"���~s�B�:�-�j]����3ۻ|�����9v-��Z�V�3^��7cQ��H��UR��uip%���u��u��88���%o���e �m��$���� �9Js�,6r�E(�=Q�Y�#O�9�Y��/�@,R5�V�O2�j�O���t4��S-���S�B>R�qb�z�D�}���~F�������:�+3�*$[\˺������y����cH��u�jߋԊ`|n����.Ջu�G��_�8�E��؂�N���l[2��s������`�5z�f�O������r��{ڄ#+ek�=2-�;�[�3��Z����a�������G�\�3slt�5s�ڕuC�e����������+$�������*�rA���$���V�5�o�ߙ�}�tT����h�Ώ�r�L_T1���A��Z,�%V���BǞ#�]�gxؼM<y��v�9Ԁ�����6�?����z��v���.�����VJ��TԼ�D��z_�ť
�uY�H�@�[b<�,p��Ԃ����l�A��k��S��ZR���ck(%��"Ƽ��U�D��:�&�I�	"�<�m	7$�hZF$y5�E�����-����'���ֹ�����P�-��}����*�"�l�f�rl�%�����'"!� ��kVd��?���N�=*ML�����ѭЭ`,����|ϯ�����mҩ��%�7�� �Sr]V��|#EN��:ξR��fx˂����K敬�)�|��Ү<���#SK�<�z{���My,"H�O�_���
H ���-K�
�:5|�KV��l��zzMA��Y��X��F}��y7ݧW�f׍)y甌p�=�������)���)�#�U^SPYu��cn;"W����vlK	Q=/*� �N[�Lu������\DA�( ������U:(Z���fWy`���DM��4���>�s]��|�� ��^��	�C�pN����u�%�4���T�`�f�i^�Z�Q�RX/ �ɡA�O����<'��V��w��\dnp/@C�A�bؚd���iFIړ#�C�9�aA!\OCMBw+,:�->��a����W  r��!���GD���X�1�"`wHe��S;i��8�rL\���:8\ᑏ��#�#>��$�2�
&�N���4�;!7='��r����D��A����~#|�[�|T�P<���2ڧ�"ё���Q��}�F��v�q�z&�:t�æ���:M�ɗ�=���v�3R@�j�x(�H���<�����/���|w`���)�6siˏ�+�f
�������C�[�5ƶ2�N���a��o࿰�
�QH�
���hoN3tv��e)�\��Pދ8�@����8�@X�xiwU���~�[�i��?K�ݞ=h�(�0S���q���Eh��<�<� �<������@��􎍜Y�9��Պ����Ru"-�NV҄�����u��d���^�k�/����4�0��N~��'�wg�:�+\��<�$E���%cB��?��?*��}<��Pd7��8^&c�+[p�;5���06A*>滨-��M�%c����&�����=�v�7�����!n4�����!kY�����+�:_�����.3U�|*,}��|��y tl��w�gH��t+H�E��7�Q\��p�S�;xI���$�Z�i����>DB��q���d��[8'�Bt.o̦��v�I�d!
���̬m^�0�by�J2�󞭃��_�YZ�i�q.��B:��#6�`��y�FԄ4�B��9Er��������F�5�&�B!jx@Q�nr��<<0_����M�G �Ys�d�b1>C�O�q3��I�3&)�sg�Q���1���!�t
�!
��#� l~�����)-l�D�m�[�S� i�8}��O{8��B#�X��	,��/�J��>W��U��R�֥X��#��HD���-yn�u�lD�Rd ���A+h��iA	��ӦF9�M
k���+��qY[�6��	T���o�����@���E���j�	��j�@�������1������ϟ�_����/.q���s-�bІC�4���"�T��ڄҬ�c�3Wm��P����|w��S�#���U6�C�uA�&��t�ar۰�oY���K0��P��E?�V^b��E�4����P�(������c�_�O�3��xp=Yv�XN]���a\͚J6�E�	�"H���<}LD?p�c�ᛄ���7o�F�v�Y=�{���,��t_�n��7��M �ڤ̣��+���e��,�"��ug�Jwj��FRnJ�Q�Շ�e�(��2W��/^����_�l~�,++Ղ���ϐ<��[(��y�a�i�'�.�]�H����y��UNdw�l��'x����D3b�s���ˎ����Y�a��<��v@��ȣ�`Aׯ3?��P4mԀ����R�������1̤�;��dt�EZ琩���p�QWf�����f�~y�ӗ�O�Jĥ܅R���R��h�n/�+�`�xX�M0	��nfZ��c�w	���6&u�����]�F� ;��������5;�&(]���7d��Y���+e@�!�#�ԆRԃ��+�	�r�9�"6�#�2I_ϧ�	�lE'(�_��!I]�.��ci���q����a��=��b�.Ņ6���>K�O*<l�
[=|I���G��E�8(��Lw�N�z��C�3.�w�$����~!�H�)��y���X���j>�3�RvF-ySV�!Z��2x�]V[(|y�W��/�,s�?/Lyl>/R�k��[�z�+����Ժ r�� �LTF�=�6N&[��r�u�����ýr�Ѝp8.���Sj#MZ�/u�˓��!�|}p��C���i����'�(,�ewzI�Жm8���=(W7S��#�k�DƜB	�tu���g�8g� �=XSЧ�������L Ǝ �,���$(z���������e����}�Ԁ�O�!���9�L s<�D!�4-��a�������45#(�{F���q���n�t����ߕ�m����u����>���l�;�Q�������#O<�AD�u�~r�t���dp�v�Ř9�<�%mo���P��8��!/3��7&�P>r��h���;�-K�AV�(�e��H�-]U�dJ. 1�|3�p��rue����7�k��?"Ĥ}١G����#昽E����T9yBs�y�-�3C�{�@5 �U��}��^cÕ<���J����ނ�{2�<�Ҋ�G���������*|�Uړ\��^a���z"�&��j����k�4�ml�qTvNy����1�"}u�D�Im�2�=}�#��I-H5xw�D`l %��}z޸�kʭb����q�tV�}��+�c���O���hD���Xb�!	��7]��c}�Zqtp��k��O&<U���<G�4���\�E�n۬�}F��YZ���Ca�G'�8w�EK�%�@;Y����7�r��8�v!�2
^b�o{��]~R��%UVCŗ%�����PwA"�E�) wr���S�#a���w��h�P�X @�7�X�1�Yu��N�ͳTD\��_eB�`_�AU���0<䱷��˧�O_�y�#����J����)@$��諡\�n.���<v,˃r�6���6S6�j�̏So�/R��xT��P�K0���(�Y��G��È��u��I��:���Y] ���(Oߟ-tc\��z�qڙ��բ�>�'��;\O�H�.
 �
a����GM�wR���� ���%�����a*�AO <�T|`�����B+*P����F��>��9i�[��A���ׂ,�|�Z �,��_
b
A�T��oF����I���[wz������4�ߢl�w�H�uO���0�z��O�Vt����.ׂwG�|�QW����*B��+Y/���(l��}F��������_�Y,�G��-�8��l����]��qelgM�]h�h��f� PS����.�ێ�cz:�2�Ջ��#`�}b�қKd�M���.��OA����Щ%U��Ȼ{W��+�6�����!)��P� %d}��}��b���#6s�}U�	\I��-�r"�N[Cϟ^�C1��pSt@�Q"7bD2IÓ����ZC<�	�	6��d��3��4q�+��Pi����5+��䆹�Q4���[����XNv쩵��K�^�����Z����Qb���^B븁n=AR��~��[}�1�ǑB�xc�-�90p��Y����.D�6�%?�Z�i#xxb�x��M�yf�j<g;?i��a�h8����K��ۇ���"�d�+�%z��hs`���Y��"��Xؼ���m�,���L�iO�,�I:.���n���Ǉ���Tc	@z�v���}�P��	��/�>\� ;�am����e}�ae:�J�a�(<G�9�ܛ��"��ʏU}&�`�Q;�9��`O�KV��E+����B��$�ш���	��z�����/���=���#.�%g`�Z�}KU�w��㌨lm8������_#[~2�:�y}rȄ�ԉ��gJ$�z�05�b������  1RI=r>\z���Y!F��Sc)�/���7����Ԩ��.�@�a�AO����^e���E_�_���Ɖ1M���	!/��'Q�gj#�#��z].on�`Ä���D>}�U>�x`73Z*�(R��[��Օ�##�
�[��[��pC'�IN å<lXF����_��	ZeըN�])�wUS�48W�o�\,�7�/O�hz��5���B�4q���f��;k؞J[:�ܲC���O��T�l�Ny���g+��X>�<9&t�v�N�[�$��Eg����̻����Oް�k�u�!cm�e��n@�<|ğ�-GL��e@/���R� =[�^�r�����]��&�.��ࡀ������j2�^���Q���)���O߹|���%��p��S��mX������B@q��+� ��0�ʄ�o�_1^�{�H�c!F���N�e'��;�$��曆��p�?�;�8� �*�.x�I/")v��5|t�gY��]*�Y���=�hO������;Z"�%ך��U Q�X����H�(�HuF"�@��E�U��<D5D�qu�.j��Vg����^h�+�tAG5c�l[�ʽHw���f~�bc�oReJ@n�=�A��,��CCr���D.P���\�;�j��3��$������鐫�a=��Haﶬ��u���#�w�e�Rې�e��?�Nj&+ ef>2fj�'�n�:�s�:��J���9��7w�gK���Eٰp3)�e2�7ҽ��O\�k�a��WLW����	K�����"��v�6|9%D_����}jo�M�kr:�"��w#����T~FQ�p��h|ы��[���"�lm�����W���=�8{I"��,ǈ�t�6z�Gvzϵ~��z<L]��4`�K[�Qd�����Ÿ�ay�G�K����2|E� �<YR�cϻǩI�;Y���Y��N-�آٔJ��sx^ͤ���8/�P�̚:�̖��i��P��uE��&A=���|bq�I�ɍ΃ǽ�ʺ=����l�w}�~�����B��uoen�I��oN3�,���*��BEwJ����/wO��X�ZP>�������*�hyh����ݸ�Q~��*����\��ڿ2�.)
{	���o�x�&�R����"�ۜ�B��9Yk���߀�W�H^_:7WYՍڍ�1��+�����:x�6���	��sR�2DJ���n3����@���[�x*r� �]�F(�'&�B��%3ݳ�
D�q��,j�¼��q8)y�]T׶0mP��Y���蕂V�u����G�����&����ft�(4�e�C�v���I]�C��Yg�_c�@,�֖P���t��n>�_��^�!c���w2(5'g������ER��ǊlBu�9[��k���n�ā�V��Ќ,��+�^�g.�)n��s�PU����(�YM�9Y�-i�����!�=�0a�;��Ί�!q@�[^�/EQ���]H"���_G��^iEU��V�2�Q6ݥ���z:��1�͏m�������55ˣiVޭ4x�+�<kb���~�%����n���;�`-#�8�y=*ܤ�Vl�ݚb�v������\Fq�m (hm�ݖ1��w�<�L\OC�üds��^��t)%��Uic��O�%��B�v��h�YE��f�OGh	������]�3�P�iw|�Ze�[[cW��{��λw�G2�јE~�S<ɳ�q�f���e\TB��@�����T������cy���Ҹ4!e4!gF�V"X�Y8]�:���4���C�������6�Z~{�_� c� �IV&ˬoϞx�L�H���$�]�ֵ�TZ�+��1�3̘J.CD-�psS}c��5)�Gv���46|Ŭ�Оa�Vԙ�oM&p��]��5o2:LD�t�@rh�@�� �I�$�l�Hk�$H:4*6��� ����R�7+=fŤz�lݫ��/H�5�/�T�
M���=Fo�����I�Ț��� K�A�vX�L����j��q؋�����>�$`:q}U�j'�q{�t8%����65`R�&r�[�&07�~c������¶̯��Y��Kυ��p����_x�slӂ�C6�L���V���>Z�X$��nw������م���^녿�(?T�ׄ����|c/�@���&M}9����غ�:�;:��F��Ѕ�� �~x���F��O�o�뢤�I C@����+��Z���Uي��QDY|4 l�t�ԭ�b�V�g�on�2����ˇ �n��J�L��/����T�F���M~�1R�1���v ���g:(�,F�g�i�)�$�&S'���F��/���qtÁb4�Ob9��e�ڝg���c����~�C�	��d� d�ir�:/�d���T/�F��C�X���s_�=�x��rͶ��3�<�v|2!�g BEaG�X���	R���Ex=S�x�UE��*�m�#
z�'K�@��Z�W�F��9�S� M�|R��Q,n�x�>g
�	�d�:m���j;V���Ne(:?>ob�I��v����{��ư{p�;1�\��r�4@�k#iB�w�.��$�-2l2Ґ��@Z�1m� ��x��?�⇣@PP���|�>1�B��||��x���`�k���'��z����x"�q[�����ÓY�k֑՟�[6dFצ��2W��T�D���s�oɀ2�~R0�>��.9���8ө�c'��V�D�;*�x��J� ֓��n|0QvzQ&GRs
ǘi��#�2�Z.?�c��3
��0�!�:NP���9!4�����cw�L��[v�)��������R�(�����4Ɯ��7�^q���g�v�[F���ʇ�c��6o���,%��Ͻ�>O�n:`�M��w��Rg������Y��׻q��!9c�`�!�����m߹�<3�V�J"�6��$��w��Ff�(�^,ѲZH�CƩ�q/'?˚�4�����$`ۛa]��%V~hMtY����i� 9�[r�F`���2�N��_�z$|h*_2�w���5���پn�Z�5�6SQ���ŝ!�����PN��R��ay�+ͽ`���UPD���n2�
�இ�6=g�rͤ�d��Yc��;`Pi�Oܙ��%���nW]#:)�Y���#;\�JF������m}���+�>��n�Ä+�@�IS�E��o`v���{Ɗ/-JZ�dt��sLp�V7R��xi/�&����T�{�|�;���`l;W��՞���j忄ˊ���A�3X�^�����>�A���?���t��:\D9�_`T+�t�ׁ[?��%[u��6���� m�(Y�~�o�8�mCޜj���.� f�m`q�i���=H{�݀�j�y}�2g��]�1ף����ϗ����qqXk�-XH�.�,���������R�O�)�L�0\���Fm�e��T����aN�t�|���@� 5V9�u�!!^=���M�n��t�e?i:7�(n=f"�Q��%-�.AS�n��r4����i<�%�LiϜuޥn�yb����c
�N5�0���ʻA��"��/�y��H5e�R� �
s�4>��%=pBw���� ^�!���V�����|uw�Y�Dk��ZX&�M���\� Kpw�غ�k�����F��7�"5�E-����`�s��E���{C��v�_���tE�l�=��PzM��7J�Z9�?J,i��I���M��I��뤟��3��(Q�pu_����t)gر��fC�H=��u)?�Q�<QY��g�z#��� �-����񓯝-��ʨ')De�
o|&��%�d�zK0�9)^4��%�X�����cO�������g\�U����$��� MO2��bFo� mosg�c��uz�p�Ŝ�_�M���u>��n��<��������cZC�l�f��I����R}�5��"&N�٧�};o�P?`D���v�N&S���[_�`-1�+��^�6��������{��0��jE�`@r��Y�}��O7�L"r�GY�4B�˜�ڻ �ΝR=4���ϟ���dY�i�2{��m%�zB�*���[�dq�7�d+c���^[��ij຃����5] �|�������ఘ\e*>p-s��}�zbn�K�JU�;8���B:q�M�v	�:,8A�4���8ӸL�o,����n̆�&~,Ś��] �Tǜ��X���!V�Q� ��h�E���V{q�O�V��ҥ��m��]�o:�;��fop|p���\����=���� @i�e��J*5��]"D�J����m
����hBe���qL��CΣ"�^r�R.��W7�	d�/[L���ǧ!І���h~�b��8�}�)�-��=(�$f��Zv��!�:���e�����Yo"�@�ن��ч����o�s�(d>M�i���3�o�x��YVJddj�$O�ʞL-m�9/� M3��A�'C&�!��JL�X�5]�������;�)um\�������z�	����2_l"��$B��K�ݐ�r4�{���3C8��'tejh���e��.ÕD��)��u����9̌�`� E�kgy��\��Ӗ�-��F$1d@���~��u��U�b�U����4�V��c2�x;�-�ئ�. �p�e���P .���&�D�ߞxu�Nd�rc�*��� �G���c�b�Ct�E0�VJ~��(F\��ʧ��$�V���]������6m��sU�a�� �)ѱ�*pi�[���3>-u��kV(��kֿkMނD�3���r�X;���T:7����~Kbf	_�Gk�%�6�6BE��O�u�HjJ�2��%H�L2��1�6���+b�NNhC�C�R�
�O�օ,O�qx㦮��_}Fpi�$�$�,T�����D��-���X ���4�n���:P��ϫȽ4��қ�WS�d�A�#�uu�>�9���"��-�9��o�-�^o���h��P5��é��GFb%��i7x�lX�k�n�pl���DJv]`/�I�U�|u3�`�s��J��w�PMףx��%���2%�2-�ۆ<"��=��[?�ȽO�e^��-��g��B����i�����c�|����yg`e7k>��%�oV�>���8H����
7s�b�CYy���)�����D�u����7����z�F&H_C���`��K�V�m
Z��v�L�-V�&��5k7�0i�
�v!��wG~,��)�A��� /��̉�Or�������6��*���FXWz~vҷ@&���+���R2��֘�s���d�6�Ox�W�[����_�~x]��i�Z6����EO�����U篈�ͼ��`COkJcJ���$-6uͩ%��0춪��R����5t�&�l0r�ZB�ԩ����աqW�&<�X������B�P�G:qG�aK�$b+��;�G����C��/���d�~޾Z�̲���>���ԱTJU�Ș
V:�ŖFG�i���G����-$�:���I`�FKv��Z�۲��d�Dh�c�U������J!�7�"|�k�[��ܻ�&Ѳ��'�t��s���Cwa�K3b��p�(cܻ�uq;�(�8���{�
X�kV��'^��(Z�/�m�w������}A����o��1N኱���9�y�_"k��\F��gcD��w�Q[N��%��y�
?�2�6
�g����'R��];&R��jc!�-��*�l�߷M3��4}��r�������Ӫ�����U��y���lq�*����%׎�N���}�O��L�a����3�����q�s��>����2��5z����T���#;�65|7T�i��Sؘp�e<��O{B���@�?���R�g��@�o*�B)}k���X�l���U�ظ��t�L���fG��-G������״%z�lU�jو�l�����3A��J8�U��!Ə�$V�b��`pB;a��z��.�X(�̀
R��� ��O�o.Q,K<��%��2(�buF2��?��� ^���Q�4���z �����RG����N���M��"�͏�8>���q���1��%�l�^Z0�8�~����\R ߾a�˹�A^�Xiz��a
�M��glTCu��ȒZ#J�6� Vk6�Q�Y���ͺ���8戗���`��{�e�ֆ��?}G/���!�R6כ�
� ��0���B3�龪1�gM�~��-f�$_�U�٨	�˸/�}j�SN"φO$�~�i�Fݽ͕Ν.$X]t=6AfI��v��˅��eq�R����t]�G7�u/��F�Ƕv�K�B����D�-:�j��/�j���(�)�2v[�5���n�>�I�l��<��k�;�{` �zC;���l���[��'��=��� M	k2W�����eůͤQؽEߡ*Sm�(���:*��eUi����N���~��]��ũ�������k ��P+;����B�U.&�M>�I�K	1�r�GR�%��?�0i!ͥ��qm���\zhAʫ�����&�gC�իi5��8C���Ξ��R�G��w�����F��X���$�Q����{!e��������w//ߕ�����l��-��	�R����	:nc'E��&腒ᶭ��|^y{A�q����<ځ5N
�G1\�L��N�Y8]�r�<���n�?G�؆]�m׎`׍|&�L�O���F��`o�	[J~�������i����1��T�B�"7�2;L�
��*�yUeO�فm��ix5R|���a�ȕ�Z̽��l�	t���7��ufP��,+�(^��"��ݵ�1���D��L���;��P�r�B04
�a��G�Nԛ�� �W�@�0�r�c��3�C�'���J�3e��+�}����oZ��1�OS�b�glx����80ei2!��o��Ja�x�nX[:
�}��Qw=41�X#��wϳ�����)����sD��T0f�ٰ�����7o�� .�"Z�:s�W���ef���t��M0��T5-�טƊ[��`������CbnQS1��^����F�;��j���9{�
����}T�]��>��PZ1M_�y��1��M/����M4�k�BH��-2�6�ܦ0�I	@���*��h�D�������AD/���S�Ot�W5>�~�������}�ðg��Qй8�&.�9���A������H�>���S) �P�]�[�1����\���>���T�Ь��`8w׊0��8�vI����i�VJm��`���oM��r�Pov�@�Z.��x���M�`�%?��_2��`�[��������JW&���G*$��(�+���J��p�b�'���	D�p�> �3�[CX �Ka�o=��+���J޺���̠��6��J�G�R���XdV��$�?�=.�����A�n�Ȑj(u4�~�Ԕ]�^�$�]�<�5K���;P��j����0���k��;f'��6��$4�H��"��շ���3�J3p=F��<�~�g`~q��Nk×�0-ͶmʽoᗟF|��PXu�<*�>@{�'p���.���Y���&z^��C�M$�M�rI��4K���m)�d��5�O���&8D8���8P_��Ϸ��4y�A�ȿ��.i��7G�45\e����;/���0k������e�����d�J���"�۴�iޏ�o�lR�%��[���,H}vJ�6cR�PJH��9�s��cVk;�ɴ�����q�)nU�r��E�Z�=9�\|���p���,�C�Lom@���f��\��뿿��^.{~����.��~"�FU�"��Ȣ�-��wq�q4���c�FS�!G�8�ҕ���e�e�+�v~r��7��%c%W�G��e��@�ҝ�ό���}N*���mJ �W�0��<��~��b�L�WI3��aQ0���$��M�w㚀.4��|jd��K�a��s���2:)6ڕ0x�[H�8�;�mu:�I̷�Y�(+�'˶�����ہ{��}D�,��C>��Ѣ���s?d` ��_����d�Z		9E(�C�q�|a7@'N��ʿh��wb��1�ֱ�8` S���?��_!<i'_� �{�`#k;J�����o���3��Z&Bz�)7H�)�K:�)��p�c�}���u=�L�����i�m�p_Cczn"���?��e���y�k��Q}a]z��凰�?�a~�'�{�
��yrFzL������_c?��H1XHgp/��y�G ��Z����NA�V$�l�Վ'vm�_|����_��D�F�o����k������<l]v�ji<�����ACQ4�G}�
zHy|!��<��9�>X�`�ZmrȚ��QY�!  ��P��#6@ܩ7�U~���C���tY�o��O�%�:f)?ǎ����6ܛ�I�����d�#Y?�p��W6R���|���r	��Ѱ�2q&��H:���f��s�@�)E+Z��|������,���bśw���I����LMJ���4��嗍|1R�Zq�U�TC:����/�-b���2�n�Y5ң��3R����dL8X��X�|+�V�4��_����	yfh����bK5��d���DGҥ��`�g��t�Øn��-�3|��ob�����u�>�[@|2i�|�����=��D��I!�p�t�S��"T�vh&���2�������-�V�` �iiX).l�k����[�W�e�!���H%2�%��`�KЗ�[�f(H���8�!}�b��X���
5�	��%ؔ䴜7��-հ�a��}�a���7�c�8���Ua�7;)�̍~߆h�ςه	��e��)�b�E+�e�S�Æ���+9�Sx��Ց�I�M I�/q��+��ڽ�(E��)�'������|"Dm�����+���f���/�[�=6҃86|�dȢ��NE��-{�348�c7_��ҫ����,�!���.C^�ᘉ�|���]B��������^�!�������^��>^KնƟ�@�q`��1�҅���+f	aژqԫA0��*�"_����+ �"_�t:��1�w�̐��C�)�'r ע��6!���Cڈ]q�����x'.f���3��: �h8�Cq�6�BKQw�����i7w]���4[�OvI;��*�0�kvnٌ5�)=��='�%܊��[<@�����MZ�YKT��[�d�/$����d#?l����h	��JdY�_r�Q,,�~|�`R�i�졶Z��6y:�R�$,!�9W�vѭK�0�|�1��+�} �F�UF��CR �\5�n_�����vZʥ���*�>�dõa�,�8g���D_�2EtBW~F7�(Q�$3B��&B��6T����$]]4��m�ad������kd��4`aV���l���w�$��-�.,)�W_�b�c1�@�_��p ���x���EI."�V�x=si�>������A��=�Y7�I���13=c<u��8�1�M�;<��-�ci���Z�nexXB�;<p��'�(�n�3 ��B�LS�v3S����p�n ;��{�M��I���.S�@@�q���C^��ی�����з,>�fA8��p-tM�m��)���U��m�6�A�!�� ��K�SǤ�y�����WUt��U��̝���ܰ�������D��"����d��Y���"�`��~Jq��og�I8u�Az����
1�k6
�}�
c���o��T�c�{��?���g1M�~~t�mdo�C�	��B��B��o�ҭ%cOH�猧͜�4_��嚎�Q�����7�q9}�j���s۾�c�y�"�#HjW����)x����?Ah����^�0*ۘ�샐Y�\R��S�z���s�_�P![����y�%C���'�ӦQ�$��D�i��Z6�E���R�@r��*e�	}:n�9T5>���v^RK�Ě�'��;p!^�U�J�5wI;�)�q+�$Z�F0UL�>��H#g�1B֡oS�0�$�O���.�o /�DG��^�'�ͯ]��PF�����DP���[�ƹYY�j�,�3���>�e"QPgI���ɔstBfqJ�0@P[^��7�jc�u�6}Ȣw�F�#�|�f��6����{��v��rq�t_�W��Xg�ZL���˩�/�����w�����WH,����(,��`r~6\��A�'L��/�(���x*c�$��@��M������
�;ڞ>m�/�G���KEH3.s�� eF�+g�u<c��Ə嶳٫��Q�}9k�bF��q��6�����Z��M�P�#�7�+P��HJx��rG����j6��}e�#8�7�{�UM���3�j��������@pd8�0�l2��=��{}���W;��+�+�;��&{��n�:Ok&�1\/2�����"����t�͸N�u�A>�@�m���Uw)#uǨ�ٱ,Q��d�~���-R1g��v-���l� ��z�VHb����g����z���̇7�{%��3p$޻w����T���K�>���d���J۪�蕛�-]Ug`Z��6�,���a���B����P�6}�
����f{��)�_-�#���р�8u G�n5e��=L[dH�=���DU9��x���M��$=h��&o��8�JA:��x���R������NZ��Yc�7aDߝ�s�5�dn�~~<�yCV�oYr������Ħ�Н���o�9�8����{¬��G��� ���#A&hKXEyo^�MS};���(�1܂(ڸRt^����h�Lk��#WFa��������I������:��v%'�x/r���-�۽�aaI��[�sm39��wk���4c܇I��䧰,-���|�����A�&��r����ag�?x��j��0��L�Q�Q�O#R��Ψ��]/hn#��Ƭ�1ڐ�3����,Ez�� �6Wh��%��M,�|��҆��'�B��:���f�'��$�3>���,����^���>g�K��(���QYJ;��SAt�5�U봷P���NR�B�7�تۍ�F�}�ݎ��RAb���a���bo�mq���"�/�oXRw{��`�`<�[W��ifz�ܨw��Ta�L����D漆��d��	"��@� ��d�O�X�Ȃ�ߞ�!�h��R˜L��T��ڹ�pBY�kK�*�^� u�X�B� *k?ipM�6�d��8�O�;���d�G0:C�9L`��s��ǟ;�1žiW�X�5��������j�7/� o�*`��~>T��S�G��������~	�,Y�}\Y�u�g&40�v��`��Q�b
���r����#��FV������+s��W7㫾�iR���Fk�:i9��f�w�Ggn9�IE�����
>F�RD�c���H�w��Y�!��Q���{��QG�I"���X�������6�^4p^*ϝ��
��t��y�v�DI��vjdht/x�-߰N$f�����C�̧���j��?�.���W	�Tڦ�Kə*�\Ό)����U��"�V���o����s�X��;Ik�xUm/$.�v��|k6�6��'��S�1,�ÀZS�݁�BoU;퉇�1�I��\�~��6��Yݲ��o!�d|x�EgqWC��v$`��4�ъG���w�X�#�Ѡ�Ġb�`�y�n p�Y�.,�x]т�w{�t�M��b��zn�N޻��r��m<y��,�$�x&%�XӸJ��%��`@?��'6{�+<QMv���,)0��O�M#)��N&�=�vq��$N�m���\"�RS(�g8�-���9aT���L�_Z�YGD�],^:]��Dn��<���d59Mk���{o�P^p�)r�3��P��
���#Ә�k�ڗ�dX8h��L>1P	�zFb��܀ A����6�.#z������}d�n�	ܜ�e�VY��R�%�IG��w��C��h�h��@�m;�z��i��^D��?.�Ӿ��.�\�JXy�@���$/7F��HѨ�OEYdE���*c��%������zQh�ȁ:k)jw�O}�?�B�5*t۪�]Ij��J�^9�pT���T�,����3p��]�@�����.��$*�t���yC��2K1��"M��?c�z��U�A�/|�p)��FK��洪M�-�t���1�\a��6�R�$G`�<\��� ��Ќ�"H_�]�8��F�H����'��
���@��	��z;Y��|݉?p�̑����"�b-��w���P�wҽ�D�?������/x�M7��A�W%�"����U�`�U�Ś�
���+_��7���jόX�-b�.�)#[W0և7O��&��.�P���U�" G��θqc�m�Rڹ�����q�|�(o���:}�D���eb��	�Q�#��FqPs8ue���5��f4j\�Vӌ��,��KCdn����e/���~ڻ��ɣ����]$�*kO8\����{�����:� �]��%�0ԃW�Δ��
����V��?�켨>j��GUxH���X�+h�6�rޞj�j �57���7�~@��1��!���և~ۥ��.�zg��Y�s{9`F"�h�l�1��s����	�J���hŷt���ښ��2�j&g��ӕ�2���f���M����i�L;r���H���o(�#%E�]�'��@?����#6�!Vv�>��מ�XN���oM��Lq����R5"r������~�