��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ۧ[���B=PKx��{�Ƈ�����3��[��M�>���.�|"H?�E�9���iͯ�;�����UC�	g{���u��!|]���D����5�[d��0��N�n�;�C��2 �ϑ?z��`8	�a�c!E�����۵�.�R�(�%��5tU�h�")y`����~���ÃCD��P��1�=�8�Oc=��5`NE�'�:�w���rC1�C]id7����U��.u�K��9_-[H�@���:�d��I�׭�TbBQ(��]��N�+�T����=ջ0&���Z�Dc���>UB�u�w��b3UF�"�k(٘FY'��/8L#%�ݱ%���X���n�S�pZN}�t��)�&S���k��X�k�G��A"w�HzFeKm(0��UB��t)������Q�;���pr[!w�\�2�Z�I=�~�*:�R�&�P��p��t�<�樨������}'pbMǟ���'��b�oYJ��گ� ��P�j�;ju�x��@*A݄��Ё�<d�H�G�Rj@��⥸s��X^�bJM%��_>�=-�Rg]-to�-%�����SKRp��(�?�Ƶ����_��,�-�>��������u|p��Z�<a���<���/ܱ�N�de�q��P���U�%���ۢ�����q|G�9�ķ��sq�/�a��6���:���N1��0=�TR���g����h��ԸI3Ѿ�y�s	p}�+�V�������-$�*�RMrҢ���%������^��Q����}��Ū#�Y�.Ee�x�vt�." %?La{��ߵ1���!���B]Kήf�x�|��vMtS�΀+).:y���C����s N��z��b������u�u<S☂u�9LuЪr�(��ڛl�^��~2䵐�[�v_����	[]�_�X��+M:v�"�w����%:}�z.s�a��1�Gﹿ�pI�I�<zz>Hp�jsa%�^�<ʻ�3Ir��,�߃s�D�)�0����/���^��]���z�0���p�t��3@�C�7F'_�hPdW��omоrS!w���\`r Zj�N����Ӄ!�'K���o�{�l��Ɛ1 O�\��')0G2d�ߊ�;�:�*��A�lF��`S$��֙j�����5���E�M�3M'�8�,댛(W�[��b�i!������1hc�ene@v����'BkY0�<���L���*Y�R�A������@�_|pF�5K�Ը�!k��QӨo�;�9����Q�/�!��ᙻ�.��=0�8V��xLAm��2�K��O��{��B_��e�2��ؓȜ�������&�js��:��Fۋ%��0�P ����y���ʿ_��v�ؿ����CC�b��&A$|�t�5+�k=���6`��Q>�Dq���G��+lCW�D���`��㒂(��ʤotl{�����0��oK�<�,�����ڶ�m��ٿ������%b�������M�UF�-����V}��l#����pͿ��Z6{˜�o�i؃�f%����{��4��� ��c�ֳ2�<���{�g�bp�ї�vy�!��d���y�\bq�z/��7�Ƌa�M	&��$��+�Yn�ӭ��2�o�*c��1�IcIR���z��蚄����(ggW)������Un�i�����s��+��J�*Ȫs��y��^|ʚ��"�b���y��"�d���C�%��FJ%�*n��?��tt��@V+��5B�y2��&�.�?�{e��5(�}p�h!/m���~�|[t׫~=p�7,���X�68����gPk�D������r|mQ�;m�%�aҿ�>abing�?
�l4C���^+Y��#��z�к��X`ӃSҩ�m��߃�W϶F`����؜��A6��\�Ǡ&{-�[��x*`��"�
`ߛ��U�������N]�w)������Y�0HH�����E;[:g7L�
�N�DXޢ<�b�6r�����{d���R���Pീ��T[�� ��r��}��F9:����\y�3փ����U��byz�-����!e�Dk&,*�΄���ׯ(��M�y�-|Ʀǚ�E�/�4{���&x���A/��X1���:�s)�&���R��l@2q&��]���O��k6.K��;�]�Va�a���il3��?f�UĭN�|�]'7Π,M5?v�Ҫ��%%�ʐG��-��n�3|5:�Q�W��i#wR���fZe�4��}�4�y�} ���<3Z^#+��hFI�R��>��_2	�j
�#�PoS�4f�����>Ii؋��������������
�xPtlJ`���rT�Ƌ/��4�csO�]�@�~�a-�0E��Y�s���4���6�Q�����S��
�����δ���|��j�����x��-�C�{���i��ĳB�8"$��l�"����c���Q��&�$�3qCJB.����H��b����J�{-z�+�[��+h!�p
�Yw\�?=22;@�=6�n��,=r5��ڿD��<W"#Ad���ͻ�5`�:�L�P��Ƨ;&��8}���%�@��^E
/?�1u���h�ϖ��3*�������e�݋���SI��Ihk�s��8�2���vXWr(�DJ���
{��>Aa��d	��gS��o.r�GH��Bx�(DgD�����c�w�iTI4Oj�+<df���)�lE��L)b^������@Ji�PA�Z�޲,��s���>��:���yʾ���(����Mƅ�ᠱ�&�; �+Z�}�Z��X�ɒj� İ�"Ax�q辏0�&'�
𐜕��,M&os�t
�!�� A
�=�H>K���f!x�/�39��
�t��#EuG�훞��l��s��!!�)��͌�p ��ğ
[̞
���d1_�,w���u\S�"���
́�95��2�*��!0������W4�Kk0��#8��4��4�}�U�Б;�-���Xc�/9S�)����ۼ(;�Z�~*W3�=|o����y�!�)�-��Hs� �_^����ajR��PP#tMK:�r"}��ʝkb��KdK����N��q������6n|��[~�6�.'�mƵ��BU��G]����*�u"(�r���SyUL�������Q����E
��+uq.I�h�ܕz�7�"�"R�c̢"�{�;-����c�=������t��ikn��#N�:/|�3�*2�\1W�8N|��&�ѱ[6�MP��I��<H�$��@�*�'�
%T���\ڈ�ɰ�W9#�+
�ۿN_�J(>��lg��[���]�SJ�AS+B�s����|��o21�z@��l�����CT��?d<z�I�Ѭ�Ƕ�(�؊;o�1��32����9/�^G<���ף�� hr^sD��j
S���*R����^P$A`qk��}�~-�{�[L ;���b���⎶9v�'�dD�m��$�˘�J�S$�+���b�C�iȋ�O.z����,�$UKgk��<���p���}�Q��a�`q�����D �n���pw��Ӳ��a�X�@s��;[�F��5S����p��^sUHu�R����(��'
2��(M
Dܗ��ƽ�ʺ����ͧ�v����x�'J�n�'V6t���˾��*_�� ��B��ֹ�9�kk��CU'�~HzgF �7S-&=cw��Z�}1zm�Q�l?�п����.��md;9»�K�x��Z�$k����o��/�|�Z^7!��\�e�O��Qi�>2�)3.J���-�gVȸl��B� ܹD�jk�P�Q8�&���s��*�����&%��Z "����/�%q��i�	��1&�D��W��e�a����h��`�ig��A��ҽ�΂ʌcku�2^���/C�q���}f�<x7N��-8���
��Ͱ� ��.�STK_B�{Kj����-uq��FP���u��;BѸ3	 !�vq���$�&�tG�������'��L�
�[�|�繖���߰����r�8�6P�l)���%�����v�kL4�·<�В�i�NadR�l4�N;����Ob��[<s	��a80%6�ypy9�^ߝGW][��.�d�pYؘi4��r$K�:���c����Z��M���F]�D�} ʛ�-|���*Qo5��<]�m�C���y���/|��y����$��,���
�.s��N㣨��O#@�JZ
/��Om�o.���A(F��@VJUFy����[��	����,*+��.#�Ҵ!j!�挳)��ti��]����b&�+��&�0c�WsHl���P�]'�˭�6�xv?䯜�|�4��<jN&B�!�ufG׃R��㪄N���8���>T2cv�_�G�=O�6��(FI��Z(�CԘ��,�`()�G�O������L���v�<�>b�G�C����g�Zpov����M �U����T���|��Y�y�@m���R��q���Jl�x��`Η�qQ#�/�Q�ME�~�!�`�.H����������A�� ��-��nC��r��@�r7���Ĝr-�,#Q+	h��{ȏ�L�'wU���k��1�����v��	���kUD���J���@⽆�p|�u�_m���%����P���W-9{�;�O�����_����<�r��v�t7 A���~c߻�#��iT����68�MQ甐�๼v�b�!�~1m����{e!i�ZӼ��P����t�=��+cZ�.�х�-R��sDP2������i|���r	0��jy�a��T�3L�߀ C������ע7��`���k��:�����t��^��
K#f�1(��v��ɹ;SǰG�K�5��3uH�1"�+iA���N��_Yڰ��N�����͘fw.E,���Q
!�wm��:~X��S���l���5�A����k\C�}�k_����1�k��N1����ԝ��X��¸D�@�4�����3ϳ<�2!�N'��-l��s���t,=IВ���_�G3�[�R�B�N"�p�� ���1	����_|s����;�J��?� ��¾���%o�Ǘ~��,�����T��Y�4q�t� �^1e�����n��HҎ��R�����>����w���x��c���� T����;�0��e�FT\tӋ�iy���A��$�sfybt��9v�����p�7WZ����
�I	2�{�90H��0���O�*��=0n���b+#��{���S���2�+� ͆�?�Ν7h0�+z��xDv���!�M��$� �J�/6����wf��1Qi��E-i�����H�?B�����!��v�'\�OF�>٥
��{Nx���y����L_t7!A��1U�܀��~&T�ק��Of�
�\/�T��M��V���!K�$h�ғ�x�R�ѿS�Z�+��H��AZ����X:�uY�)_q�M����%��hR��S�����2��9'��Gҟ� C�ǵƺϞ�pP����u.\��ɆN��|N�Fx��XF�&b�,��{��8��ɩ�;����< VN�;q�1�yJ$����
��rBD����]� ��'L�	�1>6͜�5#�󪱙�����|6�4>1�m��k�~͍�����&��^�#6�$�/H[T��i��6T������9*ֺw��'xVa�I�Y��7+�k�X�A��f������$�G��ğ���8z��$ߺkl��U�*�b���~����JY@h�D�����T���!�;$5\�;~NR��<�\�N`�{��,P�ۯ\��ݧ+K��3'A�wq�z����󲒴�(Ml��,�9q2�>YB�짴�曪!��jsE/+���� ��f+�\����kX��.�y,R|�����*��]9�F59i�O^���3��{����]�NKw(r���]%����3j@�`آy*�	�tLs��J}����ޕv��ƌ8>��Y���2Y҂�������	zY�"*{��_�%��ٺ�����k�"r��D/��@����/6�!撍�n��3�g5.ĖE>�N�� _(��LI�4�p=	c�=�3�;6�m2�F��7�����f��T;��0*	�+<����|��}~���\q����7�|����&ޮ����.�@yI���m��|�"ȅuю%̣��|�%�g����S?��h�O��
J��͐�y{X�,k�er�$B���h(�v�B0��S<70�3V����G�B����N�Q=��/V�T�d�E�R?����u��B��u�4X�E%��>�6�w�r��r^��^OO��dZ\V�$�Fu�o�vd�J�F�u��ʪ#����P�ʯ��(=sﾸ?��VH<8Ɠ"��ޅT���Z�!ҷJ��}[�$�	�N�gȚ$i�z3�H=֪60lK߬�I�(>o'�/�q�R�a�e�8h�{��]�c�Z��vX�͝����m8�F|P��BU�!yA��ܓh�$6g	H�Sx���'�K�*?lkth�%���ԍ<l�)�;�ɶ��ZR���ۛ��=���m��n񱘡]!�FD�M|	M{�w/30�_K�F�9㲽<NYI���8QE�o㲥at�}ɥ��o�-�\���h�*U�8�֎�����<�2�?d�	D)k�T��r���V�4ׄ��ju��v8"O dBFB�g���:�j��p�]��A4���W�*v����"��<��T^￑Zt����d�9[��L��|} �\�� �$����e������{��!c���<e�n�pcP�Lh���7�%�*E�_ �l�~�Ukξ<�ȨWnB�u��h�ۣ�Ni"�$��w%����� FS�am}�9���As��=�P�oy�x>-�O/I��0𯍻�oҭ���FEl�\�Y�@kĹ0iJ��}L@ׁ�D�T�oā��.�Fܘ�ymZ��J�L��Ou�Wd��7)��b��?�.�n��x�잕�8��`���~N4p�\��n!\H�~�qL�.Y�;4�X�R��G8[�O���N6�$2Q��9;�5��nX�F�c�#�����{~�;�s�`$�)��R��_�z��J�����	AM�RI�jRK�Jq��,���C�q]�{:-���L@���!Za.�cpV���A\���%�Q�������t �Pc|;8��kϾ>� �+��Tƹ�Μ�n���y�D��1c/5b����y��%`r��M�c^==�zi4P{�D��b��9�KE'9���wp"��s�Bj.=a�3Àl�)~!8Q�L�]F!X�m�@5���__d�T���1��.!B8��ϵ]���H�[��A� ������*\MWa��*�Nh�֋�O��v����dv����:6���S�;������T��ƶ:T|��'C��Y���{'X��σ.��O��o�Ĭ�	���lc:3�a,�6>x�۽b��s�S�Q�W�{}w#�7%_��b��)���-uBuл�`���b��+S�.=6�N�X�F�*���z���ɽ$>�T��IR����Z�v���+�-���� �GO����G��	�Ccވ�	E�e���.{5��C����)�jA`��c)��#9���ܢ7�ۗC�GL5�- J& �\G�/�D�����z� (�sj��ÙL/�R)d�
u�E�luŮ�>��8��"��5��~� ��= ;'�~=��4�w�meC��yX�s)��p⌸[+��H��c���Ʃ�����E�B?H��q�D�Ւ �a��޳}�~�e"����mi����=�<ny���B�Ir����m�r����o �φe�e{���5}�L�ȯ;��أ$����z?����m:l�!�9kq3�%���5(R�MA�.�A�}�?Qu��\*�Z�q�w��EA Q����3v''�OM<��`����Y�$+ۉ�'���,�R����/�
<?@�~1 �1(�rx�m�r��"��N#|��W%� $S����M����Ҷ����B�<�yc����}��B�T��ST�=�AJ��#�����ˉ�]���%��YMi�Cy4�k���oh�<����{����>�2Y@�k�&��8�����jVQ-�ߝ�D�O�tjP@��ՕE�P�&Ҏ�:?�G�Y\�KP�:oT]��a����:v����x� ��ܥ���]�w���6C2Vs����J�i�(��{��D�W��ո�_֯%�$@p���j��	���k6!M����}�/�qԨE5���P����<M�m�"s�h�>�7���/�SV|��ī�"�v�圆5�^B�Df)%y�9��@�M���X�<���ȳ��1%���込�������N��M/����Y�0��$��G9l-$=�|�."�����R}��e�W�� ��+1���u���^Tb,�rz�O�QRg	��y�|֦(�=�`�ā�9|x�?��K :����Y0;�VI��Q �?����6��C��G�8m.���GZ�K �;uߕ����m-g}���`%���B췩�/(��d�����i���/0��_�﹐��v4���Y��x����V��5;�k)��6�������]�[��@�����l�tDI}.Z���W�:?Lߠ0QQ���#����`�k��_^�p�����%?g�n 2�4�@8��~g��	<j��p( h�V�T��)BE��q˽��8�L�!w���-�䔓�w�|}�&,ޜy]��E̲r�9��������ڌ���f'�63��K򪨎��YPA9�\��@��h�?"r���]�s��b͒�
��H[�D
�+��mN������:������#lu�;��\T�������>?Y�Yp���5`8��Σ�f����Ғ0�qEg�@r���).^�'�B#�
fk� ��!o0:�l�틸��2.�-N��*�%7#��T�`m&�:ǚM�j�Љ�V������BNfkt`
fAb�*�M��Z���ds��33"Bd����0��+�.i1���������ͭ��4�s�p�7~�� ��BP	~��L�����&0]Z�ɐH�\�/q&�0��[��&WۤY�<J� *���q�z�`�������
|E���@<x��[lc�gQ:;I-M2���w$7@�#@k��ԫl��r�����]n��1����IH�ۧp��O�ڋ�i���2�쎐���4��t Sݑ܋��B;�&ߠ��5(�Z�=	�:;_�R�.���|���<cNJ������|�!�Z��LNR_��wN��:~0���)�fx�-> ���c��䰝^��&h�3����-Zj�԰�>�֘�u���X��#,3|�T��E�� �LN�!w C�D�pt��3�U<~QP�/PL�z�(��^C'���:�Ω���B_\��F������Ա��v�y���*MU��y�E�$�U$�d�#]���g���=7y9��!�H�&gaS���孙e������OG�W�9dC�!����Aײ�fD���bp��U�J�+UR ����W��QQ��m���@�9�_�J,[��4�w�ye*�0���?��EQ�%$L��˭r�%���$�6�9Մ�y6�����wG��M��wy�x�rR���m%�0�Y_����;�ֶ���oǜ�dK�Q���)=����d��?����B�-}���2�ߵ����,�	a�9L�ɕ�V����PÉtE�~+S(l���4�0f���a4��Q���vE1s%�(�h�:P �w�@���T�c�}Կ���[T]! S�Mu������M?�D��s����~"OÅ�fN��i����s$kP�yz��3|,���z�=eW��& jF��Gq6�Y�jw.�R�V�%"�Z�P8��J:�Gw�81)#�{�\:Z;d�Ǿ��&�}2	^c��kG���×
����e��dd��	�{�KM"� �\��{�'_DI�эj���jlMlIn�+ka��BV_��������4O����T�R�h�
����IJ��ƥ�HV��P~�tϕPb����4.�����P��ٝ�k��������rj�`R��c,:	��i[v�P!�+%��#�P~xB�X��#�JVg�-��z���&cV^.@�ǻ<�)���К��C9����O��0��۔���|����|Zb 軴4��@�w�u�]�Q�˓&F�TB�d:GA��8�̩	�� �U�:u�?&��P
�9��*�ֶl��G2@}MI=�~1���*lq%}{u�T�/O*�j4��N�Hs� �}(�����o����E;�eB���q�yD��u#yhu;��'^�+�U���:	�t�^Ѣ�h�3}�|�CZ�b�c>����&U:{��U�i�736a��NL��S�H�@���]�.�A�(�YVn�%@u Č���uFP�D��[UC!�7iǑT�KIz�(꘣;�P��k��O.�]�X��&��{��r�� +�CQ%#��A��S�-l���T�������*��n�>���Ҕj���.�yW�\<$@{�x��i��x-�����a̬
�ڛ^hR~DFx�`|o����zo�h�־z$NH�bٳ��k���_F"@=/�<��<Ŏ����3�pu�p�ͽ�r#�! (~�i�'�\qS�]�`���<��,S��F� A �˻�����bU^��sW�����9ʷ0�CQ�F���%:��d��V�s��Ov��5���e��$H���Ǯ�V1��䋽�
�P�|�{ �u��y��R�ݘ����yirI&��^��x����{͠ћ/��uͲ�/ڦ�u׸"]<�V�F�e��`R+��V�v�c��(�̷5qw��~_�L�Nt��Y,]�pE�	�l�4R#�v��
���u�5  0�cѾ^:jݵ��l��Е��9ҍj�y���f�TC��q��x�r���*6j��dO��2�Yla��h3§?�V�6�� 쒽 %g�5��\�b��5��
�
��?��㹘R���E͢-������G�����i������x"kY�`�˵<v�����s'ꐎl�����t�,��Ⲿ�鷼`Q�CC��l����H�B���P��=�0�?}2�a(�vf��h�#O'"� -�Ef��T�Q{�ϩ�y{ĸ���d�7v��W*y����M�Z>�mxH�p�RR>��$�*~���@���,��O܈X���Ūه�&�Q�Ȣ[7,��L�Y�^�A���L����*�ݲ�y��en�+z*�k(Sn֊���3���p�T?:�B�S���Np.�F�P+�@9����2&]K��é��{�삤(E����	��id1��Κ ���)��C���1����P+ �p��a�2�1s�����h`�xq�ͳ۹Z�m��W����ju�V�j������S#�+Z̊_�Z$�)ؿ$U�u��y��.�:2�8��;YUB}C�����9Z,aR��A�����|�=ծd�y��߸T�����V-{W�լ�O�����w�[%&f��'"��T�#��?��un<�O�hb{�A�v�.F���?g����E���mH{NW*�ѯ�`�>ڝ�z�=�銋��/���4:z��l��n�;8�����$l���<�R��؂Gk�ɼ��%L%o!���tyu��B�:`v���kjM�&����ܜ�o�s="�]r�ld|�a�8�f%<�Cr��叙��Wͷ]�%gE�ׄ�2��������!˘.�°�c��/z$jw�U�@���gq� vf􃈉x~���C+�X��UQ�;�R���9��$c������ag�T���Ƃ�޼�)�+�9�V����E���<��V�Z��!	3w��	���(q�u�B���﹢{�l�Y�V�����twY;��h�3$�J��q}�q�B�d`%����/v���C#��[�ch�u,��%Y!���ǦHܱ���)��N����t�f�����1J�	{��J�]�j�C�)��ZEiQ�E�ӼJv�'t����M�v|�^�J�%�1}�i��diıH�ɷ�<��:�K�!'o2jNH�vœ}}.�Pc=�q1�Jt������d��<+ci�7h�w�_���rՇR�������@9I��#,A)�@^�t��xd_����ο�ǰ���0��ެ,���Iˋ.��r��c��)O{�\�0I���
OOwY^���o� �W�z����~d�,_ZI.�o��9��3N�)4��^_�G23�L6�t��i��G��O�� ��Q+����rs��O^�T��_�gYlX�;T^�x<��˪�`/+�Zn�W�i����e�5�8�(�צ]�Cr����23^WsRP�_c��� g���q�u�鯉���d��l�}ʽ�Hk�ULҮ&�0<�jͮ�Vsb�G;�ۡ�@0[�]Sn@l-d�iۖ[��Q���[�I�3z��7M�P�F�4R����6|�sݒ)����\JQ_/��T�M�/��;3��'t�)�P�WD9���J՞��D���nR�̎/8�Nx��������Pt�ސ\�Ժo��'v*rG�@�dU��(~���>!��8�
�VōA$�/�j��j�=*�N�qԲ�^�zKRE��*��t���E�&�k@�]�Jʡ8�Ż�ĵ�����^�U�H�{��1{�>�|�߭�^<stj�+��4	s�������5��$�y�5(�wO���c�g"���r��׸l�(�u}i�6ܷ�AFޟ�w��A&���9�{=�X��*ˌj0��]�f�e��3���r�s��K�����eJ)�X��o�uZ_�t#�����vYp��X��)4;�6t������X�^��@	�mq���Θ�doN�.}5Ha��  B�k/���N|������v9�7�w� ���@���)@Jلu�G����'x5�t�r�m�C�#�f,����'�r�"�w�:�iV�xߑx�I�%�͛�!ٰ�,�_�!7�n�ؠ�w5�,�����Zk�	�C�ĎxБ�]�¤`ܧ~��e�E.������tq�����x�,?
�pMg_�3�9fv<2����e���{�/�:E]E�}kY����U����+�Q	�A����"[��ȃ���S �a����Ѿ��(��v��cN6�F�٠Dv��~�����9�þ�ֶE��G��2Ҳ�E$Ow7�$�
�ݳ��W����BaV�E.��tSȤ�	)Z�+��g�6��B�T̑g��˱qwnk��y��zBG}�*+��R[jJ�_��3�7��/3+�1�	rۢ&�,�֧sc�ɫ'�dPS�\�Oy$�����@�U��~��f�ؿ�B��S#!����ՒQ��&)�s���!E:6�j����o�N������i�%��p��x,�6wS�h��|[���t$B}��f�H�H��A�'/���;X�	ä$��7�s̑wb�u}F��o����Q:PL��ωA�-X�/+��8��\��Tc�|̰�𯗠;��^:ޢʨ/q}�� �$�
i�+Ƒ��U�y?J�>w�?E�uW�)��9d��Rh�ۧL<�����Q�U����o��|@)F@�ߗ��!@��%�OA�T#k-]sHu.�~p�HB�Y��6Ky�kƃ,
�/������^�������FH>�JR����C�ҩ��T��v�B���G`:������0#�dMĝ�'��j0X�b᭐W]�V�4���#�������ι�7��K����p"��C��Zh���!��TN�4�'��{ŗ^��G)D|c�QM�InF����p���*VU��#!���DL�ꑳ`�B�� ����0`?�����_�afcE�P�(\Ѿ�8�B�.*)Ԙ�Z�2�br�$�/�p?"�}$���T���=b�5�{0������Vo컈����K�Q��tÏ֣�-�m	�8�x�&DB�U�5�Xt�G5�Ō�7�������i��u�KbW)���t����X/�4�o\
/��&.[ 6���.�Zt%���%����L�q��."�����\"�kY� ,�e O�U �܉t�Ԋ�*W��_d7D�ٺ���=S�������z�g�{��b �{��T����|��L�`t��sof�1��,�4�'�v���0ipv�u�Sa���k
���1o�E6�A#��}`W�?�µV���K��*7�M �udL���Y	?6��ҝe2\.�@�I+T�o��3��S�OB_X�	G��=��y�8���I���Ol��e}pJ3h��;�����ĵ�����5�H	�f
�<)�=�����1�q���0�����?���v�HF޹�Qjo!����"�G��c#x)tk�>T_�rRp.;^g��\PK�EZHశi��.�,�4�3�/�l����]9�Y�^J	�J잠Q�c8�f~#{?))D�6���ڨ��>2a�+K��^[f���	��?#�ȣ�Y���YM��)@հu�����$�F6���������|t�r)��Z�M�=�f��:�Rr0{pAJ�ٱ3/V���d���\��)M��Z�� �F��!,��m��N8v%�T��$.-�fZ����,2*��{<�r� �.�j�7W�״f�C��Z���-��,��֗�g����QD����>e�;��Hus��"XF�N���w���t^7:^!���KR�<�eq$�7Aδ����3�Mg`�,*�m\�Y/�Hk��=Z�r{�3ܴ)���6 ��y�eQ��ιb�����R&�٩j�Γ�5���2��Y��3.�)�+�j�z�1>�����F�<�i���9�\\�n7�Uב�7~2������g��Ćǂ���*�q�슗��@MMfo!��)�b4pb�s��b9'���B�8�8��l�n��K����C�k��0n
�����b���	^��:�lv����Ҥ)��T�l��w��8���x��p�GBE�=�%�d�������?���u����_�ZEz|4�$Y���P���������ψr���JL �XIG�LW �l@3����1� 6��5�=�7���Y�SL�.a��V�_�l���osJ�����c�hPJ���l�Z ����"5;���T����"?vC�{LQ̨��Y���qȑqe c�Z��7-�]t<��=�L��UqqE�NDyT�P�#~��%�~�=&� �MKY�m�w;a{�߫�U� �'X�N��	�p9ߴ�=��PJ�]��|��Yd�n��Ԓ�K�#*er����Ro����܉ġ=m`��T��R���v�U��c*�TQ�;�9=�J�k}�*�����Ac(�^�W^��6(u}I��ndRnN��<�>�JT���E���o�l`��`����sI��e��Mh)��%���\`�DQ�d�_�¶��z��#�Xm�UtT��Cy�
M��_&in2jʈ9ё\�Z�2�?�(덁s˕�Z�Qd^!j�t����_�A2ը�?U׿ؑ~1��4����k/����o�OD��b���g*��}��W��!�&���ý����t@��{�>z��`s��"@tPh�k�	�F�P$���b������~6X��3>X�s�)Y`��.����kЪ��`���^bkM�Ѯ��1�-�@��9Ѻ�W�7�s2�yg�=8��l��Ƅ��'�����̳sc������\���%)�,0��v�,��ͳs&��k���:��<�oT)˴C&0e��.���;��1*b˹W�Q��/T�Vji�s��k�?�㲎7�͑:׏k¡Ie�f��r��о���Դ�����4O~ �rE5�?��R6�!�D��j���}�o�N�!H~��d �lǒ�%4��*�ƺd��➰��?t���4��p k�������r�_NI#ct;6�@^۹�ϻIs24�]�=d���ac�L5 ��}V�I�*���c����� 8������mڭ�9Q%�^�֮MF3E�������8!0�m���|��7�Y�ޟ���=�gdT煌���3������$�|��9g����	���� ��db�Tm���o�e7�ߋ�R`��햪�>��3x���rY����BF;����_Ǆ*(���)n�[	�3�ct�Z0�G�Z�F�s�`=�hP2tF��G�
�����ě�� l�pXö�����/����`��o6�u�X�n��p9�D���	1��Y�L�G"K�X���e����w(�8-��f��=V��>�CY�´t��t��O k5�ߖT1XS��A�4�T���2�qU��JcW�
�a��Rr�V~{#'c[�#M�(E券^hyk��0�z5V����+Z&r�$bE�;bm{����!0��i,|ʞt0�h�~Z��<��0��D��A�Igng����j�^0�b̢�h�jӫ�u�]9苞�[��j.�+��Moܒ�odr�N��Eh���c����� ��+��yc^�-��i뉩K��
Y��p�>����+�*��d��Z�3inn�I���
���'��ѳ�C�`�<ٖ(���Ft�/�#R�T��g�$�$���f�=�fI4�0���sn#���=�-��<�e|V������?8����H)� ���E�*��d�3�@]�Q����LNw�7c�<�'(����	DaKHe���-.r׽1�* ^¥��K~8*WQ�h���v����ht���#k-FC��~���qă}����s~:��H�5� Zn0Px��ފ���3��o6��D_���u���-oe������>��s{"�̫z�=T�x�A����_��N��P�^��(�On=�{���\��_2�]�w�a�)o�5$6P6e@����ٖ�����������N__��a�"��VQw1�L��� ;WF7C%�B���̔���8n(KZX�!A�=������ȏ�|��*9�߯ˡ�-��5̵�����evUJ�'HH{C�ڽ?�Z���m��p^=�j$�v1[��+���߶@�_�G����z:K� #\��x����?N�ԨRU��Q��k1*���E1��=:��Ո8T��k�~�P�����p�6����x��j�C?���f��ݫ�;��U�EB�t7���Hs�Ä*���m/z�t�1��T�9��l5�4�ᢈ�� �h(�����>�JOU���:p��G^j���H
��Y�(��d'��WȨ���#[���3�Z ��<m���u�NǃoS��9)�Gߚ&n��׳�oy%�P��!�R%�@!�<��^Ǟ��c��&jH6�;=�!n��4��c��p?_�A� Q����'VR�HT��/G���/^2��C�w�� ߸��к�+}�bN,���ع�_�=����X2(�02G9���������7�j;���oA�L~��r�$0#� � ��D�,R玱:�����b��3�r{��k�0���:N���~L����ق��sy��J;H�Ls��₝/3x��W?�An#�"pzE���G�?8��՝�[p� ��M̬�������/�'2L���5���4�BEG�[.0j�kT��>iإ�%B6�����9���������4���|� �@	��<�C����l�gS)��!:��IP!F�qE{\��������~�ה9�1E��v�8[IA\�~q��Āѭ�1��?��s���G�9/i~��ە&@��ƴ�՝ꋭԼ=�2��V��>�a�R�ݤ�@:)�,DVvs��[^c��@Y�5M��"�ܻ�5��n���h�ޭ����͞�n�Sk���{W�K�[J�@�)�|��x��G�'|T�U}:���8�vL�b����{�z��IY���F��� :�\��Xeaz�t�L'R���݈�;7k����n264'DB�)�5�Ŷ��:�`�@q\7�v;���jY��s}_h�K��7E��u&��kmj3�X\�BU�ͰPg#�_PZ��݀;0��0)W�V�@���چ%|�Tm�k~}c�\�W����A+$V)\ґ[��ʖ�����u��	ՅC�Z�������Hu�gU- ��:%1�@��=8#����;s��0����|�W[��d.#�@�-���߂TXSUֿNa}2��K��0=0����_tvg�"����������}�m|ٟ,�~��z�?�շ�c��ps�;W��-��5��/�3aHf���꼾!4��XZ�(`�Q|s7�"p=�%�e�x�1�e���B��{sn�t���kj)�jg\Zo�B_��]��KױM��n>�ͳ/$�ψ���?��h$�	�  ���n��e���q�b�[k�uwh��>[D�IzϏA2�ߧqK�NO��P����D�0'���ڛ@�*��K�"�ٟJe��wM/�$�^��+3������Cs�h��pE�����Kk=�~m�	+w뗮D���:��#�a/�
X*6�PGZuE�K����������Tkgg�d������>���1�TV���M�W���K[������E�Ӝ���?���5�0�G6l�#�(H̼	�Zt[5�
(���q�4vX���	Ō�k C��_�SpqD,��e�yo7Q�/��F��ړ$�JT�����������˶B�,ʨ��L�X=� ����'TL�c�(ʿ��{k՛�VqZ��*��	9/S �~.J�{Y����>"�Թ�J�Dy?)�^ܮp�D4�<2H���f�8FtM,ӏP�w��� �e\d�] ��u��ݿ��)f��޼��0I�2��G��3bJ��;������"�X�����QT�$֬�F��� �.zi���J��e��q�N���%�� 4t���K�$K�~�R�kQ����n�Rjr��ө*3��b�v�0��feO�<�!U�r`����� �ƚ��>����~���� kR�r^H������j8��˒L�!��� �}w�rd���%��>�¡�]GQj�A�u��;i(��i���J}��p�6�����n�E:4�K�R�E(צ*p$�b^d�a�A����`n�9C��O~ ���>�.h�bB�Ҧ�t�Z���V��68��#[Yƚ�����9�9H�R�5���1PJ�Q(�>��cF�TӁら>H�!Z� ��&#5�BM�K6{zw|�O���}�5xw�]�$;�&���kJo L�@D�L� �����>����c7L�ߒ4�����Y�>�{O�l�5ր6Qk�`�y��k�8b/���	s�+���D�l��}��:_���zs��z-��״Ae��w���|�,X���֝:K���׃��T2(��a�,~8g }�G{��_jc���,��������s�Λ|%AC&x���0"��7?{a0�v��f��C/�[G���k�sK���
�3\k�g����T0��$8���a�":��M���pܡԌ��x��U`�J85�H��~�Ge�u���R�"��%�Ύ�d��.G'��4m({��%q�?ڊ�@�6�+���H��0Ę���²�᏾y��?fg��0�H���8s�).�yIL����ԟV��s�C�G�T_K*�^Y��%T�fkO/�i'��\E�R�HP��y���j������F������ډ���3v�0d�(�M�z�U	z#��!�g'��kj:�U��X�&�Ȩ8���́ᄾ9Gj��#�ٵ]���ig
~?vn'-e���N�O��4�0�>�@��4��6��������/��Oz����rp�'� �x<�?7H��(y�
�U�uEy]��=X��V��q_�NW�	��L���@&6Ǜ21RU}��4�Ŗ���5Z#k�wte��-Y�_V'c�R��-��PgZJ.xg"�i5�Ɏ�"b,��9Gf�/�V��&�V����(�����d�D��*�d�\�THL�k:�����.ޢ�LO
�KAN�Q2.~��;�O���~��P��ݶ��ۑ��]�����_�<ɯ���S~mT� 2R���P8�`��ܘ�]Ȗ�y�NU��l;$gQ+dm�$�зB�.
L�}FQۧ�1�q��h�bP�4�Yn;(hbM��3؆q�w�+�	�a̢B��ed�bU���j�����Fȇ1����G�����'�o���Az�L<��E�C��+�Yۂ�ivό\Iw�$PFt YJ�pWP�.�1~v��v[PI�ǌʪ�gh^�q/EW���r�XͿ�pp(�A�?��f��{�͠����[�Qv�3K�԰��%yi%S���������T[߹H�GAL�!Hm
l}�j9�2��Q4�a2���TB.�8Mko�)�;�s���P��e@���d���/�}z?^�h��$��#,����S���}�N�Ʒ�^A��	u�+��`�NAdI/�e-�p��O�Dp�6��e"h�t����2N�����>�X���$�J3���)��ڦPaa��C��)�����떆�
��Д��O� �A�Mٕ���֟�﯋�ײ�&�<8[9fÎ:�o�iZ���'E��M�4�P��PPش"D ���l�-��j���_x�I�4B�Q�DQ����ђy}q���b��t�D���ϐ#�%�e�`˺Νy���Cg����5���O�>��kz,4�b�ӝd��ļ���>�4���ejpl�<\��u�`���|ɀr���������E)�?��2��i��3Ւ��%������n�����dq�ԥO=�ؽ��S�Z��5���S�6:-���������������G$�Z��J�M)��P�����$��]��G�}�||�2
�V�2N�G��a�����IĪ�΋�Z2jՌ}��c�E���4����.��9h�W!E��e�zX���c��^MM>�µt�l��7l�SI�J�����=\��1g�y�{�r��P3��N��w
�\S~;%m������x~{ �%q���ϪQ����,O^���n�XS"��5&��q!0jJ�����)�Q����G�����L�J���b� 4ȣI3�|���+�t�M :�*|"�t_'$P�(����+72��6-��M}:,���!������1>R��K���aЛ�Q��1;-4���k��S[�'d��J�j�(�D��Dzq;@��:!�,�T��J����r%l'O���=�M�(��EW�/M���-kp��44��K�şe)�K�e.[�{�2a�#�u� F8��@��z&���y���6�d}�V��Ե>���n�nE�7[��Q���Ӊ�+ݓ�:N����r`��s�&<	�ᎋQ�<��ٵ�5>�R��q��p�U��3�ۏ;,�6�K�+��&��y�?eOfksqCm�u�HmS�q����d�ӻ�(�OةM��pl\)W�&o�d�E�4�g��<� ���;#`ƪ3ήoX�����#p)��	i��/|��繸�,�gƚu�����X����5	�i�}"E`�wOO=>�*| �^�oo�9�2�Q�0Gv��ôx`�@m���	�F�;�6����N�J����Es[�g���� �@-���I2��7�g=���=]��S�^�,�Π�ú���FA����H���\�_4�^h�{��=��R�¿x�c_��5Ќ��s�=�0�I�C��Պ4��_��;��ϫ킝��f��1-Y���`0e��nE)��V9w�i��%���E�����,-������;�%PX*#6�%�����2e�.��oB��j�����h�i�����3c��H�O�S�6VQ��ހ�_�*�ε���PP�e��xXRs��X#����/7�2�}��n'�p55�YŹ������Ԃ�������@1���u,��8�����,��vho�(=kʽ�/��y����8�q!������{Q��|�e2J
�a?	��+�jH�^J��{�3τX���=�лÓ���R�On[��1��ʡ�T����KU��z�v���ܓ<���H{oHd�ʞP�|��a��� �o��'�z13�Th�q�+ۣ����&�d>�u'��G�g �B��d�������]���^����CF�1�\����e� ����:��Hb�j�9�/�h�Y#�& x9�^_k �u�R�D$C��B
�{=�d�9��Z-M��Pp��
z0J�i)�п�QB���0�C��Gwye��
�dzL�ʄ�)����'r}���D��QRB
��~����խ���tM�?(�4���1�$'�P����c������ZL�B��:L�=R0)~׺r׶���Ke��ᛞd�8<r�R#�̭7��G��]Z� ��i�=��Y�� ��qB+;B߸aX(����cqρw/�e���;�*z���%]-+l�う���*w���y����`I
���DJ�^����ʁ����5\mdr�6f��gLL�#���KI�`(?,?b�q���>�oc%� �[�"cnI?��x�P{}ˈ�끢|[��M���YzEJ��rx����-ñ����Ư��g���{�*�2#�o���@�I�i�����p��V�=XM�ɪ��$�8iWV[�����Ѿ���� ������?����6�g�ڮ���w�sԖ>SrI��Ϟ��<{)r��mT��5�xN[���1�+�q}��nfd����ɛ�r���)�/�Ͻ�3e<"����kF�� ��˘g��%���WX	�����,�*����_?�l��=;ɵS���N��〙Ft&;� ��[V�g`tK�@��"�)p�W��t;��A�4M�I@��0#�$�TP��5����+@8o���|_���J���mxMM�� {�v`ˣ ���j�K�!�,1�(WI?ָ�ü�XJ�U�p���K�a�3�l�������/�6��h��:�G���R�'Щ�j<�	�-���tRχ�ҍhP�j���Ap8L��p����r���W���]|�<p��ƒj�)M�^mґ��� �	��""�3/>ƥm�Qv;IP�M�����~A���̱�O�7�s7�AK�ȝ���].�h�^pZ}�6�����ͽ�o�/sMYg=Q1��rdR�hy��d,T��0>Ճ��^�t�$�Z�F��$�Q��|���5l�%�MP��bkC��̫=�KՀ�_BY�#����sdJ�@�~B=�i�����ee�
�L��w���$?n�
.$���+2P T	\�)��SA��e��^�jZ����q���"�ܿ���s[f�И�q��)�k���\z�B'�.�0���Z6r}�Ǐ�i��Q�;�:Y	���O��������T^����;�m�Q�x�����4}V"N�q��h�aKum�����^����T�� �0�'�+Ie}z�������L�p�d\���~�%��|=��mWS(�����$O2�Y�m(�ZLW?`���{��M����N�նWH+�`:� T�˻�/���d�O��p�>=�/k����1�h{>p�V{	�״q��c��E���ֹ�&�g�QcC�T}�/Y :c�Aj��w>0kv �1l	,�/��0��s�~vZ�ʀ��8�8�~��1���k�
�2w�_�8���O�֝������li�T�.�n3��p�ƚ�s4F���|.��v� �0l�!Rr���GU{ �Z5[����wtR�f��M.`�jY���%��z���܌�B�E�m!t4�ND���M$�@���v�V��jn��wi�l�6��(<6����7�,W��A��j�霛����q���n������=9
]�G�fᲪZxR*��O� hq�QLqˋj�������w6*2	�J
Yr�*�jn~��U�h�oWZ{=�TA��pR��X�דsC��Y�l�^���	��=��g�$��/g��",kG�]�\X7�=���	W)�I#!=u��W��ϤHh-�i����N�*�Γ�ڢy�cΟ��q�����<y
Ҏ��@_C�ow�����Y��]�b�|�(���	��2&B	�������B��	��ņ�h��$���0�:���v��ҧ���>�3ʝ��=F��@�l'��ECO�e�;�Bv��F����p�M��/�~�%W;I�]�뢷���ԝ�قp���
���b��k(�Ȧ d�A�3�ى�G� 0��0�-!��zŠ'*��-dH����w��W�u�@�Ȋ�R����YM�j)BkI^,E����$�]z��ʠ�ܖ%��A��E�p�fe�P��W��a����{����y�`8J�S���-�3�իܢ(���֝?����8�/�0�694�`��e�Ż��y5�p�F�qajhlxC��-Ѝ�7쵝�x���cҿn�d�������4Bj۟�j}�q3F�Q4$�6E`"!I�i��w!؍���_�'�K��=�SV�͹�Ƣ�e�c�X2�{Sd�fȩ������o�4r%o�:��#���,���K��B�o~������)uJ��.��*� M�($x����s�����0�mf�QÍVi�3�ٮ�Q��7�iV� 9�N�[�(����f1D
����9�Z8�2#��)����0�uf���?M`�l��^��g�_�@��,�,�]$üْ���XQ
��3^���ǎ&%��ó�0��u���$8�Yg٫t��t�i��F�n4�m��tN���a���j���fW��،��ctA��P�;�OxM`]]���M?e������(S��4�@R���ko]퀞��ё��ς���|�+�� �=�,tl�
��&T�������Άg$��وd��:�Ym<)<�0$��m�V����y�v/q<K|�HB�|��3>�UvOM_4�Ԓ�9o��4�|���`��[��hzU���;\(p�.B��p���7��A����!d%_�G�*��AZ�`�,�4�.E�3,��yذ�u
��ɉ'@��D��%ԄYz���7՝�=x�y�Ҷ�*��c& �9���!��dM��4���k�P�E>l��RE���K#=~����HOJ�F����6.`���ᕞ��gl��ɳ��VM&b6����#��tU�[����͔7<L���'D\�m�,��xBY�y�	fwT˔'ͤ�"�P>��t��:�����D-��;�������	�D5d/佛0=��|���/�9�l�H׾����lƣ�eM����IƖd�,�[ԫғB $12�ue���:"����%�����F`�4���.�	(����2FZ����!��'>�E�I���_�5v6���.Tg7¬\�٤t�P:H+ !��m�B|�݄��<?�l�g�>��QFo.�E����D���o�,�[eJ:>ʭߟH�k5����g8wn���[�6���S�,��]�v��l���s����L|y"%=F�&���p"�,�R��o�=iʡ�\��
~7Y`$԰K|m�����f;�$D5��9�:��Sl���a��� �/7���B��Tt��g.�>�pt*�[tc���C����U��6%*�7H���z��!��0 ,���ȷ�`���6D�6 e���p��$�}���A��.���&Q �ރQ�����Q���U@o�y�;��PCې�p����')�k��@�S�y��Z?`��*!Z^%��a�"�<�������,d�X�g&1h��������vZ9U���|+t�@a��g��<�m�-=kބM�m�,���k$���vx����N��d�h�r�ȇ^"!�d��m��6��n-���d" 
����G�A
�����c� �>�K�CK�7U@��!� ��K|�Kx3��v*l��:��exfaٕ��{��b�W2�sf��H�QJTx�tך[�0j�?ق
��E�@#Kpˮ�S6��-xvX���v$��0����6JL���1;�E���{��s�)�_�L��7�؞WD���ĵ���"����m�7��]��{ް:
B5.�i�M!c��rn:N�Ż�|}�I)��%7$��u~������[ ���6� �qj&B�VBW���� �&�K�9i݌C�6tŹ�О4>!�]N�&�4g��X;a�C!�D�$��K�)F� �[8cm�0��8+a�~z$��d�5�#L޻���F_�s��2Z�p"f^�����4��M1���u�Ӳ<�ӗ�GuS��vQ���?�s�#{Ͼ�}MD���{�U�q�R��#<�#�|��&�SHb�=�<�g��D_�	3�?���W;^c��5�&�ؚ�5?��'�39�?�U�i���O�͸������NI�V)QR�%j[0���2��KM�swWC�2��w*�c7cY@�N�?މ4�C,O
�X�ilz���9q������:�!�~��UW��٘^�Z�y}�`2/-��-�P�!j�"K</2~�z�$���C�����U�E��b�����@7���F�y�W��iKREp$iK�V��ي	")�!��9x*�3A�WPC���&Sm
�DW@O3��~�V��u�(�.�!��R& �9��/̌�Y.��w^�Wx<&��m����U��Ȗ�=G�������ڭ�v�"�i�aR��ҹ笏&�x���2�}�����(j��,\�m\R�7䌉��Z�9����ǹ ���kgؚǡYl\NA��l��Y%*o�9����7X麴���̙t;7���y��F��.
9H���B�I���y����,vs1۸d�k��]��H�yT-c�C8�2Jp_ ���T{d��arq��E��,�d�%�Ff�ͧ�g]!����s�� �U�]SCrvK��
"2�v:���ߢ�s�;�+�CZDb�M��zE��*z�9�]=Obm�}����p��q�W�t��/S���y����J����,`�l/�c�;��nL�a�����1���?.��=B�r�Ĕ�%�f���	W����~���o1�b�a�KYj�/�u��3�]$�)0lp��&�hBA��W��K�墟�a�\���4[t�1T'4�!8�0�'�P�"�Z�v����Ó4�%�T*|z2���%3(�qJ}W�2b��Ul{&$��+9����mW�!cOy��c��5�*b�,vzM��</͔#Qݻ���sҾ1h>	C�-t[K�������܋Eo��p���s��a������F^3zs"A��k 1&�/	� �Ug���e�&�����&��������D�To�S�V�T06՜��?����cK�Mr����7�cr�b��C58���2����с�WWr���{)6: }/���c�t��ah�	so|�:��3��_*=S�-���,e��Q,o��W�ۜ�5lsB �f�u�V��n&�	v搪w����*2OϷ��Λ   �d��?���������~<�6��˃a/ �v5c��бXeҘD��0��k��a�����?��%v
�Z��<W�F�#j�E��8Lt��^�[|���Z��!� ����>:/�Թ���\�����M���%;���Qq��	}�;P;�#�Č7��}����y���������>:��|wr��_����=�Q�"��@;ÃLk���Ks���Yr,`W���s�`~��a߃�;I qk28|������y�F(g�ā�kA�|Qni�.�w�����Xa*��ګ�/aJ�ꖒ�����I3�u���,> �z㘍+�~N!͍���� �t��$�����Z���í��8Ϣ��a�G��"a�ʢ�R�:\h	Ҭ����dmʑ�a���܈!�e���J��hD�|�p��U,X����kQ���68\pV��$�K�>��V78�>�~���Q�9ϥ�}��z�H��'��oD2�A��H��!Fg�i�ݬ�l¬�����ìE�L�նࠫ�C1~�8rHS)�3����~��[��N� �)�\�o���"w�넛up G��N*�9�]�<��gMn]����x͵�|�=�z��3�`�g��������H��9Dک����T�&]��ۦM��a�T���L���}'���&E�?��Ǩ��}�Q��,�y���X#�f�-KT�oQw�Wr?��i6���z��������a��oJ��>����Af�ˢ.�hkrY&~j��*���K+n_��W����r?W2K_�-��p�'��z]�Q{[}˫��U�	�p��d2��&z�Ga�h�:��Eo2�b�Gݫ�ՙqJ�#g{�e�sְ'�K	4���`��u�E9�W�1��Y��3�˘? �Ó<[���ߜ�F7e?��k��y��������6�b�!=��d�p�.�W�,`�=�����<�t����˯P�w=V���.w��|��uz���c]�V����gU�
js�r��f� ����������j^��IFHj�o6��Q���1��6�GV`[B^|��X2�3��z�_4�b7�fۣS���g#U��F���Qw.�S�EŖ������=b��v(��?�����g�Oʟ�nٞ+FhO�E�!2�o�kgn���e$��7��0�7�$����F͊�l���핑ЇO8\����Fz;�L��Q��/�2E9qi 	��+���^�d���ze׶?�@��-�U��"��!���0��!7D�:���a�y��KD�7n�vY�[~4N���v���4.3��LSi�.IO�����x�sR�א���������3ow���6!(�@
�j���::���~P�+�71�\Oƺ1�k�p1`�=[�|Ƅm��J���+fZ�L.�o�w+�@����Z�Ac���/����0d��~99�6^�u�k�ٺ�܏ � ��0�����]�;Y���!�=;�������W�d��O�W�n��r����d��6�щ��wF�¼L��	c$L�t}��*gxl�<ac�C�)Nd&���#�7mDpAཧ��ʔ��s��2�u�s����T�zQ��ɰL��fC�k�S�;N=�6�یXc���9���G��OQ`�X�~��ÍQ���_J�4��2,��_���R���K�����fNV����+�*��C���vq�S����Z+�i��#������0�Ww&A�M����*�o�q�"��Y?=�=����+�+[���o�J�6��-�;f��o��ŽIU=�s��P�����.�KY��G�C��!�cO���P��P��m p��v!ݢ�1��a y�ua �=&`gd��#��J�Ԭ׋��](x����BƳ��~�����R���5��|Z��7��h����,,e�3{V�����:j<�9��b,$��@�N��kC��l�Xb�A�G'���I��w'��	~�VUA�m�yQT����1��j��<��CP��qY��.�fx��=�,ꇍ	�F926EU��ؘ+q�������H?׃S�8��,�;>����'�9����c2�'��0ήa�ӃR7̱VW��k�~�KC�RBt�5y1+����v�g�&�x>t���:�љ��R����`��!� "�Xo�E���8*hL$w>�%?t��!\;���1��r�OKu����g>P�	I�O���JtZƿ�]b"���S}���>F{��@-�1y�d9;o�_�NV����c���zY�����?����)q����&3�C/�b%�׫D�'�?�R��)���%�P*9�@��d2%��I�<�i=r�oKNԑ>ж��"��
ϳӯ�K=x�@v_�,�"���w���P�N�g�o �PAQ��VQ�*�(����|1@�J�'��+�%�N���+N�ގ��Z���"��D%,w���jI���@|�n�ʊ�`�x�y�1�����RK=	i0-Q�O���2%i���n�h�U��V�uB��Y]�}� ��u�ʔ@f���4����m��+*JM�m��}_³#�|�t�	��i@<���͑%N�·���D�rc����eQ��D�u��gL!nxn�ʹp��)f��-׏��2�]���C�x�ׂ(��e6U~
R��1�'z�*u%f�|J!���q,"�+��C�*wH�]s!6��9�5�m��������W����68J���U�}��a�p����ݤېd5��D��G�]�t�xO*7lfၗ]d�t��u�3�Aqm�O0҆�Fhz)0�;��HGG����
�B'v4U��{��A>�/�w����j�羁��J��x ��2�<���}�mω{�@����ѣ�>����sE�����V���K��Jdo���ON�Db"U��J��n�q(0�7ͼ9�w�r��8A�[�S�[h7�7	�a��2SD�Ʌ��pR���2�n;6�|����:L���E6�f��K����;�v�<�0=�Y/X��r�a�"C�t�z(����'>�L���t2o�w�ݻƥXL���4�X�+�O���ud[L�)$�E�F*P�jϤ��
�<��� �i/ÁR��ij���Y
`r%�'���e:-8����7}����c�5TT�Zآ�Dk����9��G�TЂD!$:î�k�qz�ť�C;f�(o��T��vށWR�>E�t�s�w�C NC���Oq���J혷��K;�G��,豼��s*�_L`�Oǣ�� �ؘ�`��Zi ���̗�����A����]/Cw����P�V03"�������U+SΕ�&g��:Et'�`�1�pQ�ԍ5�ijn~)�m�Dr��&�'����`nf�!���icd%ra�eq�T���ᖻ��iV�zz�"��N\TSA�\eQ	��G�p�:���zQ��3����a��T�� ���y�fSl�D=�8Z�d����ߡ�`])� �=L~��ONg%��N���<�E���(.�c_ʷ^��ǓO��H��$E6������, lХ��FYc�dR[u|�sl�P��5bŹ�=/�'J-S	l�}�2_J^�ԯN�!_R������������:jG�8�]"�W��/-�ݠP"�M�m���#��a�ѐbSk�1D�F �7��,����q������ru�]M�, b�zN5~� "���\s�_�b�aKF�q���]^>�аa8e�G~,�o&I��w;�>�)>zӂ���cK�T2/�j|6����uU�I�@m�=�k3&3�_��z�8�ힵě��ŀQ���T2�w�M�I���U\0�f��G#�L�6W\�zo�,����1���2JYV)�0�l����Z�_f�=/*���+ߦ��Q���ƦcT@އ��r8ȄK�GA�T���]"0>�d�4���P�d������aq|S���*�UM�N�=ݥB�.�ގs��T_�wB���������q�%�7Фֽcz��5��J�/2B���ZI����`�@��px�|�C������,�١�eF��đ*��q�t�ԈǷ�f�d��q˪�Z����6�(R΄Ү6�|_���j�q(��Th���d �2Z�\���#*#Hh�ě�쮖�#Q P��u�Z�q]�3YEN�W�$��H�ճ��{}<ݞ�]S&Y�Jۗ�X���h��N8Ʈ��(����~��-���|_{��#?T�i�]I���.T*�Ǔ���HC$� i�`LB゠m�o�ȼ�V��l�h!�)��`�ՙ'����4�L`��Ru��_��P<��ʟ�[J��^&�ޯ{��hNZ�f��)��ǘK�>9���s40=�m۔p<٢�]̜���E�=��O��Z�v���n��B#2v w7��8]�M����/��^Ng�?���8Q�`���^E���2-M{����T:!�Nf�Dɭn�@P��RZ� ���/E3���5\�dW���h� �3�+g����`���.����M�C<����qŎx_I����9&5Ve�Bk$�#Sx.Wd�;��"�'�Hn�4[���˘���KR`Mu
pE_����p{}I��g�	qѥ[e�Z���Ft�\Z�_�H�\)+�Vq�:S&,�>ӨJ5B�5������!O�|��wV�=��
t��u(��Ø�"�&��tegA��Ɔ|獵o#�7b���n"j1hU6���g{H��I�8g�\̭���SU�"���~�ׅ`�d�5��/u`�}X�H���"�2�
�^��E��@֍D+�;0+U�3\��~��i3}���u{ޕ	�yFI�|���-��(��[3�9�z��$ﳐi���g�+.�.�">��������S� u9M��<]R� HX x�6��m�~���)��X���nTQD�.��+`{��_ ~Ԧ��+�J�V��6���G�g��,hߺ� �FQ�M�4QzΖ��7 )�pg��������M5{���k^��=M�S�މ�S�ЂƫM��ζk�`rt~ ��%�q�̴]���%�O=��'�� �튒/�{ӫҶR�,"�-��~��躎@�N6��,��\��u�B+��27 ��,�TX�䄢 �C��I���~�%�i6��U������2���%�]]:�S!^�$�0-���j��`u���A�o�о��)s�Oj�Vѿy�6������q�<�B*�����)t ��w�H4p���^�"��Ƹe�Eka�r܃�@� �lk�SOJ� hAz�!0�U�0�eb������������$�%��<ۨ��4�cR�7C ����tx��u�mCB��4����e˰���?��xz�wØ_hg���{.+뷭����\c;��҇�- 
z[7dT�~�6����/�i��P���~�%ڤYE9	�KH�]��,�3�t�K;yi���'��5��nࠦ�G4�{�u��;�Sy�"�U����]�~B����q��~��>su�������!����5�V�����: .�ka �d�%���5�*32�}Vִ7�[���>)�;��)�1M�S����8)��1e���Ӗ<ܩw1<[�^���8F�	������n ��6��E�����IM��&X���调<5hR i�=�OKϼ�X�m�,������#�&�4�-��ۓ���u���=!'y]����*����c�ä-�[�l���^���?Q��m^���1�ss�z���<G��ɯm�|��T�&�(��4�zh�Z��6a��� ��$}�
�&�}�&�׏/��,��/�:!v��&��:�`�;h_�c�;7h�z枾�N��h�G��s�F쌚��4���,�6z���Fb8�_�U�����f�;3z�kUF�5;�dW$���N�<MҖ�9���Kl���x������ױ��o�����x��U
u�w�wC�4!��5�w�ΩA���O���l[V�*�"�#_<w�M�܌Oi�,դI��~S��6R�W�㫑�Д��HcCa�[Q$��d�	|�v&B5 3 ��a��\(;~>�1�N���Kö$ǋ�6*�&u\�{gm���Y�Gؒ�A�8@R��L>��!���Y�|`٢�Q�Uߴ@n��y���S�!�{�[6��i�d����I�AY.էe�������Ƒ��BEޢ:��:�rL��;[тt��"��82k�znfP�Ӷ��\~��<���m쨩ƾRnX��WA�w˔��(�{@(@\��\��ٮ�g.�O�	�7x��Ρi��Ocοe�LW��k��|a(�u���xn�� ��ħ@����w(%��u�[[��ߐ�,/�G�v[���@P���[GD`z*��ݫ����\�o0�nWk�� ���o�ay���rV7B᎒��(�p�1&JWK�`��C$rN�j~wEy�kp�����\�Q]���f֛;io��=�&[�A�^Q6bAD��Y=)��&7����}^ k`��śy��x�d�K�z�A�!ƈ12Ơ�c�Cg�mz�|"5޶���2� N�/E���R8��ݛ���1 %�٣���J$�����Jg�Tt��ئON�懈��N����Ŋ���׿����u����4̩R������4̟��i�- c��h����g�Z��"�u�{���h�@�FtUmze�Y�ْf���u1��>@hة��>���������m���vC�0\�r��,�دܽ��DM�ڳԱg[�3Y��q�&W\+G���Q}�0+���棟�ha9�۟��:���Gu��U*���L���Nע)��X��,�ü��I"˴ª� f�+�ky��l�Xh�w�	E���3�� ���>h�t^^@,-$���,������- ��#�(ku�m^c����F�$�V�v�
݁��6�j��Ǳo�̐wU�my-�f��=�[��\�/ݚrX86gw^�4� �9�15J���!�f�(q�,�	�Mm��l9������7ݕ;�u%[���Z9v���e1o6}��y`��?B/�ʷq�I�m �_��xu5�*4�`mO��������~��I�,h�F�G��|V<�,�6o�9-j����v*��h@�Vv�M�y��a8�f�2><��;�.��ԇ�0ә"S�}�i*]P���Z����N0_�5�0$E�/T� Z�~�����nN5����5�٩�r�_�<
�V�}68Q��h�t�a�v�I3��v]�'�����[o6ch�tNɃ%R��٢������N�4�X�7ԌTK�����%뗐= |j�i�'�
����"o��P��xr9O*�d���T��2��e��]H�x�v_�p����f􁌴�w13��8�����ʑ.[�ξ�����Gu	� =
�G�,�T��\��r�oP����X5iy�(�d>6+u*�H���#��I�F8�6��J!�>�z���S+�B����02?�SP�i��CIۙ����z�kk�F'n���D�O6;Iь�6��x�,R��?�EP� Y�Ad=�U�?X'{P�5�#HV3n��}B��A�[)hs�N��ܞ�[b@#�̽I8�ץ�nXuSӍ��O���2�������7�ݫQ�7��x�/?7Yt ��g�}�HP��,�N6�zM|�X�3�TCdd�n��*K�ZǱ�r�r���2�C5�叕K�kQ�ͭ"U��zJD�i�ٳ�͢��%(`=��Ңw���Gg�4�ȟ�HWq����a�vE�X�8���؈i���3���1it�$Rl~C�X��T�������F���y�2Bu��dم5�%ـ P�?�,�;O��J$~����l�*�ϻ:����!�Ly-�%�ʛR�鏠>!@rΆ}���T���D4W�b�@Yْܼ�T��'�t=
�'�8=hHuk��E�����T������=E�X�>�ǡ�;f�@���ZO��U�
�&�>�����rH�.���N�/��Cq/��,}�EO��#�Ø7���$�U�8��e[(��,?��1��M�� �;[�}���B�]�6�1�e͑ű�Pέ��7�*L���^��|RˉFbq_[;3o���
4V��D`AF�ЅZ*R�z��(R����ꜥ���qJe��/Y��Lr��䄐�_�_�	@]jaq-X��T�9_��^k�%%����lR>\�|�yw��['�?d��G���T�V)c���8�0F�]���5,p��/]_[�Ov�F�C,%�8T�:����� A�W����������*ҋr����u�('��ѫ1N�H��/}���B	�������2�|�.�����݃�5ϯ�Zu�fD�lO���}��ۖ�ru5)�g�R��Q�.K1��9p����y=u �wx���<�#@��1
�4Rx��W�_���������,�|&��\*F�=w��=m���M��m�����#�L�(MTFŉ��A�$��k:7���L��Qs4��J{�l���(�~�n�>6B�s�4�Y�������L=�Y��Vl�jcP��Fe"�؏��.�����1 '�8��;�y�Vv���W2m�ⳙ��ߴaG�}B��;��զ}!z�P� ;�[[�5hr����}�|c���Z�Qa˔V�r��qO���X��Hs��K��&R�	���:C���r�c���sM!���g�B�a�6\M+�R!��Bs���n��	3_xמ�±���9�څlV a���~�ӡ�Й	�j.����'iL�D�����!(�F7.�g?+��g[�X�q��ݹw�q	jCHJ�5v�v�����#���T��eȳ��o!^gJ���z�Z��2F��)~���u�VTd(��2� 5M��d6��&t�[]"i�}J�,�l�F��P$nJЂ[���<�CSq�2��S��j��Eg�����6�������]O��.���u�F�[B�O1Ȃ~��S:ԇ�IJ��US��)���~a���������q[�S�����?����S2��I�ɛ�� 1�t�#�� ��}'@D�?�[Gi^i|���+����\N�q�L|SN��D��7�R/7�����0�e�������'v�'Z����g�0�.�Ye�4E��,�=�i�$�mV�q�׶�O�MiS�q��.�ӣM|�C�N}�F?a�$�҂�CVq����|~���h���[�8�h�@�&�9<U�ܘ@���� �h�Tԧ��U��qB�W�T��p�=aT׉�+0�y��Y��F�|�w���$���V�-�����
~,d�=/7�}�\�s�ǝV:���?�} w�IA�{������ʺ�w��A�b�+��$GV�j,���~��fs�4!t3�[�fN��8�  ������z�s��$7~�2s#=`HJ�O��K�!�Yju7誮�Wf�q��w)�a�+!���OҀ$��<������s)�hf0f-.��[x��9+�����Uwp�K�䌢8��}ՏHF׋"�<}�6��.FJ�$��9��9b$oVgb�<V%EX��)�sL�\�p���T!sL"�VŤNpp�0ԑ���u��%���Z]C�l��m�r��!��x�\+�Z�������tq�d�9�|�G�E-<�x��x���,��6RJ|-LR�{��!>O&m},Qu���Fj`m�����f�g�q�5��.��'O�&�K̘N�͕W�ˑ�,<�`
`ӉhQ��֋�W��6�w�s0�RQ2"Y��%ʫ}<�����I�y�>O���*Bs,�k��I]IԎ�%~r}�V3�i�6��	�'�~����-�@�#~��z��rz�3��lg�B(��Tb>��<�:N(�`6.�f��Ǡp���	� uEI-�[�pݖ=l�L3�1��9s�	t��!6�O5�a�E��F)�!ڒ-�o�8r�S.#TV%t�M�� )_����M\��V'�� ߽���ǔ�1��t��Vu�����I�S˥4�w�1�i�h8��Z��}�?���Ў3�%+�s��/�]�"6��:�K+����9S���i�������&�j��]l�ʶ�3cy�[����f�V�Ȅ�a܋76r�%�����T���U{پP�:���X�������?��)��2�w�*�'��q+B	?�:]ԃK�3V��1(R�dY��Z�L-�D깁�^�j�/���e�]8��D?�}��� ��DKJ�����Y�Pr�}s?a�ґ�%���!!��cJB�ɶ^(�&��� O`- �'����E��� ���>���Xi�����ObTU��XgZ/+C�*��#棢$�?�6�T�T�7���3W���RE�n�Z�UC��Zu�#4�~0_�P�:Q��	��#�mݨ����kX ��~��2�`D#�'�
>,��;�A�0�� �пf�[�&�REv��h�Ĺ�^r�]�ܾk��؜=��	Y3\����3�L"�E0΁B�w��*JqҔ�Mv���{�{]e��Lp��� `(2\�E��@)W)'���� �`��g�I󵃄��m�ВI<��@**���:��q��\��>�UZ�L�N5JE�oWb6)�d�K��E%��R.���%V�猴�����X�'@�n�v�q�c�W�*-h�!f�#�"��6ڸK������y>��g�\c���+�R�1Y��4b�����p �P��ݿ�Sy�����R;ql.*�LbX4?bQ�?�_�d/>1��J¨�X�5���	�X�ciTHI�2�Ƶ{�E2Mz�^8��b��P�������x��	����"7D���A�A ۴L��ƫ�Y�$D#������@*.z���#}�����(&�sy�T�H�UQ�I)�8�m'E#�/�@�$M|oN�GQ�XB0��iI���(ԛ6�{����#�7�IJx��������=n��v�;�#=�[[#$��:f��yJ���D�hVc����"n��H%������ )%d�kv�̷�K�}�6�L�$��Ip?�a�G8hN(���������آ�ï �����_�e��&�\8�u,m]Hc�@�ZUS���S/���B��0��cګviFgSN�9�)�\]��Ÿ �!X"��U'�:�[j��B��� ߱���~jU3�A�4�~��Y��e��@@U45`E�C��+����ܒ8��Mhrpg�5��Mh�m0�qU���~m�\ޜ���K{\����E꘡��ECn]r���< À�9kyĈW�L�A� ������+Ȉ3Ǣ�~x��O�nu��;�RȄ:	Kq�P-S�+5�5lt �����'��h*�;A���ˊ��O�D$RI���_��I��'��ǩK[,���솣h�]=X��h����x���]"a2i�][��[���� ?$�syf�9b����ĬO�щ�(���-&���Z��"���;x��������%�-�]\e`(� ׺�Uh�)YE��SA=7K7�b?5-���c/[{�8�q�rBo�	�Y��2�Z��hҤ����������Y�X+'�(�gd?���zQ�	����X`OS|/�35f�|%�`�}�r�.�g�m-��a�g�-��R1��N�8�G4給$�VO����K3"T*��䌪�N���ݞLX��Oِ�It���.�2�J�pm
�����ʥ>�q}q��!��=f}V�b����[�B�*��p��N���jiv������NA�=�0�=�ؓ�F']1��Ԏ?
��^?P�$�p���%ۈ裗c��JT�Ԕ�Ⳅ���Ќ�QGMd�sn�q^�5 
R�g�m�^��3���EF����T�+{/�Щ8̪�+ȕ��~^����H��z�a��	CY��E.dj��::�:�=zu��f����i檇�sj���>�q8�+�٫�/��ݮ��mג��� Y[�ğ�!�U�Ln�D��&P7�$�)��z?���k�N���߫1$��sM�lV�f��V�����
o t���+Yޚ�E1,&�a�i����0!���S^+jMI��w�V��e3�?o�=�)�u�Ԇ㈽/-%��������t���]s��GV¦q.�/�ur�$��{7��7#}z� ��:*�KL4Q��K0��RW-��R=�iY�b����(Q��!��E�-��ڡ�� ,/������'[[#��0%3�y�sI2ykМ����_2�U��	�З��.��泽����p!�؃� ���|G�}+�L��kV�;D:�H�밂Y��"!���Ҕ}f���&?+�JF�Q��N�Y��,D0�$֕5�)[�+�*��b�ɑ�g�as||�
a8N Vnϴ[V���R�xi������y<]⿢�{�F	OwPܷ N�z��([�ڤ�a�^��{�0�P#G��A9I�s��b+��~�y�\�gxX��^g�^M�����bx�r�*� OVi�#%6�@r�������P(z��ɲ:�޸LBC[�I��&���z\q��g)��	����n����[��:eS0G��9֓�ñg������K��1!��},����Z�u�����<�� �����?D.�y�q��v_�s��@�h_�HoA�Qi��_:9+�W�I�(�y���X?S|P}�/��.]����Cbs&zn��.w�OՐ4�͟P;��6�uz�p&,Xч��{Rg�;�s�������l�6-���d�����NY8�4?���r������h�~16ؔ�vD�g�VU���j��Q�١m�i:.���UA�N���K|,�&�47}z��9����:�T$-�6�^�������5�8����T�RsRA����TI-�G.P�;[_M#���]�D�[='�q�>f�6P��F!z��sJ;�m�����d�ҡ'fG��q�4C�]_W�1������:F�P,Q�I��O {N歿\-a�4������D�́On�7pk`.�Jm������$h��W�ǰ▪���Pqf2�+�/Z��Sv��	Q�:J��#29�ۋ?�Ui��u���������<M�־i<���%k}yCG�,�A
�7
��"tҲ�������Η.����n�p�ECn©5t�Ǘ�5����3�h�3�hꀥBR(��ٲ�ئ�%w4v`Q�h���вԥ��&��H���BY�@�0��Z�(�Hi�->���؎ ԫ^f�9��K�_΋8ƭ��"�N N{QUѳC|ݷA	���S���pG�1���E�8Ò�!#Ny�u�� ��Ⱦz0�1���0��p'b�#�ޝ�2�����,-��2�m(�@L����Z ��ɋ冔�uM���6���]����_�������2M[�?��b�p׭%�~���Mn�����i�=�D~Ӫ�Z��� 0����,5� m��N8}/
CL�4[�����U�17?,4jY�ҰI�m>���Mۢ����:��Ŵ����HC'�,�dw�g�(}��xBj����Tc��7��P'��J��Z���x�!���1����՝��mI)�ORt��k�7�R..�UbvQJ.��r���D׏u݃��\�s����i��!�A����np�)9� �b��l?(�1�3X�.�x9:�eְ.��2��w&���l[`�$J��a}8��*)��=0�ZXIj]d�k��i�~�䲷)%aC@V�yP�2�iD�[��԰u��0r��F]ɵ������s`�g�)�����j\�p�������6�njFwv�C��� 2EG�R�;���9(pZek2��;�h��J�ͷ���v1����ɻ��ρ��著�����g�h��ے�O������S�?@ߑ�Kº���~�6{$ ���۵!�F�7����8�W3����!+ۄ��*�YH�|
8�����!�����\�P�'��H������iix4Q�EPL������NB��w`zL3�`]�T3g�/�յ����~��6<��w���Zޡ2	��8A�3!�\V��|�Ibֆ��p�G�ӫ���a������^tO#�����3�?���2/������	���U�N���Oa����C���Ҁf��9Ih�-̨��!��OR������d2� ��o�C'غ�6���
��y�_��ha��o4PS���4
׈��Q[�8V,-=M��>��q����{D���~@,n\�'��~�zp���7�RjHsҲ�^�)A�c:/	5�d�n�=A�ygV��d:)e���q��G-9��T��Տ1���
��{8�˙�s������#�|@/(;��_4� x;UB��cQ|�� i�<��a��R�\n��"�A�)`wH���bv=m�a����R=�L�3^��=����W?]�#~����nqSu��ߝ�xPB�|���hhKZJ祳����hß�	�\QQ��h8X+�͜%0������>�Ǧ \�>�xowZ��	�R�-|̹��^�9��j�Y�Hħ��Du�B�[+T7���{�/|n[��+Q��J��Rv�Z;�/!%�*AF�2����{x���Vy��c��B�h_%�#�:^8�(?V.����;�#'׹�y�#.���ä�B�lwO��sZ�'g|&A˯,qE D;{k䝌"�}�2&��9��U.��.��r_�bf�Υ�N�p��4tdY/yH�;�V�,�^���"�Ȅ�o�]jYNWŕln`m)4�����%�ViM���p��耋b�ƒs�{��y[��/��,E�w���q��LQ�.�pb༊�f��&\Q�tD�����m�&343ɿS�� Zc���~�����>���n,�in��>��3M���S<B	:sƺ�1H+��fD��ˉ"�D?0WY�3�&�W�@}�����C.{���m7�K������So�L%J+�5��Lf�P��3^�t��cܸV=�ˣ�T�l��A��uz�� a/�v5hz�"�����K���?�z��Ep�ձ�n@h@΂s�a7�1��+��ox�f����)�;�	u�s������,F��>i�՟�h������l�]�9�To�_S�B;�R*��κ�T��m�I�o(׶%�ہ�VN����y��Ò^�Y�i@�#`�5_l��db/����M���=��F����%�K7F�i��m �B���/�����Q�MKX�ǀRK:�֮��H�}x�����(ܭ.I)9�Y}u���$K�}��e&���MȘ��~�|�Wy�Oj��z�W&��P���^/�7'B?�ċ�gbߵ�,��Ne%6��O��Uo����d8�%�m���:DՋ (�0�*ɓ���������%x�1
6��S�+z�B�a����:�"�QtE{�?�@���ǔL��Nv��T�%�v�iV����F�����mr
b,�>���˹�|���	o��N]p�B�7H��G��I'$��t�H�2���n*�&G��ӡ`u� AE�ly���HȊ�w,%! I�����~�Z�������A�0�3�]Zy^���X'�RuX*�.���p��<8\Fs���$�y%��H�ry�m?U�g����vx_L�{.�XB�úP��
9�D��QF��C��!���sI+�A�!�[\Ӻ+=E<�sR������k��p�*l�i�#�&���t���b�U8)��G��h/�	4��_�[$m~��xxD���I�ZJ�X�yh��D��.��'O�Չd8�=D)ql̯ ʉ~��J�g�iN�h�w��]Bʲ�"�R.��$h���%;�]��6�M6~A������rf����/�=��Fr�YH�I��'���>ʆ*ı��M&��\����KUí�e�I�	�1�
rg��U[���yU�nS/U�4�?�$�Nf�fk�!� egM+ �wږ��̿\ n(M��1�ɲ'lqF��W`����\�ȴ�_^G���HP������#s�BR��UԾ7s1q�~��Y
D��NF-�aꯋT=��eG땽t�ڽ�x�q���$�ױ�wF�MH�D�K��g�Z�����{�	O����DI�+qCuQȍ� g�,L��Lu�o��s(���E��
1�n�g����w�B�i���m���+�E����+�A�԰0	�B���i�$׽���Nk�y����Q�-zǧqFG�#�`q�M{��:|BJw #K��
A��"RO=*�_�H�bO�t������;�X;�a4R2��Gu���V��㴹N�lt�k�7���y^	�٥�#!y�kW\Z�A���ڋ�hˑM
+��9}}$]64I"c)�3ǉ��5�"v\��YhXWF?Ḫ�5��;%�����:��c�I�4��1��Y ����Q4�W���/�;<�]b����!H�tM�r�l��j��э-;�'�<� ���Ob�YTz�)!0���UK�rG��gf4۵:l�&�c�7�zIR�@z��gg>��
�\���D@Y�;º�]��i?PH�l���#k+�X�o*����,������!�-��آQ9#�N�"dZ���yIb��d)�{���D��e�,8
p�<�?�dX�����o,��ryZ�(��_*�������C*�l�,Q-�Z�*� ���z�Nl�ŊC�"nkR��J��*���P2Ihi�ə�G��A�{��kwoF拫ɢ�7=�n�>�8�m��ȿ���8}J����&Z�����rH}��op�N;��a�GtKl�(�ƉM��+�M����er	�eu=/l`*��j�7/�c~q1��1X=��t���.z^��U{8�R���l��	����� w�'(QG���viF����ZD���Cr>�۷߽̓1�D��=�T6���c"��zU"��q��^�Upۥ������Bt:��3N�}V�@qL�-�d^�`f�^c�^�YԱ0� �� �С.�}܁��e�ȆG�����\o6|��������s�$h��l$�+��2*�A�dqy���b�f��k<'ܣ~�_z�9��"ED�!�S��Ip��kK0���џ�i�[��(
W�yt�*�{.r�[�Ƽ�`��b<)D���������]�M�'��ǭ���8���9E6�霏��X�c��M��w|��K��{)�Bb�~|8Q6S@<�sX������j=>C���6m����Q)*�|�'R��鶍�{Ll�B�˱7��Ȯg@�(E4��M^V�`����l'��?(d�]>)�'���>E�0)���*7�''�Y����嫤c�'�&�ݲzF >�0-��:�z������o��jN�3�6;������?̲[��^���ǹ��H)i�Ed�M�wwS��� CպwT|���[�YT�!�J��.�X�@�z\x�	�����u@ 7U��!�vԒE*1�K��C�gX ���^�偃ab����D�%�����}�2�U��S�[�F@:?����n�?"��lx��5hyu(�v7Κl҉����WѸ��8���N��P�H^Y�U8*+?��B�S��)ͤ��3�}M��`9���]q�
���b�����E���4��l#BL�{	C���Ij�J�sd|�J&�r��/m�U���]�<���5HW�TҴ���L����J����\��!MFA�<i�n��̵�8�<��}}CͶp��62���T��Z�6�JM��%��~!�H��3-����=A+�3h7̓�4����t�d�j�5O56ĈI�%~�9��oS*�l�2oO�u׳�����M��}��U�mtb�Y���_����Q��}'���q%b�/_ok
�>�q��R˒L�&04��Z�6�q[?���hd���c=*$W\,SI�y�l��7)ɪ��J���&@X�
��@�.P#(��}K���lUYQIO�&�"rJj�(6�\��'�(��D�����e@<���!��䒆|������vLX��gFOEX��@Y��??bQF3�#֤\-�9�ϔ�%�k�?!/��3κ?��
3�ۑ��X�>类�0
f��f�*����^�~��	cIa��ɧ�)�b�=5d��v�U��h�4���|�=�[X_`أ'l�Gr�=A����nD��I>�`��kr��g����?I���9*�έ'.�X��;�����я�*'�D���g?���cd�2���WЙ�;�(��sOF+��iAP��:㬱1���
���˔� �\�e,>������{],L۞�{�jt�Y :��/��/��QZND�gޘ�Ў�&��u^��[)V�p�׀�X�g}>�HJ�Pi�\�}�1��{��	�#z��������ZU�cJ���􅋦|�z���
�D�݄ɗ#	�Øw�,��o����JLSK��`�(jy��(nK�XwE}Ş��j'^&I���VT����M�Fr�F����p��a���E�[��7��ߙbDZw�̄��j���]#������>>��zis�.����Uu�� ��R�3�֦��c2�����\�e�G��
�K����^Q����}[���$'@kb��`u�ji�]%���O�?�Sp��ǰ�b�<At_�	<u���G
T��ײ!y?�/!�b���#�dsPY)�� y��-ćR�J�yi�����t��%���76p�w���*�R��FRO���\N&��)0J$<�Έ[��.�,m��V����X��z/�[,#�8,���`�~wݹjj>�ohW�I�����0�n ��	ic�9-�Nr�����waP�ھmL�\Mx#+�;��NSҸ�пGf�bw�jÔ����R-�OV�=WC����#���i�15wm���z�6�%����u��w4VNȊ����Ys��C�y1�2_���������'���9}�T��r�	W��yZ�Sf�y��M�&��.�E�w� ��	͆���Yv^���	UwA�:]���T�e��3�*Y�WSC��qQ'�����*�YK!뭐^��aN%�}uR]j�	���۴I�x��I�[_�Xs���<f8����B���Ԋ�����6u�>��P ���Gqu����Ix���~������hH�0/���<�td�s�;K��8�c_���R�ˉĜ��-wݰ��
���7��XQ��vt���U��ɾ��h��PAQAⷎ��F�ࢆ��{���"���&�Q�q?��ꠉ��\�O� 8�3V�����
M�pv���+��<4���4vuֽ���'�xc�Õ=�dcK�{Gga�7��9?l��D�	mع�'��H����й��}��͝z�`�lKn;���
�"Y�7"�E���%=s�/Φ��8��٫�
�2�<;#!p4����F�GFI!^�'�6
��"Ρ, f�	̞�wo�!�5np}"��}��"� u��&|�8s�HN�������Ɗ|3<?�R�b��@�va@�c<����wl���  �Ԓ"�3�[�zL��Jw��㶔K/�W��#�.�������pZQK��ڼ�������s����*P� �IߕI{6�CL����Xr��b��r&�ޔS�ޡ2m�!�W�Ǌ����+=�װO����$�(r�]�_��v(���Wm.����uACߞ?���oa�*� c�.���CK7tC#P��n�����(:`Hn��}c����lU>K1�^��.���G�;�uz�l]4*wq:�����I$Q���E�b�����^pö]E�I�-�ÜHF0f�+�
�~��B�۶�;5���DPb�2����=����,�޲�2�X�;4T���p j ��v��G����g�4N	�VN[楛RS�3S�V���9v��Gt�TI���HJ��y�]�7ǈ���_wuu�a�`�o�BZQ���M$��^�	��g���M�)�V_@ܕp�s���p/$�K�o0���o��G�ʉ���(���:��6)v��ԉe��4�����]���o�|�S>�L��� ,x�$�.�!f`���#ݙ�T������R�qRi(�N���7+|����d8��-�3��������ܕd>W�$t�Vf^�+C�o���s9��t~k89W(��^�-{�h�u�VZ0"
ڃ�V<aUN%_>$�L3��t��C��y�m�aH�2� �i�Ec�A\#���Ԫ�3�1@��O4�?��zYǹ`[��Q��m���y�p=��h�ne�4 +�n5*=XB�]���r���6͋N$9�lI�EO98�";�^L�õ�1����m7��n�n�c���p�DJ45#��'��[#j�2�`��0̧'���lM(3�d�<1����� �:3Y��\|���D�z�*G�M����깒�^����M4��未����)@Ts
�Z2O�b�%q���*BWQ�a��� �o�L!��B@��H�E����`Z�kK�X��R�'��o���IJ;��z�֍ѪL0�H�Re�S���>���[c���9�w�%aØ�*�O��Gg��"hh�,��C�ҿ�>�my����;�|hP��ъ6B��C0�k*��j֞�={�h�%r씢���Z8�k�%�{G�ג�{�W��7��B�)Y���#^�]���N����X���=��}Bi���`�N6��ia؉�?7�������{���BXA�^��t�j�me'L2kٺUlDd��>Ȍ�T�gP�Kl*�w٫G 8qe�a��zHb�ͅ�2?����%cNVR�8�{�D��iħ��3|΅0Z#�h�������\N��YZ]�G����D^m�dZ>�u'F$
�&��@D�1�x�
�0[�����UR�.ױA����Fz�1�}���i������KIV���{Y�J����*����Vo�|���>6/���$r32!Ɗ)726�*�?�
��w�O-�����n��I�l<QY<�l�Y}5�В�N9~�"�������Lw8�	�?"w��qW�W�D�&�I!}�`�5��Ҝ��V�,=����L�TF���7kV�{��0��Pk�� &	a7�PI�a�.]W�e�v����L�9C/"b�8�
r���=+�z��f/!��r��*2����xvhW³������3�R�	��a��� , ���q������P�_7�PI��ʼ��٫��p�_�fߙ�=|FH�!�u���-��7��� e�{JG�灆�����c��Lw�[w���A	ds�iq�rjklsA�A�/�v6ח�����$�;Q;hO��aCJ'��j�p���-=l��ꏚr��,��hcż,��`�ʢ�¬���	�n�!��
mW&�,i�{ef�!��13׈�%�g��gܞIi����bY�j�H��(�K�fW��%�l����~*��YRU��h}yi%i����w<<��gBKA�b�`�� �D��}�D8h��:����e�q�p�M1��j���i�G '�`����
ʳ���>���c�c�`