��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�x�W��$�oC�Lw�S
�,h�eԀ)�CQ�_���o�E�'+��l�����qz%�[LըMū��ş��Yz�g�#Vz���E���_�����/��'�w|g>ѐ�=dC6����	NwJ!�
�PΙq����F�<hŚx��#��aT��R��`v����*>wEb�3�4��	ηto��b���RQX_�?+��M���C�ӛ��/�7X�FՃ���W�"�Wa�'_ ���0��a�ߛ߈"�|J�0�g�w���r�~����"0-̦_DoU �0�,���-f��!3�!
\/��M�;�P�[ni�s� R F|�h�[��UtNi�qDۏ����F�N��Q+�9����f&D�����Ш�q�v�.x�a󖷮�]g$�3��|�jWu�m�lB8nB)
�
:�$�y]��Uhֿa�dfp ��:��b��Y�ٻo���i1߾x�B�i��F�"�<0A7l$&������y�Vk����1 F���C�l(*�]}Ԓ�*H��*PPm�>�Z;8~[���Z��{H���^��-���؅��ʫ9di�����K�vk�E�:�3^t3Q1F"�K����>@�H#����]է��檹J���7
W���Z��c��<?��_�[d{�ч��Ϩ�lB�����A�捳�pf4{T\K�:j��.~�����l)��r�^��y�u���s�:$Hh>���	��'xN9��yEySSKҐ*���L+C�4�]j���*�ŒqK�KYeU ��	���X�Y�C�v����]!'XK��q4"�cE>��q9�����2įP����?(�"�{�����,l�{�?l�7�`�@k3L'�����2u[�*R�����V�YN� g��}&U��KG5��[![�@��bH�<	�� "����ޡ)8��0>u�$�U ��F�Zd6��E<b� &S�|�� ��c���i�ڑ�A�h�'��vS��y��+,a�OG7M�ܪ��̮2��x��y:]�/���>5t(m绶Q��
NqC�M����a3�@IHb�).[T�|���L�ʻ@��rk�6��˨�S.xU��x�	��uo��Bf^�-�;��J;���@^��I� L_N���̀v,�Дm����+P�-]��2���$̽g�*��w	R_I�q@Pdj��:'��am4y;�$���D3��
�"%I^	7���%��oW>��wU_i���״������e��=�����w[���%��4/��,T���h�`��Y7L˫;�VW[Yss���&���{� �al���ۤ5�J�U
٦��o��=��6�9W�h<��2��8�����R�����A;?�m.r�)�3�|P�Q�]gC�;��GY��v���@P���[��^-�1�����ż����S���'�d�zv�"H:�`7M+/ojT�3!>g)������N�F�����#&�m�Ͼ�ɸ�2���ۢ�컬�m����Gc�/i[�@��};� �ug
�/����}�F��:��[P9TfZم?B�iE�	��ˤ��������P& %����Ր�L�DW�L[N�����u����q�����!u{����O}^י?����/3�cR;=U��cN��Z��o�v�g�b/3?�-��$'g�v�T=e������q�K%.l���k7� ��ZLUW2f�J0�2=��~�|���J|꜃��k����˦LR�L �x�"�<9?�uʍ� B+���pV���Ue�5Fl���1�������=ę2o]Q�L*K�)(rm[1�Z]��*������ڶ�$	,F���P[�"�D��!��%���s����/=b��!�h�W�ۈ8���Hʄ�{:[���M�l��$v�a�P��ƞ�g�5�}��2Ţ	�n0+�ȼ�l�ϊ'\M鹌�q��N�?�F���%aG��r�`�.�'��Q��D�}l"�g������l�p�?��旀��p��a�*�ǽ��A��M�/$j�Q#V�R��,"�b��d�?C]��5|��/�{��r�{�wN��ɥ;=�?��BK���L��'I�38N��b:�J�
.��^�\�z�a*�TO���*9���x�	�ٷ������]nN���^>	�D�����tP��v��؍�E:����	����%�L*i�#8XBK��������+ܬg��~.��`��v֯۽z��$��\�`�����$`�_�ֈ��`4Q��+��-��d��b)�#5������y� �����K�,7����f�X��`=��N����
-/P(P�-��W8��UEz��E�ZBfw�SM 9����?~<��W6��)+(���R�Do����Tt�%3^�XEJ�Z1m�� ѲQ��]��F&�S�)~�F�t��W��i�#�8��Bc4��ҠE��%��i��p�����N�]����v�.�e(.U�5E���E�M 76.&~���my���-ZΘ��noV���#M}XG'-AZ��b������V!?�} �W��]��<�W>`���a_"y�����+̳Q��8X����Vg\����B��� �'��L�J�A�H�.'SϳV�>��E�~�|'�>�� 5���>r͸ﰊ��V����O��䛰6&����4�Y>�@����%��_R��S\I���W2�Zr�f�e�u@;�)�Н:�IR��J.�{�Q5bx���a�u�X�I�u+�(&!��zL6��x�%%\��t(�P��V��
�s�_OJb�����[}�HS���ct��ї�`U�& o����@�F�^�����JP-P�?�%Čb��1��J�]Ow��G3��tQ��>���b��=�<� 捇�0��
J!j?*g;W�.%�
���y��'	l?��z�b}u�_�Vh��x�9j�5h�+�{%IwX�Ȼ-߹�����,�?LYT���[�Nrw��գ�Ds�<��Mgj���]��p�O��g�b�'��}3`?�H���4���K�_ݿ�����!���%�t�f�ɥ��w��!V-"��=0�xh��D����#���Cr�̓"��;�O��]��6�' d������6�9���[���ed@�����4��)��ޫ-��P�+Ϛ�m`i3k��-�.��A���w'�%[�R(�2� ��ٌ��󺇭��M������di��Z���\A^!<�+��,.��y߿�n���_]=�f����o�O����[���WM�=��}p�7|��*Q�#��T������`:{��R�ܲ�DеQ���׷�� �/�Am����GL�%yd�}�1z�qfb���r�1q�v��6>6�ř���e�j������s":$�؋h*��m����ъ+3��:r��R��]�VLQ�&�_
~J�A�|}n u�j��t-�]��T��/4;���) @�`���T�l�XHeǪݎ�eqd�
�~�nyׂч�ōiZ2Yӟ���Hև�((�P�e3�f�y0ˬo5�u9�	���N�(�����@�D8gJ ��}�~S�ɀ�mt���Um4��$�&唢+����`;�;ˋ�a"��	:
=m?C�+��fǳ���3CBq�J}Q�Đ#j�#��VA>��ե8o�p�S)Z���<�o6���cr�a�4��0)7�긛�P��{�w��:�-�j)B��d���� ��R���ឮ*꽩9��19x��j�̶w8�(Z��ե�-�GN�xy�Ê��Xa㈜r�Xh�_Џ+�Z)O�L����=�Yk ��-�w�l��P|������]��D��B S��~�������г�����Lbb!�A$����j�Y[�g�3�g���-������8�n�?V���w�vh���%*/��"�7��,�4J�@��u�{����T��쐸���>$)�U��0�×�ـ7t��Y�Sb��61��0��_0It&�`�ٔ[�PQ���'G=�48s��C�`����t�V5�e�F��!=n��0��Dp�?�}gߞӤ̈�5_լkM�軇��}i��A������e���$o�SQ���V�!z��WBPǽ��wq�U�������砐�U^u5����;����?�
�3�wv*��Z�'o^+3L�lqI�?��O�v6<{��
�̢�ҋa�q; ���J&��,Qq���D
iᾮ��&:�ոzF�>�j�Zg($�{�3
C�p�Ш	��&��L�z���_�ȡ
nm#^���&�k9F����;�I�<;wɂ���⣱�w%P���P�u࣎����P���z�DB��Z�nW��8K�U�)�l��{*9�pwDt�ٝ���w�4�B��/�q~���ӽ����:�ϥdv6��jЬ�+�d��Te�<I��D�M8`f�