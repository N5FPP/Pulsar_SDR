��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��e�ik3�������w$����g|��J^]،�[Hވp��L޿�e=�/��h�8�,=��2ؾ+!�r1O�uN�&��`B4�Y5,�hp�AJN �@�@��#��>�z���f3Њ��b?���-�>z&�H�)w��ȍ^*���(�>��N�߃�+<�Ѓ��?�^��J��HT�K�R��K�3�R�vf��u���$�10�uJ]�	xF�Bg ���W@�mz�60���Ґ^�8r�8ÝS��Zmp]}�Fn�{�g��#�2��S���K�v��@����-u��������RC�T��j޴C�!U���.�ک4:{`7����8"�"���i��R�v3�H�b�xAk6:ߧl��$v,�E�JLʇ?
�P�)�J���~d,S��7z��9��<�gO��n�x�����m忋��]Y�~���5B�CI��Hp��zA���#�%d,��D��w21��@��z��{��}��5r[,E��
��G�p[+mI���r>��;�£��M%/�5.X�ƽ�i�P�ɔ;?Wuٹ'�s����f-�$6sɹ�=U]���ֵ��]��-e��G8ѭA�R��vЅNx����HP	�Z�Y��0u�W��KL�!�h<xhe�Y%����}�薰�����#��*��v��u������ι�rl���r=��^�<��6���"�@V��9˝��S�^m���̄<�-��D7�����%PI����AM[�z�@٭�!�*�V��;��mh�~��ʘZ_P���4U\	G����d�	4nc_ț5��B�����lczl��-��N#�C_�����ҊJ���Ň;���sN7Q$�!��,�F�LeϦ�Pz6��)��'
�3���y�����[h���t��H#/g&�Ӊ2?[�21)
�^Јc���Z�P��a��Yq��3�w\�W�69R�dAT��0�\��9��F�V����?�ӊ���&8菖O�:R�n�Dk%r�P���\�{[.��H�*���̋8mý��W�,�{ч�������}�6����)
�n�l�'.��~���#Rq4-�3W�qkҞ���9;��&T�� ��I:��QD��+����s����������ʂ���./�[�@�`�}�uL@a>��~9�9�F��dn��kno�G��u���9՛��	$��V��� �*)��fi�ڥv6r�;�ߦ�s�DI7��i�p�ONdx*�C�d��E,�*�N�����cJ���V�>���8~��g�7�#��d'C�3�NsX��V-Nf�q*oN�w��f�9Q�y]��G���L�]2�3C��Lsix8(ފ=�(J�������t� .qR����Kx�w��ⷬR��h�y1�x>~��T������)Y#��,*2`3�0�*��ǣx��h*�ZbڙP����a�����2ǉ��BIȧHA v�<�{�v�&�6�-��I��.��]��B��dv�W)G!��Ht���( �Y����[HK�d�%�]�C�۟�p�`�Z���ә����'}�����e�|.~�,��'}9��?���C�|�͛�l��-�^w��G5��ËCV=5�Cjx��a]�{龧�&��M>�H�A��}�����������^��K��L�\�J[f@f�v�H�C�������o\F����BYZ7�dw�,˶��-��jH�7�}����c���u�k�#�G;��n���֘��+P�%x�N�,	�#����R���i'���@p�|�;L6�C���Q%�ZI��D��3��(�\*�(,V��S)L���5����ͳ�.x���mއ(��bc3�IS�.X��.��h���<.�mM�,��}��s݀m�K�H;�A��m,��[ �S���,���k_���b	�ncΰ\�4��ߦ���-j�Tn$W�����^�yOO&d�N�ij���e?�@ϩ�EG��R�E"V2�g\K>U����I���p0��c1h?���ۥ��M�Dʩ��}Nw|R��+m������=�{�ބTeL���ۊ�j8�r����_0�.h̚ �d�`l;��]�虞�U��p���6��DyA'��b�{)�|03�}*��ۣ�?�e8k(N�S}��A��#P1�*<�zx���ec�)��x-G�$�ʖY�P��TG�t���/�.u+T��97�§.��պ�#j�?N (%�	9�������>��Y�"����?��^f�S��&O(�a�����<�-V���������s #���Y�ۿ���ʯ�I��5"4�A��e�	2���v愘��<�&�<��Y��c���E2���!VZ��[�r
z��'Fn�!1	�HH�Et�ɐ��ئJ�@n@�$>��5A���M��_#7�{)'G*�*c�9�_ ��ٰ����6�B8���X�q޳� ���Y�3���`���[8��T�ٷn�>�5�o8���5�My7㑭���y�ys,�*p���=#�V�v9�V�4��3�[W�Pf#1��;�u����ڈ����+PUvW�_<{ul�c!��hvT�l��\f������%��}1u���p�̅�]��[���Y����Wf.}�/�D�� 4����=�-H(��Z���#���̎c��8�BsY��^����Oo�:��Xf���e�Zo�������#y�n����������Si?��/�-:�a� �lH��ų��2����C:*�
>���Z�scǈ�sJ�l��՘�0H7��F��'V�����k
���!��2N{��q��y�&~~x�����ۂ)DdTE�]_�hD�fg�	��٢������$�EÊkq�F2�ORT�����E�>��]�m��ded�I8�p��nX|`���P �W7FE��A 
�i��l/^]��:���ؘ`��LZf�������SXr���Ϟ'�`��η��3���N�Q&a4�>����Aa>�s|�G�Ǔ��u��Q��_p�,�6�5�(G���3��&�0�7-�㤉4xݧ�H�	�oA� ����:vҜw��Oqp��>�t�+Yqe0����3���Xi�	��9���0�䆂YU�}�
w6��0`y8.����uB��	�S�m�^�wu�`���a����@0v�i�߁�����>���'� :�JVP�f�<����r��ý�(��K��YH�4�9�EFlD���9��sG㈞l
�5L9�3�i5��]Ԃ���	`O��ȷS��&"�"�[��vD%�YݣUn�p���"���x"3eC�=�Ùv�3��@��gkߎ"���.��4��|~�~�;t����rކ�Kf��M��R aYO��A&=��g9�xv����Ee)�-��Wd ���Üi�:Ybqݤ��kz��"�m�z+@�TB�Ns���T|~�v*a�.({&�i�Qrz���ܒ`�	v�4����o\��e�8S�����5����@��n1(Gn�}��q�<�OaB�̻��2k�{f�>��%� ?Q���)�����54$�b�[�J�N#w��C|HO��ץ�3�
h�ǚґ7n�8�# V�Ho�6E�����򳷮)�J�K�<��mzF	[����\�[�.�5�]��WMB.�r��\ I7�6��|�����ڂE�:2��4�a�Z�|R��?&r]��;^P"�Y����҃GV��65:2F	Ur2�����`�5o�Ɯ�;$�=$���ѫR��h`�cdh`������}�u���*�f�r�@xP��7�I��
M���|����s�oK 6u����6������<�X�c���L]^��$p���[x���{G5{T̩VGXJնI��b�<�fA�v�La�`�Ԭ~�2�����}�A���)�C�--���U�iκq�m|��h�7�qp�⪗L48�]RQ8��So�P�&��,�T��jÿm�\�_6��0b�$"A<�T��l��B�5���0g�|h5�>d�Y��g�+s?��?uY����� �s��a���I܇�����@�<-��B(�g�&Õ���O��5����+g�dU@Z�TfE-����9��H�ek����wı���aj	�ߺ����`]&e)�O>B�~���[#������j�\!�ڋ��QY(����&�+t��RAQ@�����vSv��in�V5۽��tܕ�C(�U�2*�^oⰵA��G�3��Tex�xՁ�D���.Dq`��_ӛ.f%�}��ߎ�\e�F�E/[-P�
NCK̀�دtT��6I�[S~O�]�c��V�if���@�G����|W�>�uř5E�$��U^v�D��z�j �@s��f���������F��rX]S���NQ��x��p�W�>�?�f�M'��N%d<�n����C���,R�{�s��_�` e9�1�%�/���JC�!$��d+�2��D
��\/��[���esWԷE;�(lo_e=���d�2z=]��U
�Dq������dٸ��D�`^l���ZuW 74mU�o��0����+IJ����5d��qK(��4�� GGY���W����$�NU������Нݽ8�L9�νU^>�pT?t��˙��w1z��>�/JҢK��C��P�m쏎OT����'��c犸�$p�_p��HF���Md6}�6�Zy�e�4��J�(}�P��0�>��K9��g1�QSQ��C�
�p����x��d�.i=��*��Q(+�1�}����^1�$�
ʬ�z]��^*F�:�����6��&�p���Xk$3E�D��"n������������.������ʀE&����l��#j�[?4�0��j��n�E��P�v M?���&BHuu;�,h�~%p�F<�t��p��������T��q���������2��Vjt�7γd�l��%I\�{��i��)�p5
]:�e{.���#B�6)v�p�	Z�Y˶|}��R<���5)i
��4�}18v܇�r�q�?�C�������@�/�O��J{F�`dSk+)���)$Σ(��m9�\ca���,P�_�%?��n���ߵ���	�_���s�.���Z-Zw(�)f^7�ZY�I8�t5�b6�x6��b�,Ǟ���U�Me�Ӯ I�S���;'+Y*yaى�`���3ݚ�">���D�I4'���#��͙{q�磌e��>�*�"�ﲐ��\���ܒ�=x-�>,�����?�Y+���������"+W����7���
�|d��?����t�F~�j����5#d b�aS�8���1�4�U���z����r�L��@�p`�!�����[���ē�u��%K׽G�yk< t&���� *~��m� !�
�'9�e�i��W|x��{��ܔZ.{{�xt+�+m/7�L;���yt�o�F���p?�E;^�-����������׼
��"�@5����=	��ۑw�Ҷ:�|g�N�'c,�`Z^���AV��1�`i��y����CǼo*�4�Gq��å����(=������7>�
�L����9a�y ��V �NS�"�z��ga�C�g��f���ۺ��?�הk�q������Ț�[z,vf���� It������|����ı���Q��Q��\�D�Џ�K�Hrn�� �@w�kQJ�+����x�H�o)1���7_I��Ev����t����5|y"o� �+�nԒ��(B��f�U;+��-����}}��rE�(O�����B[%�~<��`d���L�M�����p���m:���J6�hg� @�w?-�vh%M��k�bf�#zp���d���d�Iׂ�Y
r��s�hE�u�m2��<d���\�>]�{��\���d up!���#q�1bQث.&l��+e_��^.CV`@ ����0�`��g��읒Nmm,?�b�l��9!CV���$<[!����HO�-șL7��厡�e@xm��~���l�%�	�D9~�hP�n'������>�w 1,��?t�m|Ӳ:|��s�
 �ߗ)_h���z���-����o_�9Ǘ�(O�^��[��V��ɷ[�oi�I�� �a����QR{��A���?X������ Ǉh���UN�f�وI���L/����Ŀ���Ps} 2�@al?�O��&�W�%Gk�����^�Q�h���Z�	Q_�,9�(V�'��*��wr��7W�Lz�A�>
�)��_փzZJy����D��u$�|��~|�W�4V�4SM4�.����hL�Iz3r?���F�4�Y�J�CHY�
 p����S���J������z��R_�u�)�2Tl'Sȣ����JD��L��,��<�X���M"5_��eY�h�%�_P��Q�~��$[�|j書`|����D���"i@&��@��:��\m��)O�Ri���07��`Y��	���9����7�K�X��콇?�1����bʂ�1��r�í'�/���f �E�)TI:���L��~��G�!�]P�s��T��x�,��K�s�=5U���EFt�,�jS=0J�g�:���|fz�.C꺮�=���y�$�s`�n�!�_��e��%��#��:x���첣����||�\8A;����d���-E{�QF�Hcͩ�Lo�N��/"gt46	��Y�r��Z~l�"���(`��\Ҟ�7Ѡ���8�h�׽��MQd�;�0hv\}PrGloH��S���>(йF�@��|�g�l�{�0�ʚ��L/��(�b�5&�J�e�h���qÝ�)���=��:���t*�5h'�I��g��-1m!U�w"D\sIyC�,u�k5t��:W�d��ﾡi�j|Ő�S����mpP�xK�˻tB��-�89�U@Z��8=�x�n؊zM:��G;>2f�%z0GK���L�0Q+�2�Q��_4x���V�T��:W�a�#�u��z��� �@��]	�od���ɲ/覕��lˡ��^
�W���=��r��"������m`��H�i{������_��?�c�,8����,%��
@}�TC�C���w^l"ʀ>�؝W=I8�e`�4s.޳�9(�P�u~U��5�/.���Nu��)�">��������\4SJ��ԧ&~=����%U]��h��Mfs0�+2����ʌ�]��[H��0@D�%�'�_ˎ���W2�D7UN0����C��`C�0������g�'�x�6;E��mv�����[��e�y��A���'ӻ�8\�H�K��O�B�k����*uD	~����Zj��e^��N�m�p��ݻ�q9&��?�Ɛ_��W�ǂ�O�?��Z=��=�eqw����l�c~@��7��:c�T�|�)ޯ"Yʓ��2�'0��b�w��5������DH�㸢>�)�#Źe%���gF�t��p��+a<
��K���`!?g|�.�{I-�z)�s��]S�w��Dŋg�@��Ӫ<=mpOG ��;�ªI�]4B���ұ#���ie,��D1G�� �~��]�����%�_�8�m���{U4|�	_��cmD1���������Cfj�\�Ri�es��?1H��(F�G�E&�X44I�i�?FlҺ�
e��ioA�i�/�}hT�����Uf{�.�#ͯ(2R7�qk�Т�ȐGm�H���,�)��E��a �Q�����J�6�N�D�e3�^�����X���guO��h(7>�S�΃��D��I��_6�ր�[��w7«�zMy��p��Q�i:%�������Fe� �#��d�;mH����(ت�&�a��1���d�#�r�z%���AKmtXj�w�ǅb�p�`�����2jx�cl�����ù*��W���p�P��:_��s�6�#���=K5�
�F(��C��j"ͳQ�\ŶL�gữS%7�o�.���#�;�VMh��M��[�N�tG��n��X�N\?ٖ �_��ګ�9��§E�5��p_^s�!��Y�7As!��d�h�-����-.��('��hȵ�FpQ�>�
�؟�Gΰ����N�Ͼ8��jq6|Wy�F�
U�{�A�F@�d=�O�&F��9�#� ���E��3e����m ^��E-"'�5�kas��~%�4�vr�	�18?��f_e8�7X-���O맢���O	+����	����y����(CI@֕+�0�z�n.U���ۙ���P���%��o���l�Υ�{��\�b��
�vC��To��w���r��c�k�u���h��;�pw�=�
����]n�(b��?_]w#�/&��߯�f��Ќ�3�����6��|���c e��}�=v�:��ļ�zW"��|�2�1�_ܦ�������3LV��Y�<�Y����E�{�ƌ�Uј]����7y�b���A�|��rﺈX�e����A�cu��9���Nʈδ]��������4u(j1y��ص�'���t�,��)c@ɉ6gA��m�X����*^�U� ���e�u
�ք2|׮�E�,y�3�(N�,��?=J���V$�ؼ.c�G�)�ހ1}���ѫG��0D���%$2)�����O��ne{Nd�%�V�2���/5�?ë�6�=J�!�?�1�����L�9ԡ�;{��
1El�\o��'�π�Q C.����b�N83Q���(М/kx�/��qa}!�����/��]��pq��p�#	����t0�������͹��v�Kc�|��T��ny��ɧ�X����RC�P1�y���X���#S:9���U��toF3Ď�f|�"�1�T�|F&�V0���VYt1���/�����Aמ�t����,ϟ-�;�5.�y���Y~�~I�\y�����ti(*��p+�eyd�-���A��Q�-7��1r���'���,��WQ�"T8�{@�V��9�
�� �實��P�> %n��T�R��n����!맙ݏ*�H�m��u'Ӄ�oj>P����h�� ��m�~���F3�=���Y^���CŮ���f{S�6OZ˦^��#b�C�h�--�!��d&Ѐ-�-k:B����Orfl��eL�FkP�S�=n���<Ћ+��Ic�&�pR)B4�%��s���jh�'�����k� �<��_lP�*��0ӗ���x��1���@RB�r�	�<̒��^�Ќ`RCcXox/aӰ������)�Z^�[��$�4&�!F���y%ϯp��X�����?�9��?�H��ra/�zD���I��Z���%���������U��	|{���FB�ρ�>¢��F�2A��tZޖP�d����C��=k�$�P��m��V{�k��p��_�j�[��{�K�L˲�G�.7T�6���0��~����E���K~���uns�3)��i<����a��Kb.!�r���(�����tP[/�l��',�JY���}��X�ǹ���$�N_>5�\����� B��< !��"Zv�	�[���;^�w�p$���k�e���t�>�s��bM�E��0�)����<�)=Vk�������\�c6���T��H�-7��v��	s��ID����D݇�i���X�9ˤp-. ��m|���8,�ЊMe��T�v��1�nSr�j��
�E�	� X�N db&1���DS鈹X	0� �$�ɝ���%�.O�D*`ܲ�t������=�r�e�л���,�5��U%�[��z1C̓��@7����#�����	��UC	��X�y�[8<xpJ1c�ў��w�=h�#b�:��ְ���׊T$9�3Lu��q��ЮF���5 q���i4�+�@$�`R�D�>Ğ-P%D+���__�=uobG+��8ث&(��dL~�^~%a�f4��r�vs)#�B]�3�׻]�F��80<���!���R�c.�F�w�EJ������o���B�t�3���
^W�Z�l�t0��-�Z5��I>�>[��C�µ$8�-=Q��-��}_	�&H.��F��B����<\�4U��:�J�S����˘�y;�������Xj�U���\w���^CYfn�"��,V���O��I��p�/��Ƶ���`;S���
�zcw�F�^lM�-�@�q^�BC�����Bއ�ս�,꫗]��'������/i�1�_��{߅/���-�o�_D���q^�pe;�x�7z�wY N�'���hw�{zk�:��Ւ��Ji���E^Zy@������\�Xs�<t�7R�ck��:���/��n�qwػrߌ�N�@A�T)�!D1E�@́G2���v���5�#���i�"������II����14�&�2��T��21�.LH٪���䤶%�.v�/A.���C�86����P74�� �i�U�/S�Al���2r$���8q���
�ǁ�҄�:��V�h��Cq���ə����C]������U�����}����� o*��eNY�l��57��pH��[H�t��jO>���.|Z�*W�y�<D�e�/����-�%���f_��a;������i#��� K������J�2y���vm�K�٢ŚQ��}Z ���s��\M�W�Y"�sM�7�t���u!��Iv��Qh+26'2K;�z�	��M0/q��(����Ϣ�}3^}#�ϓ@^ٕ%p���靬�ax7� Ѯ~��FlؒӒ!N�����|��7�LK�	{챫e���a�%c��+V !e���cX��.ݒF���Tz9`���It��ci=&����I%����D��
(A&m��,b�ݹ�y���-I�Qs��X��Я��Z%�:�Wm14M ��Y.OF�Y:N�L|���|Fo2�5l&�DaâC��Y�i��@�R�+��ʼ���T�����^[�~MC��e���!^� �z�Ɔ���3�S
ݟG�Z��,y�4Ue�|�7�i�DOB��i{F�=��lr��f�_����Pv1°��@Z�#t~:\�S��ˢ���d���������ρ�Az����Ь$	���p�eU_��� ������ʃrO��"1�ϯ���X�"�+�H�^����I�����*�����oa@�&�êXp(	n_�eN"�X�ڄ�.�<bN�
+� ��-�a
�)gˮn4pV�kb;'X��k��g��U�$�::]}��Vx�!�e�q�s�+%$XU].�p���ꧪX�n[>��T\�\׬�TR�Y(�K�����b�*6��EP~��W����P����A�D���������e������2���mo��k�����N���A��0*���A�Yf���l���uŸ����/����0*Q�6(�PQ�m��B�e�ȬdE����cj�����x9���OI W�D���t>�R梤>̌Ѕ-C�u,��"��ԁ� @�]h�c�W�~q����u�M�v\n-�� A��>���H�t���~��A�w䄙$}a!�{��\QMʺ0r���"&�;k��>���\y������GkkS��]�3�Y횈��C.A2������� �։�VO(��iZ�v����c����O��f�E�5;���%�F�E�;D���d
���G�W��[X�8{
黓���eE*]���=M��P'->��Wx��TX8�!�i��o��8�KJ,O	�����V����z�' 6���ب�0����)�^�C���U#EE��ãX֟���T�w�?0好d����X_�! >6��zX�#�*!i˳�$�qY����|蠩~�s�v}��?-+z�٠d��Wp�&�hy\�ѓ)������?lnq��^A�ж��� 鿈#��V��Ve�I+�����t /R�Fq��b�X�W������=��'z�K<%���(쟤=͖}UC�;e�:��SA��3֡#A���..<�fr%?�D�^IHi�,��R˦>iT�b�\J�z��՜9d�V��L�d���$i��Ü�����!o�o[2;J6��R�$����۳��C0軚�fq\��1��t$M|�dJ�#� <q���RD�Ks�*MD⺈�)�'�K���)6����Z�4�O�6$�7��#�Ɲh���C���g�� L�){�������]�|I����!�e1���'�LS���g�9���T䙆[/C{	�����˹=�m�j��"��[�
3��7�h���4���x�Q�1ӏ|�>�|�$��Kl�/� �E}y���PO/�OBB~j3��ؠ2?!μS�	�&�g��BP��H)��8�������T�P����)�;/��
�x�9�ƀ߾�š�|�@7U�)�y���9>��.�o��� �^���g�G�-2���x�@[¢��w�G�J}�J<@�ua*fɻ֓N����bF(���f�T�r��QG�R��RR�"��9W��y�F]���f2�+�,�V/�2h�7V,��o�Z��4�ʒ��"������l�ϼ�*�Iw��@���ǝ���� 4Ј�#רR?�!m ���x�|��w�#%��{�$67��A��i���o`}�力'������i�:7��`$"��K᱙R� gg��9-H��_ox� /�Ѡ�ڜ�JA@A�=nm�UI��]�n�-⍇��=�)�m�Up��eY�9]��ы���<�#��]���I���'���JA�V�Go{��@�}?�-o·���,�F�gdy�@N��K��F����.���<�
{A���<~��3��I[�l�b�A@��RL�w?�xT�4.�\��#�aK�jh�DN��� ���g�����'��ɧS�&Գ�O�P�ѧ|ґ������/�a�x�tR ~9�!i)<��G���U�I��9�t�D�akAgv�;��|�ڹ&D�LP�H�]7/����k9��=���&���`ϊШG	٘��� s�#v^��ƙb� �����u���w�p!j
Ӄ0��Ұ1�g�闽;�{H) cA{��������(3�׎�Q,��3L/�b:��
C9ڳ�'�}���\�'����u	�áԨ�`DMXÿ5Ì=/ƚ�k�{��w����bJ�u&|�FJ�4�����뉮(<I��qOl� �c����(���t���&�۞Kx�pt�7�/d���9�Ό�|j��{������j�n ���;q�6����+�*��$4�,��7�qĢ��m=�^
�4���>��f��4�B)�駀���; ��w�x}�O��{^��t{��/�ّ�I�6�I��0�7�r,1��~S��Z���dVd�'pC�q>�>9͗��u�t4A�%	'�U��d;���h�St��r������!��V��^v c/�Y����S�(���1}��ۡtgW��ҽ6f�t�?R\�ÛچzeQ�����Iǥ�6:*���C� Rt�6�����RE���y��_M�M�:d[�M����Ox��,	��`m���y]���/"�.�2��vu����8m�&�65i��K�8~�G�*�m2��=~�'n_n�$j� �M�q���67?{�[�%S��mQ��9����6�5���V4�\6������MK�%�Te�	�`9��,-���r��h?��r����TvVk]���:aj��3ۗ�u��q9�0{D�v}Rnp�wu�ҍu����/��֧w ,���`GyA>i.C��7�Fy�l�%،���Bx��g�#Q��o\1�u�����l)*��#�K�6-��f}I%�M���w��Uu�
7J"e���خA+������8��?t�ŰŔ�J*y9���P��S�dyxʉ��8sX����ۧ�_�Ν�\��Dj�ˋ���"R8E�{T8fT������I��L�G_�8��r~|w�6`Nؓ��4��� �h�,�b�o�U;B�=��$��wzQ��dl��!4�κ_w���"��D��������8�{�v�+���:'%~}�rl<j$����9ō(����<�v����v�V�Z;9R2F^����[~su3�/jNI�	�q�d��$�
��I����o�s@t�s|?^<�����RIZ�Z������Zh�e�w���62�ݩ�r|�Oq2�az$�`Q9Ŕ]\�#6e:�ZA��!�d���-�]���>�)��xe�;�$Ό7B(���G7�����ZKF�@�G^ĖC�컂k7*)W�UU�Y3u�M�W�2�j2ubU:A���l�䔬q�B0ޮ^��ҎcF�Zr��ޒ-�etiB�%��O-��y��p��Ǵ^a��Zf��6}����x�t噆So>�<�,��w���*�k���p[	�r����=]�X1A�d�ޔ�a@k��|�� ���k�u��������鸞m��~lCS�,)�[q��6Z�*���Mx<��ʧ��f���U
���=C�6�}����'��" !Ns��������
�OD2��.�1������X��?�t���-0E/���W����%3._�5b��F�?Z �E5C�q�M�A|��e�K�ɹ����Z�1��'���}c3Qf�����iE��]�6�r3�0�>zfxy����"�*��yzھ`k[Fc�~��x7.*m�^W�X�T��J�K�#�F��n�y���	�;�\��*�#&C9�в�%-�7p���
���1��bg��"�1Yy�=Mn�S��Ds��Y?�^��ov�Y�d���5�Kќ�@��"W ��a|1�j��(]�ǰFA�IC��`2�o"آ�C�LY��.�_�qPD��Cp�~�B�@w���EU�ǣr����K���ī|���A�y���J��,��2hqkL=��
��i�*��
)�D��
��\eң��oi^�qt#�B+9�4y S
yOz�ԗ!��dHG������ W�,��a��v0ֈ�����$8�Wz�!���<�a��N�%�?���3�w:I��@�m�QCnw� �
^�G�9}]��f��3=�7��2˾�+����
TzV�4�7��e������;Ƚ�p�O=b�v_�9&��PB���/u�����xna���4��kZu<�aY�Bg�y���G4�������r�h�DLU7O��o��qm�FI{������m`�b�����2+8�$�N�;64q΀�(o�&��7OG�ۮ�}� o\<Ά?i�v�@h�e������l�UJEƓ!Ρd�
/�GgY&fsr7��.���sQ��W�D��%�*c��Ч�2��Yd�Vr��Bƫ���o�7���GV�,}���E��OCz!��W�H�E��S�Ip�t�mb�)T1kb\߮��W��3�c^����:20ޚ^p)h�w�@p�΋��R�,��z�ʑ����?��˟�90N�-
lߤ
(�*8X-�П�
���⩪�D�B����S��M�nU�\)���Aў���r·1�2��I�II)�IӐ����,dkک����Q��h��Yz�B(y'	�ێi��A�K�z�%q��1:
�� ��͇���A���H������Ｂ�����<�'S�^�랻D�OPD۬�|�Ի����?�$-c	;��l0��2ԘL�G�oD4�]�c?,ʠ���ȏ��"��F�щ�A+ot}�-R���~���dPA=M�f�á:S���. 88��3�yƧ�'�c���akΓ=�]D�	��钅��D��"���$�E'��c8 T���v�Ϛ���"��հ��Ǎ!�W�L���{q+��\`ٻ�ޗ��)�ْ�G�N'Wt��h9��/#z YN۪����ӯ�x��
�dG�mCו�-�g��mb�t3#��4!�6F�Pv��-��\�����u�[���3�$��%�����(�Be�'AX�]��F�a�C�pF D���4)�c�o�������l(�{~��7����-��M`��f,�:��*U�r�3�B�ޛ�ŗ�vuO���@��"f>#�&Np��ɡ�5˜�?kE����9+Yq�s�Z&��nIy9�����X���D���y��Q$���P���t4��	Z�qo@d�s^.9Z�J�(P`�Ȩ\؏��r-��v
� (��:�1�WG�M>Zڿ?L��>��y�bJڬq9����p�+9A�M��S��F�уl�.Wt��Ί�2���/��ٱ�f]XF}8}�8#�f!��/�9l?�K�cQҘq=��%!�-1r�u*HYrh6H)�	`����(�H,fy6̛�D���=��\���z��.���~愈'X�c��4@Em�3��¼M]YcY�c�y Ѹ]�HڜD؜��׆�;8JP�χ�݇P["[2M'D�Mf����k~}����g�ԏН���SR�`3���T����(F�O�+v����~�&E�݄��ۭ��q|��.[Ⱥ��g���絮~��2����7d�c�-�'�.�)���K���A17(�;�`GE�8�$?��C|��Js4BD �w�X�Hc�%lK��<�r���*��b��X�6�F���L�?�ٜ�Q
�/=� ��Ս��{0l�~��쐩��y[ �<>Bn٠��³�9�&"y�Nr���!���U9�\�BH����}�M�L�����u�\�8N���)vm�쎨S%��_;�� m��8�/�k���s_���@a���6�0�7m��tH=P�����8�vUhE�� 1jڃ�Փ���AB�Ah���fǝS���8MV<݋��?7���k��1���8X.�&��
ꉵ&~&x+�(�}��]����K�=�������Q�#�˽��v�$�3y߳ ��mpdV��|e��7�tD?�w!�D�3�8��������M��_w�c�����[ҾX�H��[L�fz��cm�8��V-�ȭ��H���#={���q������qq��E��rX�%�{�:\	ZL�߂���cx��6e��R-��}~̒�sQ�4�74���X��}��V j��J�����uxO��y�����05��@o�.l���eh��Z޹���۴T*��t���&Kƅ�<�(��[Q����?���e�x�LK����a�H�V2r�f�k��K��m-��`y/ =���4�[�L�N� m=C[��\$�:�E��B��7�M`�b�x7���_`��3E�b�;�l��Ν��XⲷΘք-P"��0�^#���y{������a�>�&(}�o7�tI�tԓ� ~d~���s`I��Rw��x-�{�l����!�� (P���
,o)ɛ�q�q3�z��!~cۓ~�}%y���+��kW�i|(�s�)�kHAߋ�0������#.�&�����f����Ooٵ�k�:���(=E�g&#��k8���l�Q��6x��3�y�M?���w��BV�(����H ���9Z�p��H\O�S�mi�Z��.gb_�g����6�|���.�����Cz��)ȓJP0�`'�߱������r�". �j�ێ���f�{ycZ��L&UrϦ��%��Ƭ
!�����xҤ��N~A���qMmx�]�ҫ=�@���UO.E"��0�X3t���R� �Y��p7�v0�a5��G4*\�N^ڈ
/r\�p����ڀ�x�j*��n"V�Qk��h9I�ʽ��a;2OL�$�+�'x� M[�[?���XF >�
Ø3y%�)2��L�����(L���D{"ѵf�����MD�p�#�1Z?�	]**��Fk�����tsH�.Ɨr��l�I���ݸv�<�l���8(�ۂS����"; BR����{���=�Ȏ�Z��E����p���w��m[\��^�g�iO�!X�&l��,T�v	s:*�h����*p)�M�F��&h�˄3�U���*J��ۑ"�NK���`�l����D��;�mbG����$I0�5Wvި�M���U�j ����E1���L�O�U����h=������n�t"N������=#/d�#{C��o�_:��";��jB�Lp��F��H]��n�'�]�Z����?|Kz����@,.�/�0��OY�1��9g^j\9C f�����版G5ػ����wj��hG<9�p�Ǖi�u3RmS��u�-(����y���\�BGX�7��N[��-66+|Q��9�jEn��a��h�(U�?#� ]�͔Iޞ�m��G��)C�^��۩���8pG+pں�
�|��A��dZ�6��{��_����\���s:�tA�p���Ը#{c�]�ѽ7�a�2��	�
�BBۤ9i1��Ǳ�b#�(�V�C1dɹ�1�u~nCn�����|��2w��Y'3�kM��)z��OnnQ�!gJ�r��z�{��Y"3��gtX*j��������`��1��M�V����DeO�
�`=�xL����j�}�o����ˈR|�+�����r���x7A@q�����a���}O�d���Rk{�j\��M��7x�W5��}c,�Zא�Hw�ȏ�Y/(�\���x�&z�>�e�E��oʿуc��c��Y�Xk��.��`���|D|���/mX)�&��]��L��;�Ujú�A�@��B���uӫ�_W���*���cc�q���˔.[1��1�i��L	D��@�7�J�t��d&%�����Un���v�&��LQ{K�$����ʸ�+�D�^~�����������`�ͿN��`�æ�艞�	J���61r����|P^�6)�*:��_���_��NH�͏q��!3�m���EHL�-K@)[b�$�涳��Β�]">����&��(�u��1z�����\]�/|w3��!�G44�py�ڑ-;�8�ץ�ܣ�?��G�������g:?SA�TRU�֋���:����-�m�"ܒ�	ynUIؿN�0DO�9�ʷ���״g���V�7�`��#�=�4���Χ5[��QN{�}���L�W��t��g��s�ZfUd�� �u�%/�',q��9�J�k��!aV������D�y��gt���w����<�V�xu����������Ѐɢvy��2�"'z�Im'0l����(c�y����Zðf�J�:cu	�<�����I��	�X%DYVC/���^GAU��J0�������D���E6���*��]~ly��X�u�_i�::D���F�樎��F�P�?���Jy�`k�	Lg�
5����b7Kb���%?���fZzJ7���Yd�m�xL���AC�<Uc}ӓr�=��ί�Յ�fs���{��o�%"#�8��)�w�<�s֌M4�_�:�����!�	�o���K5A�i���K���	�ݾo���$���fӪ�x�D)|}�Qp�}��/ݢS�FL�He�]������;5�%�qg	��}�����C�S�q3�1'�	���dsE/4 �t6�E=�1��R�Y'�]I� Ǩv���r�q�(BD�5f�Y>��Ѭ��'�R�Ql�X�@�I�'���]�l�y��h����8;�noK�5���_�޳!&���t�Z��+�ď8o��+~���x׃�í�i�[ٺ�4�:�j�Z^
�l��]�eêS\�)!�������h�=.��]?�:�;njo*�b&�t�RrB;��y-�,@'�#}sY���p/1��d��L����;����_�����Ж���^�iV��F7�+��������5D��i�;�?e���ꗖb���RC����.+��.q%]l��Y��xI�x�iFdTǲ���Au��;�(�����_qZ�����MZ}'%���}/	*��L&es�IGt=�IQ̾,c�ڪ\.��ܪ[�����&��-�Wdx�������b�Y.ҋ�3ŃZPT��N|%��&�;1rȖ�{3��آ~�t��Ū������W��w%|�	���:A[��\����^�U�I��A�4_�������Y�M�"�(�ؽ�8y.c<�������^���2��(�w��"�r�Ʀܴ��;��ᐞo15��Lr�`3�`	En�B���{ف����tg&����������i+i��:,�mY{���=�8�q��'n����a�^K�W��#�<
�R	���G�Ö-�F���4����3ҵ�m��!O���K���b� ȣ@gJt�� �EJ�k�~'#L{����I�΋��m���8��2��E&>��a��ȵ4�����Y�1��_��ig�#b
_��;���נT�9i�6Z��Hg7/�E-N>��i'�y~��xA�m���)���Шǹ��+F˙J*+Jh׊YOY]a.�j�vTwZ��F�\f��C)B�q}!���]��������o��P�&���*nٝ�p�����^�m�\��{���<�uW_���Lc�`�}ߑ� w��J�m�O����늈���a�QF"�꧓�&b���^4�7����/���n6&&�R�{Y�S
�/���Ƭ�)����	�)���Ż.��^Z:�C�쨕#sv��1�j���lVĴz��?+�!'r'�bvڴ ����Gx%K/�;sӽ0]���^�~\?�T�aX��\�m���py�r��3�ŏK�ꭂ`�Q%׺�HK=���rLPxe�*�|H�	�^�/�AMA���8ʇu�n2Gհ,X2������Zi��H��Tj�N`���R�6��,\�@����0���
\x%�:j���î��u�F:����
P&�{�m�?Ie�c�ڗ�����6�tl�̺vd�����Z2(I�SZX�Q���FL�`^�.~��_.���ӟ�����} �*P_�����c	�w�X;��x�h(�|wW�;��Ⱥ�
#E���V��R���_��㶒ݖ;A變+��W��<܈�!,�b�@�s6�'���1��_��U���	��|[�^�B�_M��켌���jκ�)V"[���q��6p]3���&*�Y��Gypd|��|ǟ�j>}��"��H�5���h�8<ik�ο2"�.�v��yC2v6Iʯǳ�����*{_6�Z�j�쇥�\ ��o9CsY���!5�|�.!a�
8Gt���o�Ơ\��9�~ÿ� �[��V��X�kK!��������|'���+���*�����̭t�-h<����G@�th�?�ѽ�@ 9��\{}N�К6�.n�/>,|z�bw�~u��Sq��8#�{{��}��@�uT�K{7
��>�xg�&-�UDh�F�fy����F�έU��''�P�"���{�U�)�	�����
I�&���sO�ZP�OG~�pU�`F�6����6Ĳpd]:��I�P��e�Ѐ�B-�;f�1YJ]H4����ijM�"��!&�]�R�n�K_X�%�N�R������Kmss3��a_٭"h�"�ArQi�7�������֖�n�|��3���H�%T#� ��ӫ���8����\�쯀P�l*����b��C^�貨����?�n�u�cUe��~�Zҧ��uks�N��{R���n�C�ګ���3 �<�VN�>�V��O�v"�S���#Q��k�V���-��ی6�ǿ�d�9�IhO~7�c��u�0�iD���E�~o��#��G����f�mS�Y�诇�.'�!,���,���9qܢ9�d��7��v'�{���|� �B�Mꗯ�����_���^���gNb8���в���v�
���r���D��#�[Tæ�3IG�gTUN8���׮$2u��H���m*��s���&�J�d���/I?��Z����v�y�� c��p�QCnDJ� �@�#�,��80,ǟ�����O/���I
��4(�}�F��g��6;�p�D��?�wp����e�FP[ϐX�f��o������R^��@���2���SU��RoA��r�������?X�roj"�A��Yj1�k���1j�S��ݾO� �:� \*ԐP}B3�(�7�.,��"ҿr T⢲X��5��m\�mAf{��k�ů�R�yY�̘��g�K1�]uW���-��l�O����E+��X�֗��x=�Kx�ܴ6� ]6i�a�Q"�T�Z]�cE��xK���1��i$�*N����!�����zM��J��t�� )3Af�B���O�����Al�~��ﭞ|�󹋱��7Z�w^�e���C�����4h�ܙh/�09�s�G�'�$|�J�ϻG	<f�i������ɏ��<�0�Ќ��I�;x�T�C�g%��?��fL�I�L�m�i�L��sq/�b�O4r�Vԇt}?�V�U�:̓�k^����Q��v�󿇬t?d�)>��Kff�-��E�m@9#�a�<:Jz	rcs�u}��	�.%�d�U���{�� ���Z\Q:aNѷE���`n|���5m�k�p�=2e,%��"9y,
������ZX�h��v�emIc�gџ�â��v���ZS�\�yg̪�������A7��I��b�z����h�(�`�ǊOiw��?����z^������2����p!��`��tzQ���c<��m��E:X]xD����J���c(��8ɡ�:�XnAO	i}}͏|<��
C>���|�r<#� o����#���aۊ_	���
�L	5O,㔚�o����~3}�� �	�R�� 䜚�Y�?0����`�n�^a���H1����M��͔���R7��v~�L��xE��IChiX�Så)��M: �������_AL��������(.�I�1���>Y�Ћm��/F�
z��q):�@b�I/�o��������G�լ��x�8�ǫ}��4j��o4�_��78����I/%L�/�dexb����|��2xj�`�q%@��L�z鈔�����x3�%5�����}-�{=:b��4����������:�.|�����^lo�H햂�y'7��$7���@�GJr�aF��E��\�qI�~YG,:mEK]C��j3��%��D���J+��'��%��3��̏Bs:�P7��Qe~V�b9h��4}?ǡ3&~�{�67�1i�:�ɩ-�N�9�6�&e��+�Z55߃�E�� ��r�I���&�j�Ն)g]a&���畳��߈���՛���Z<�X^�%]�9ʐ���E���#1ž��v�9����̵l~g�E��?�}���}���D~��\��(I�1Z,��&�$�?zGW�S��������o���/�c�:M��̑Bd�5�m��Μ��hov����L��P�gB��cQH��(9�>Yw���@&$�V��N!�J�=�l�Zu@�W��@i�}�E�H+�@]���Z^ȷZxv�'�"Lp���������G������]�4�v!����q��Oo����Ne�1<�;Ͼpb�qj���Pyb�rE���}{��y �[�����?N�:��.��:�Zae��;S�q��W�f�����G��m��8$k8���:Z�P���X�a)�&t��c'ȣ���-/(�w0I�L���i6�mR����/"���W����,J)8L��bG�:&�V����;���&�K���AJ��%�k�HVFr��t�U�y9(�#���� �K�sw{�3��,��A3��kDt�B`8�3��\Z�r�b;�!�'Tg����FVS)�5]1١Rp�ĒxÔ��,rZ;�*J?=ôh��\���ң&����5��5���r�'ok![���ۗ]�I�^7�=
��vNs�N>���ߏr#��������
�h�x�,��*�&��KO�t���b��Z�0�T>�s�-�e-̲�P��D��2������07���9���\\[}��x�v����Q�p,�zo���dl�S�1�z�R���Q�T�`��RCjӲ������dȖg��w�j�\�p��\z�9Y��2��0��Q�w2/����N�3R�C3&�gm������;�n��)%:�AS#���W+�_��`<��d:�������눢��~�:3?-��[��|C��L��b�%�,����>\�q�0#O{���9��W��_��a�������I$�?M�����i�^�j�ڜ��YV�h[i���������j�1V�r���N���@�t����M�y<]KN��T�xg`B��32;��2+���N���	�v�s@N��B1��,��A}/\l eRW5�B�x���v-�^�O_|����8���Ob�) |0}>$��VM�7�J'����N�{�I��]��?��/-Ru8���ߝ��%qшe�u��0������z��o)���(G�[}�q�����Q�rKfG��.v�U�|mbjÎ�O�č}Z�^/���["53���_��t�029��ڞ��{�˳2���V��P�Kiφ%�uY�,���5H�+���;��g���<_骓O��>X��O} �l#ӛ��$tY�U�)%rI�@�;�;�-쐱��,)X/��ApN�D����o'}��1�/�\8���rq��C�M�M&Dp���Ǌ���S����菵D�� ĕ��~(�,!BC(fš֘��<�,���Z"�O&1 �Ε�� ^���Oj�F�@�q���Ԡ�o�f\�!���"���h��UP�A=>�EQ��O^�*犗�3�X���q�ﶜ48��$!�T�k@�P��jC��_�D��D/������ yUi��](hL�����d8��&�b�
���k:�wx�������O���r5<
:�%�de�!t{�F�WDk�`�1�ۋRy�~�?���gF~o�`���-�ذ������LFP��y�ac���1�h�4���㣙Kj�NFhi`����JTQ/`o�6H�n���4����$5B�:����'S
�t��IR�]�O�i妦G������<ۄ�>]����ت���SR��D:�-�q+G�ids���9Γo����D4]���
���RA�gf����9��t�f�z6��X�(��R3���r�u��I`�CT�����=!ſ�ie'JU_>r�Z�6����)?�%�2׺C���,��?�D	ϴ�_�!,��f�R��5ށ�5�����fhŻG�w0���$#�[5���������c�$/Q?�)�_1��&:F��rD�'Zx*Ε���I4�[���r�P��k(��x
�mA�	����y��&���%��k,�v�Ma���~%Y���K���JΤ�9  ��7����C~��,q�D�k�c���;f	@�;����<>�&��	�<�|`�r��b���Z��P(@"��|��[g�M�+����,��V[�ԙJN�|�Qw%&�q}'C�ut�x���?A��$�_1Rꖉ�	�-�Kա6��{�v��1��$e-�sZ
�9�f/_{8'S;��Y����dSK��晉Cg��J�S�pEQ\ſ:��<��CI_������@�&�>�;��������w_F�ow����q���6��l�dҁ�@���f�O�jT����(���v��*|�KH��#�):c{��2�z�3>G)�Љ�� V�Zf�TY��5��i�W��@�c?:V�FT�V�
<��7�C~Ws�hĬq��kpB��l�9���6��������V�w�|lX�e�w�1��U+��$������C�����C��x<��Q�[�E)��[R�� ����*���ɲ�հ඼���o�Ɍ�z�o��b���ot8(�U)����ҭ���ڌ����[�Z��r70M�̀��BZ��s�%շ;[F�#�&|�Wje:����P0*tjR�oeo�۸'=��EgSY8��4�B|�m͏���'J�YD#�ݫ�qA�6�J_�5���~׽��.��|��u{�A��t@az�G��ș��y��XE}����r���aG��VXշ�HxX#qDO��1A��n??��7D��J"Z�^��ߐ�|t;��m�HT5\�n�;��K�n�(�k�y�Ov�A���#c�_*i�tW��������Q��"��O�<:2�R�.h��.�Bc�N9�s<a��,��ӁoZtI�̝rB	c]ඬ���L�� J%1�8ӈ���"��D����pw��$��QJ"İR�kQ}|���'#���,����P�m����'�oi���]�9�6���
�)��3Ǉ���yfk�)�͕-��b,��Is���@�\4a�����n�`���O}d�n�	�m�Ke&$�Fr�ʽD���#}'�U��]�l)�YTa"�]-�4�j=l?hR�� ��qJY���NI�*�Z�V M���֖5fo�i��۝���j�eUfHR��Y����+3=Z�vÑ�8I/�0��@��M
.��Sݛ`8��H2���f|}H�Xe*�U}�ΠJ [��r�ܢǖ ]��x�t�Gz��=)$��:q��k�~c&8}�y����7!vB�aW,1��߆W��6��:�*2�4�����a��N��t�MT:�t$^�Ʃ
 ��f�,�?�Жv����on���p&R��u� d.�!8Qx~Ku 	#&[c�]�$��..�L3�1�]�Ð�Ei�����$#����q�����b�CC9UZf�_�����ż�����C��۱�2��Mr���4���x���n!$
놔�ax�Da	�j\b���cB�Z��l~z�g����k��SU��TiA+])�g3�2U�.�ȁ��g[��#���bI�	c?�J~7M�s�͑%�N�+ヰ#��j ��N��>!����>�����lKj�Y��Mk=#b�G-������y��'�"V�};�	@P��|��2`�[$����v��?a�� �Qk/��'Ou��^��Ӣ��H����� �4�0�	�S�������o���me$	���������0����>�{�=%��w�v��!�k���Ѧ%k*�BJA �<�gm�6� �{�xi/rs+N^�/���ИR���o���ǌqB�GK��n=��G詝H4],�l�l�'��"�|�a�⤄}��"�>P{J[�i�/�7gz�x��:>����EI����s����4��Iލr��=D��u�A֧rY��@�M)���sh�ZQ�H�{�Eћ�f��?�)�Iݡ�4|^%i��V&��Ke�£��I��jO!�Ww?"�}c	8sѷ��ذq2v(=Q�������@Eդ9^%�hny�2s����6�g��-t�EZ�0$Xc(�BU�
�v�{�W�h���P���*��n�Yޝ8�H�dIUhjJR~A��S��Z�I�t�Qx����6t2�#�"��:~�����'��s�Z��8���9�$x5�\Hn�i8��������˜��v'��i����q��"Ce����A(2�~�|�֒�J�-�N�6Ot�t���Q �s4O�$�i�L ]��.�>*�c`����-Y��H���)U�i9�[յ��z�=m���R9�UK1p�����\;��)��o�L_{��EIY��a,�K����I���8���}��}�����J����IҎ�Y[`%4��Ҿ��@���!���w�%&JQ]���O#I�i,qM����Q�#x�0F�S4���	�_�w���؏��8X�����1ͣ��>��@�X�!�\#�r��|�����Έ�>0�į��3�X����sQ��5�<��gb�#�w���,�s��|p�zB�Ε���rK~��
��8f�H��9�V]6 w5٠��%Dd�=0]��Ǯ�Pj]V��<�[�r������%k�B���S������S���R��{ZGȠ��Z:S��|��-�`�>Ou��b&5�]D]O���ȟ�m�C�[�`�>$�H�./�c�7�O����{E��p�l(o�`L���@�{�r����
��	"��8˜�<��ߧX��@9�-���M�S("M++�����B	�ԙ�>���A�v��}�����c�A�턇c'�b8��Al~s�fh�0�x$���d=���$�ƃ;�9X>{�������>7e�nX�(c��ʣ���d߹�f�g�GǛ/���P=B���W&�=����ߕ��.���	�x�{A�c���?���v��+�ن�ZTUG�l�C����ߣS�?���D�ˣTe$u���������R�*
K��� ���"��q�o�'~���v0�C��/�iX�xp��^���7��u��5?O���#�q��M�|��O�����d�"�N܎��Y�`<� �x�k�S�`P�T����@ᒃ�Ň|�S��~o��2�.�9x���y�[~�E�Ң���of�-2���ì(�$vA��[��V��a��(�_W��-��SH����e=�e�I���{?=<�~�X>��Fx����]����C{gT���������4ѺМI�9tuN��HQ�%yV#9�/�7�x�ޑm=M�;>��)�����f�k������!G��W�4ѧcW;̽ܕ�A��d��[F�t��30+��1�R��G�+�)�a�R�{P(�B�>�_Pߨf��%��0&�nyq_��@ū#����g����,V�j�?-V�����dq�Lsc~��oյC��N��i*-�$V�=ˍ�����Ӹ�P�y�?/���s�5k	�!�Ԍ;����e���)e�@n������U�b�����O�g�� ���"�R��*�t�_蚂��n!���N��v����S�"��D�Eǭ�}O#��'�La�O�������s�rG׉[l���q�UҏyO��6�G'R��R~�o�ۯ��`�px*|�t��d���Ե(W���%~�|^J�@} �v���� �RB͞W���	+��Yɣ�1�WQ!���[�>��8&s�O�L���9`���H U�E*�7�(v?:pRaIX�}4�k��s�>30sv|�^�R��5�4�o��[�R�zy	ag">5/I�՗3�WE�^�D��㝊��/�Y�����T�Z�{g� �"�#!&�"@�*��`j(�,a*�+�n�t�b�2��w;�7�é��'������f4ip���&M�����BP&6�������s|
`R�-S���ϙg]{����G���&�#����Ln�N8z��8�}"����u�$���R���ˆ<`��z�D�q�z|#��OQ�3^�Sϩ�P���z���.΍y���9T�����/X�<���~�f���j2��ٰ�>E�I��
��'PU���VV���(�(�P�����A�&DV���,o�\	��F�D� }mF��Sc��'��g���;<�������h�ň�@��T?��K��Lŷ���CxU����[m�Q�j��}n$�hޅ��m��4 Ʈ��o<h��FJa��&�'2c=����zB%�H$�;oPR���r8��G���T�I\D�v���#�`�Sw-�|���v�@b���y�x]�=҄Y���(N�ߙ����������V��G���Ե{U����ۙb7�&?��,)�>�.�\�*�
z���X�����MӖ��D)�U[��Q��! $�.�uw�s��A�������<�mD1j\�9�Ns^�7���K@1 g����1���I��,���)�u%�\��ǸAv��(H&�)P�s�E
�_��#�x��;�(�RK�색��	^�@������Ϙs�l� d̰��}z�c�)=pϏ/[��I���	I�S�_�.b@'�q��P�ps���4��k�.	���ګ��_����zQ����{����'a��f��lC�ë=�S�?���ҀY��J�2Ə��ݶ��r�&ȺȌ�ǻ80W6�Ⱥ�5�H�!�K�����U�u�&����ɍ�ʀ���D�>��wF�[NpR�I�F�d�͓���[� M�>�݊ 
�2q����������K��o�]�"j�7\��'&��z��n�3b yZ#�F�G���z(c���|�O�hC]�Nb��i~Y�MB�-�~K�7i+}�'+�N�.#�VT���f�'"�D�%,	�`rm����W��l!N���S�մVj�@*�|姦�ا>"n����.741uE��/55�4d�/)Zd^�W&��I����w���:�N#c)�>!Z��5�������k���}'Z��?}*4�~�R@n���VC�����gE���?\��6Uh@�w�N�s�կP��>i��5��T�Q�M��r��Tg�n��m*.15�FB�p@s��M�S���7� ��r$��nomj��������'�"4׀�� �Ș�$v{W�?�!&��0x�d/�%\ �NZ�E�Ǥ��#b�_���npS�=#H����]��:j?�Is�J�a���w�z���GV��v��9���6���_E�8�U��$����&(�wR����H���-���T���`�� ��أ.��ʜ�DmN^[9��L��F߲U1T�_]�;X`�c6��Yl���ld�B���!n2ѐb�q82y�Owi���L����,p"T����n��ј�w���AD��a�l~�U�f(Ќ|�|��b&p�)=_-}^z�7��,(�"!��]eֲS�KA�q������S��4���#��,O����z�I|��)��3J�s�����;��
�[��VfIdbq�_��/�]���~�<ـ�t����pC>��#����nB6Ɓ�#Sg�R,�rڞ��7��V��������<$^Lji������h�
<G���~\*K���[cT�}#��]S���靋"��Z�@#�&�"{ܓ�o�$�E�t��z�sf@9�h��P[��	x�����A~H�p<�>�a�Wܥ��F.�#�谏�	��VC�2�5f��F�cϩ<w(E�]���cݨ��]�l �
�Ʋmn����%�FH�m<�$敖���ԛ��h^��I��O���|����91�[����U�:>ky��X�q����o뀰�v���t���L"��N�.ʜ��Ȁ.�Y16�r)�%n�"�f���m�5f��҄�I�*1�0:J��B{���ŵ�=�v���~�=��p�s�<z\u����`�c��w4
�ҷT>>5�����s嬹���`g�=�Cnt:L+|ԿM�;��d��{�?�(4�?���{:Z�����3���[�i�]/9�u�v~s�i�HO�{ؽ��*:<����K��~���q�%T�h�Hb�]M<@䲩Y|1�?��c`nfp�ƙ��zH����d	��X:J�	�,�.�M�#G����MwD 	 *�}C�Z;�՚���0n���{�9�v��j��,r��2HA#��HN���$[�pS];�*�g�* �};t�yy�wCm�K��j-<y��8��%���R�U9=a�� <i�Lt-%?����ӱ�rΆ��
�`�$��#3���r��_>����mU�R��߭#}��F���C��3���O�s��?cL$��5��]������:c'�[ay����@3�u*+���(�8\ǎ�� p����M��m# z��U=����g����o��ϻ�2��+��ف���m+cj�&�|�l�>�|l���v\/ʽoP����p�	��WA�C�<�P�Z1}��P"]�|�.����g�tӪJ����Ӝ�;\Ψ�*ȳ�P��M�	���;�X�*�+��D����vPcԦ+S�0���ԉ�UI�4��c�Z��Yd�ͤ��o� �)����x�?����l�8s�����wk�+?�C���½	GIH"�������^E��>֔��o��p�`<;
�/�����d�.��Fc�F�ػ�7ּ+�c�!Egq���A:'�/2����c��դ.����l���~K���0[Y�}?��t�.e ���k.̌}��W�g>�=��=����G�eg3�m�~U������H�ئ9��}��RhQP3��e|���h��ꘑ��1�!�U6�ق�[ԕ��̓��U�r��0�f���?�m��T\�����*
�� �i7e�/h�����IQE�����$Y=�׬�����n4jg��-��䔘gdb��1<�?�\8L�ڣD�w����Xk�}�i�詗�Q�̈́��~Z�3L�gAO��Į�7@�L��A��8�T�T�ƭ�i�4��8{^Y֡��{5k��[���f�*t��lz'� X՗�3�T�v���I﵇�Y.������g���d+|fp�\��h6�*��AlT�2��F��հ�~D"]��`Hn�ĜY^̒B�3���c��%��A���ْ�ߵ�3=�cX�td4Q��=�O�NR�DڥHzLv����٦o ]�;�O6��ƕ�̳���<H�v��Xޠ���sU�9$_��&V*&?h %�<�}EPӃGc7�J�mD�~G�Q��S����/��k���>]��~�0���P�:�%�E�;*.�yw\7ˮ�!쟱�b̍�pv����1���šH�Jw���ɍH��g꾱*�U�qyg.O���Ũ��q� }���%������ex�{�wӔl������$Ұ�J(l���^�x�����<=sI�#r�w����#�^��Qw�\.�{��zS�F�n�w�|�H�O�y[޿lǵl��^mk`�L�|��:L�lc?��Ԯ0��gMJ�	N�a�M�6���QqW9"��k��$�+@��bj�=	��#[U�lQ})��h�-�LEF����P��9e��r9�h�z����>�zCF��b���p@��Kŀ� 
�c�~<z�!��[�"�SX@k(�X���c�Z��K�y�ȕ>m�;ٝi�B����M��1�ugQg@ӱ��7"5/஻���F:|�ӏ M�F2aJ���B�ɚ�/y�� ��5^<�����b.��{��k��N�.���X���7����
e@���=�/A�Lw��g�9�+~���*�BtD´P-�����*'�p�ӴaEd!�F�����ھK6:�����ތ~~�|JR��0�q$�*1tSO�X��t#f�Z��D	V!��R*���7?Ɠ��n�(�<�+7����m!�eefp��FfN(�*[���G�m͎M$A�1 �����=Ӗm�t��ƺ���$OS��#,�
��ʹԓ΃�N��F���ݚ�qCT���n��(1�������4���d�\��&��ir����R 0>�"�S�W��}����H�����E��Es�� �_���{'2�P�h����\#'�@��k"����$N��٬���XY4>�S���#14)�0�ri��;W:WO�q�La-��3�\z@�(���F�/+�����mo�d��'��</�)��v�ZS�|��`�&�-&�fOYu�Eg7�����dLhq���ۚH�F���-vs�<м�����r�P���?ړ)W!Z3^��H3��}g�;YЩ��r�����*2f�����l,(8�Kd�D�h�8���1u)�M1E9�X(�Va���|L#�B��?�[�6z]�&�� 쓰�������.�p�Mx���<Z�I6�
���r����;,��~�U�m���̷��G��4�?و�~,�4�-tP~�קQ'��\z Q�n2�ܝ��v��AT��P�����x���\S��bd6`�v�:�d�	�={j��ʒD��ڎNVRr�:��U��"�Y���Q(���=�����G^;G����(���d���5��h������i�ҙ��q��8�N�O}'+#/�8��SϹ!;������ܸ?$��q�V^}����f4މ؎D=���v	n���L!-�?���@�%Xd��`�Q���l��5%�TY��6�"�E(�1�����,�*f=�2_�?��$~�(5p9(CO-٠Ś"�s��	o�a��2�c;�]�%��o�Z-g���22ƑP�v �ش�ޟ��
���K�˪hdn.����ɮ+��h�S�\x�VOL��3�H��:($S ��9b��)x��6�
�Zϧ�juJc��RD7���ҵ�S� ���;?�=�����`�X2�`d�����N���>n�>�ZZ��MıK0hղz{aScRL*7!〵5�κ���n�qv0���gީhՔeK���0��c�~2N�Qȏ�\���ǉe(�=tD���1�_�d�FtMW$[;���+��z�I�r��D[d����&q�n�D&/�S=<�#~�!�y�O����qf�ߖ��*�ݠ@��&s��1-r-�ٶ�����	p7�;"�F������NMa�F1Yi����?�����o�L{� rASjC�q��p1���O��v�dwq_�t�Xr�@oeD䖴��y�ab�Umh+�wWs@���D��Ab
�]I$aAiװa�ȟ�d�����^���o�D�tx.Aq� �"��tGP�	��ht��`iw�J���Kb"~Ny����i׽�R G벭�`�w5�7D����\�Zr��J�T����x��ck�1wݧ�����A�����lN�0D���	7��͵kڕ��0*�K^���m(�k�Ý̎�*���r^$
���_�z�+��St�AUZ *��z�