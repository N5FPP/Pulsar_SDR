��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,G��U�	�oJZ�@�z�����>*Q�p��~!}8~��m��sDmN��3\��\�A,��y��,�y'Zs9|�v�G��Z��J;���������!�p}v|)�pB#1�F�hZW+	��M�����^ ��RK��d��$��BB�a�����*(�y󵘔�IYS�0�"8��M�px�	�'k��}2����p�Qc����t���[H�(���H�^�X��"v�v��L�p�Qd�ci��H�z%K�t��	R�Ͱ���1�&�� N�%�ju;�.�b�LO������!l�KWȐ5=� +C#Z^~*���J�J��r��c��B����l�<�޴_o^�`�`����^U+Л/B�t`�&����:Ȩ�'&i�EӅ+e�j�Y� �e��R�Y�h]d���,֡&S�|&�*�J	��A�L����3��w�=��<J -���}R53���R���@���ܔR۝�<�X�����~��e\����n���آ�rr��}s��""�ʬ5��s=��ƒ����gc|��0,'�d�L+N����=��Ik-"�x��&`�?���%4�H��׌,.:�Se��	����%�)�E���@"ɹ&��]�CB���dB"c��_Τ�Ȟ�rr��[�Ac����}{5�7R�{<1e��A	pfqF�^���L#�NT�� ��v��?�l�YH,iQ���_���m*{�nɉ��tKi��\��'���d���g�
Ϛr3NA���Ϛ�A�nN�'ŕ[�;���mF��}X��q�	�8X��*�����3YE�:�X��%@�����%�8oTx����=��O"�G ���I����|��L�3Ϟ���&��ZA�,�_p,L��dA���eJ�����ċ�a�Kj� !<�hzn��O��|?��OV"�.���5]8- �|��Qe����m6R
�����Me��
F=Йr���]��_e�B�Վ!��n0>�	�b���\.W��Je-$���o���吢��ʃ�'Eҳ�<	h��U)שhi8�Fz�06�D5�?��I;����j�V�{�����YH��*7N�+k���(�y"(���SsD��Ζ�:�_�(7�:��܊�c���SeO9����G��#E͊�ԋ6��W<G�D�H�}��6��%�5*ͤ��n�߳�C��G���h|3]��
�����2��e��a���R���UmVy+R�0�j�.���"hw�PovͿG(���A��.4���k
�,q� �Că>�5f�%�\��eN�kC7�?��E�D��^��Ji-��`�1�������dź2T�zj/y�sP�u5�N^�UE-T	�^��6#V��\R���`��i ��C��#}��kEn���X����{6�(ӵ�����$P�/�����3CI(-k����U,�r��z?�A�aE���C(�`���曾_���/ŕ��ܒ��B��?'A1����H��]*$	��x�a8c.KD���s5������������i���ېd��ZePЀO
r1^Z� �wЁӞ�br��Ls���|i�C������]j�1�P�o��@�ͯ���cj܁�:3Ӕ�VH/��J��2}����&�g��8�C��,�:��Npn��M�Ȟ�S��4�.[��+6��x����m"R���Ė�����t~����L�3�w?$t�"�[Mv�C�L�it���$g�S��3 �x��J7�"��]����ok �R��f�?��F@�i%U��bQ�ٵ�`����^@p;ڞU}I��[����?���1�I��ARو	>gFL��0-0�wt��9���d�-y���'���|R��<��<�z�U���w!�d���O�F�6H��V����P^+yhQb��Ek�o��s�2��*��ŗ;m��|���n��1�qSy=G}���X߸|� ����.	�+��(i&�������숱�|ԇ��b�ĺ�~���)E�Fq{+2���Y�%�x��vp*!e�q�u�8�C����\=l�`�o��{�L��X�;ߐ�h*<�rt���RJ5�qie����A=k���.�����^Gq�~Y��=�9�;IV��z���-���r"��6n���V�R5�:����wTe8�A��"��P��2x�j'ퟠ�����O��t���@��\6oUw����ͱ��)��}&����wٿ�\j=c$��cBC������]��*u/�G��> ��k�&�,#\�m',��^D���(٨5�9șn�k��;�b�9�;t�\�6��K_��N�`AX�����E���@�12�]��vQ�s`G�O��*g|�i�?�R�:���#}؞4r�2���&�[�S�6r�q��ّxp[�D^�wf��\z���ִ�V����e)�>E��Κ��K�bs�*�Q߂G6��=޿z�E���w��ˤ�9Xg�-y��wf�"Ws3F�"�E���W2^.L�)�:z{yh����� �����^4�4�O4U��$2 �M����v�]-mPCM|���A��%A�}���b�;{ �%b��¶�E[�!fFL��c>�˼T0{�j׼1Fs����SL4��jY�l �Ȧ��h��3�F����lP�Ct�*e�&2M�2LL�b�a� ������)m]l�{"�gҏ���N ��ցm���E�/�B����J E��^� VR�fZ�X�)��@m�gf:;	"'�X|��`��
oV����[;]�ƶ�A�N"���~�ߺ��x�E ��ꩍ�G4���V|�Vx�2J����H�rd��@��g��;��]���w��Ӑ{�)�W�\	���A-�F�=���}��1�М<�IpuH��H���G�C3�B��\�K��e��uOPf�V����:+���Pֹ�_��#�U<�ܗ��Y�3ngF�{M'ڂ��Dv ��6!��pA9�g4nGD��FCő|�=b'z
���TJ�s�?�P$�>�ztS#��dLرb�@-�%T�2�EM��R�q�0y�s�� �|8]4��;��?1mj��^67�#>�4�=o�`��"y��#;���^X]q��᰿g�®�Ѝ�Lu9į��Z6?�Y.����YwX�y���Ӳt�d�'���X䅵��Q)R8x+�Iآ��9<����|�U݄{$��b,�^�����L���`�p���pDe�Z讁^�2X�i�"�� ׌�DP�Z��a�2	���FZ>���7�=�!eh.n�oNz����6����R2�=]TL��A���'G�!��)�� ��v)��K�Yoeĸi�K��k��<�GG{^���&��9���F{� ��<��N#�!\��w�NM��!Q��H����i��p��H�EcD�#�l�T_�Ȼ����O�!�_�ڳ�⵵�y*�H]�9��.�>n>Rp!1S��=~�gt�i�)q�vp0��[��0@�
O���T�E�dk\X=
��w�L(�:l�5�>����,�&FPte�T� �pe�Y�T��fv�)�\#�?mk�<� �����}��)g���:��Ԫ�!�J����n���l�r�ّTJ�_�e? y������Z�ex��FG�ڤ�/@�MLk��:}��Ҿ��,���[�/��<���n4Mow9�-.һ�.(J���5vp����Ǔ��-ys��7�-Y��(��'���i� I�!r��|�ۥÜŝQ�ز-o����%�"�Mub��	V�'T�?A��,^^�Vìr��ǳ
���q������	]�X�1��X="o��:,ߧ�6�R�@xA�5Ņ�POc�IJ�D䭪���-��t��$�m|�W����	ܳ�7ۗu����{ō�]<B?�ԘOg��oV���:E_�9��TV=l��}$���&�Ԋ�ϊ�H�1��D�DT'�7Q@���N8sX�Hba�=*�H�D��k�~�������®��Ն����ꋵU�h��\�9P�J~�1=a</��SHKDq�����9z:��\H� .9���\��r߳YK�BZ�8G����!�(�)cqG���|8=��t'�I��I�9�Z~�afD�ֿ�׳9�?�]��Ka�l�F#��6����=���}���(m��@�)k���3����rq}Z�g��Uee�]�5��o���8�y�D�����n���x�)��!��z�֔A=��B�.'%��f7y7�M�$g�Ʋ�{��u�iTa�	能��O>"m2o��0�A�nȬ$�p�"� �mi���I�vGĞ�T��>�}&ylޖJ)4�I�|u�|�&����p��C{��vx�I��/�<�s�_���݀�eJȯ�4�m/xX\�u��8��kx�)T����>Һ���ƍ. ����� >N�����UA��^҅��: ��[���Y� K�Ñ^-��>v�0��0e���yml[�>��)�\bA��� ��0!\d{��!����ǽ0��!���摔O2V����p� ��]�3���a��nF�D#�����+)��7�T^�>Y�Y���!)i@h�L�+8����5��#�p�S��{��s7C�.�8F�>$��?�}i��᠃�_����[�š80�	2����N�q��*��R"�\?�4�%,�s�t��{��X�F��iͳ_m�Ǭw:0ǽvFK1��uǤ ��ٮ��7῔>��'0�����*͘�9C�}�$#Eҁ���T4t�u����\�]%��]�kj����6z��l�Rݠ46acq4���oe�
���W�B���4/)Qw1�Z�!B���^���d$�>b�̈́��7�ە�KDT��I \�U_B����]�UVv�M��M�a�"y+�L���/7���Me>�V>{����ߕ��A� �-��=�����w��.����II�${��X��;:H�B .,05����I�N���&�:Mi7�7Z�)|^�6�YZqN����~�T~���I�.BC	�̀	� �jUW�L���p�]�kEQ�n�jL����7��ߺ��1�⥒����6Km�=��36%�Ē�~U��+�H������B>/K��B�4�*�eWz��7ՂN�,��&����D�d�d��ٷtb�_n�7e>�~�X��a��4�ϴ�����%�G쁰�f�V�5�0���,0n���p&Õd)n	�������F�ȍL��ty������̳J_+uiI��Y�L�9�"n�"�lK()n����[mL}�H[g��)�ǌ���g|��������!k��u(f��j-��*nX�L�8�6�ڸb�Qq/�yf�
���a0c��I-��k돐aʙ��%��:�WԪ������cdtD��Y��u��"xn[X�ݵ��|��.R�g:�e�����mp�cYL�E~�ޖpw��ti�u��y�*�� �������wO���!�/Q��ON�=/���&�y�N�k~P��{.��c�R�g���,�6���u�3p�9�N5��M�b��u��5>�68�-<�n�Vi�+bm�
���b� 6rBV��������:��j�3�qaӧ���]8GL�ԁ�,�p]^���~��_f^L]=2