��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY����ﻅ�#����f�D�&*����}ׂ<XC�dZ�p�6�6��nX�������q�N�8tjǻ����wAr��!<�3��i6k�|-/���8���$ak�r�L����yr����#�t[]�+��X��:��'@F�^	 �Qٷ`�X�
�e<���>9�����~���.i�ŉ������<^�g�}��۰P&_|0�����k�'u!p�r^��D�ح��'J_K���f�Q`�b���4����K�}�;�V��^9��Y5Tsx��n ��O���yߜ�j��xo�<�8֔����0�gf������5ŕz��X%c��#���
����$��.����&�P[���c �g!�H�|��{�\ӱ��i'.���BƘU�=���|���\�����)��~n%�a�_������̝�p���2���"s�,�9
\�CX�qn�40�D�x&fL;�7;��P��w─w^��RiGeĠ�nb�l�����Pmmo?����k5�r�����3�V�S5l�p��&|ӂ��Sx�F��� apj�:��?��˦Um�ԀGw{G�Vl���G���2�M�fxaB�� 9��".�X,���<̀��2T���v�>�����<�C���@t� ��HL�zu�D(��B;G����8���q7��h��<	����k;��Z�5q���R�!H}�_{���KTHp���\��꾤�ݬ\��M� )OF� A,㚃�����~����+FD�.�����8�q0��X��f�`��h�V��:�UdY&[�n�ょ��{��yL��:d4G�&&��61C	`��P�w�����S���my0<����{�-4����Z�m��(G��C���s��%�*��e�\�pk6"�/*.$�kʹ��tÅ0SgjK$C	�+2���6PNъ���%�
�G�K��g�����@����)R��k��j��xlH����w��ϖ�@�@�9�l%|Q����("�Ȥs��#�m.�� +G�J�JW���t�!ŧ�)�9�
�ע�,H�`�~�D>�kU��OǊP�}�
�E�OF��l3�[w�7��j	\��`��vU��@���ޑkO����F�5��	n>I�U�EIx����@�:��t�q1�
��y[xG����g���\+ʛ�URޣ��h�<[fP<l�a[Wu,�y��<�=Љj���װ?9�oڒ����:�K�1���d� �TZ3m�z��gG� I7 T
���b"uu��}6N4� �0b6�H>�xD�4 ��ڥ���г��4��rR@�S��U�3��e?;��78�����=)��v�3#c
bٕ�e��,.Drn�;��	��#�=m��
CL��f�d�ٌ��͎ /,��dd��v?�חF���m��.gW��z�C��(��A��Y�_�4�F�4���E��w���� D��1k⫑VOGUi��A��8����b<�hVb�W(��m�/`\���HZ:�,k����a��yݾ��hJǚM$2Q\'��f�Ě��(56�����-��3�aA�ⰿ�Ϛ8��ҫ���y@*yG����ao1�5�r��WȟI3�,m>̋J�o�72Y@Q�(�_=q❸��jh#ʲ���9��Q	�5J�$
�A*���_�\vɾ��R���C8�g�		$8ݚovom�K�Q�۫q��En�Z�(g�⨥`�o"�:[$;���loN煶�YAߕ�`����X�h��r�1�%���5�.g�3�y�v{tk�[G��ط��$G�T�R^J69��#� B�dߐ�d��_����������o��#p��1�҂/��(Y��êall����qQ�2s�� u�܆r8�=+䆝٧a��/G�H+��iX��^cd��hw���9Bx�e�^T���Sa+������ӿB5��tZ� ������|Irf:���I��e<��ΌS�Z�+�*l��r�|}�0�@~_O��_Qr(�T��LHl��̤��d�I�0�٬�!�n"`��|�r�s�+/_�@���{/�5�$�6�����m��x�g�d6	�/K�����/��_�]�����E�V�ko�ƕ�9��P�)�*%"ȗ�
 Мk�z�G�r$<'�� >�9�۾�&0�g5V({B8����4i��M��^~�CX����B����1S��@��}�G�b��6�c����$C��7�Uw�'��&���@}�-ꍘ.��#��׏��=�ͧy���/v��qT���`W���<���ǌ	�N��\|�sRǰAEx����	�륗���I���3��]ԕ>ZiP�i�y'Y���+�Z0b3����KrW���e|T,`P��@��R!L�42L��]7i��sDnH�I����GY6T���86;��$8$ѿ�lKRO��~����d>�7@"@�xØ�i�VC�~ҽ0Ż\�g�?~�����#L5�h)���zF���Y��Ŗ^�
_!,ي��o��K�Y����/�2T'FG�:7�G��\r1�m�u v�G�ɱHG>��'n���׽LF��i��t%����i2/�6IԸP?>��+^�DigƷBx4-�#����D\�������]l��]��w[j�xb��e��|3���f ��w�=�ZJVt����;yD��E+Ŧ�')?�� �����Q���6]�2�p�ʲ��j����Z�fj3}G����qP���>_&*����+�3m@	2N2Ű<��#,!�0����@�Q�ƠcT������c� �~�Q��/5��վ$�n>�7���Xnz��q�P=�˜8�O���c������>��r�ؠ�u��s���oJ�|�&�V�n2�xo7)I�-y����?�C����5Ğ�߼w�4._
@�b����v=�~0�hifz +�*�������6m�����O���57�bP�Q�<lX/`�ZwY��m�O�&�ם_m��~`�u�v�!F�y�g�"�M$R�{���GQ)�� '[�����:��¦��ס3�Y�Uݬ~L�
���Y�[RT�;��^]�%�]^�
�P �aY��*C���>��6�՛����������
�8Hw�	$ܦ��⮒pE��њ/5weWY��٠�F5�3:�����U;ߦ�9�7���׾'�mp���n$��յpz[�g���z�3�I��!3�og�xIZg׈uz�"�B��x�E�9�X@ؗpx_[!��r��cI�&��l	Zø2�ɺ��T"�¦�(�b���;�]���pN�&O�(��΀��6���p��A����N5�6� ��6�y6�w-��Ls�v�O6[Ke��I�������[9܌!S���_
�!ERq拏�O�t�8��񸌹Sk���B)@���a���[de�CJu�3�uFn�UcH<�8�L-A]��sWgC(�\#�N�x��j�ʊVnXl�g��Zl~G��� W�"򳱻P��нY�%@�#��'R�n�߯�{�AfwngB
����}?�3��4QO�3␾�z����6�+�5Lz�*�ힹ
�Kb�B�RrfN�$�JF�`w_u[��~�v	�M��]�_n����I7�� �;$������Ĭ�E>; ��OR�	��u������U�D����:��1��TS�g�<U���\ԡ�]����ݾ�e����.��}��[�K��q�����ϝ�ذ����Y��(@��/���$A6OO������x�Hvr�����kW�l��ڰx���~2.jAհ���CeE�{;[7;������a��٠Kk�`f	�d Z�~fk_O��]��NF���X �v�n�C^�G�'Z6?����͡����x�$[�?���-�g�[���������SR-_����Yo!�VIK�z|�q�Ι�G�^P��������6�����k 
�|pb�,��)�d7~�;2=s���Q�аh�Mt�	�l?|m6��`�5�m<4����=��.���?X�F���tsQ|��z�9��Q=V�z�w�b���<:)ޢO��/��|G~�]��Ǿ�:�c��*da0�K�K�#����̀�AǞH9�ڔ�x�PI��t����Id%Ul�4U��n*�N9�#_ܵtB�
�Qh�m���SH	k�7��q`f$yl�����C�+W(���ں���,����n�[E�N���`Xc)��&ͧ���f:�Ԗ����hn�Ln��Z3�'@�/p�.��J,uW#�G?G|,�D+���~����>��QCe�����D�4y�Q��Uɒl�s�74W&t]�C�Eŝ�i^�ЌM�����m�*/��把��C��1t��F��N W b GtJ[ƣ�Ч̑Ι���rQzZ��/�lB��K�'��B�O�8��?S��"���-���J���̮�uͭEm}�v�����A��S1���Һ���%�	��)L�k�9����Np�汜����.&��I5�x@æjr7�_��S[ҿ�#��H��Dt<*9�rjO���Oe<��^,��A����[�Fs���'�=!���y���C��|o�;�?�0g���������0�E�۴7+���d�.Q�s%C��Ϟ�w�y�f]�^������`[bS��;���@��K�9\� YL���4�����ڿt�]|�<��pT>���g0�TK����
;�ʍ�k�����1��s���P��~��$��-�=�g���\���p����^���,���N�Rd��������*3�C�!�*�Qs��P�{����UlaF
���{�I��
�g2p�v�X<�ݕ����e���Ii��R��LSU|�`�|wГ���X�g�*[N�_�n{1�©Aa�}�/-�4ݭ!3����rNL�G��~�;[�ܖyk��?rg��.�s�z�e���"�mn�H�W�b- �P��E�\��S}n;w��B����fӥ�7%AO��Ӹj���ocn��}��
�~.���ΉJ<=�_� Zz}��˻�֮���Ο4��͚{UL�����%T�Z�"�il��UK4���vD�(ϲ�r�y�7#m�t�su?�vE��(ٔ������JV~��'��D�{�hȉ����Q��=�1J+7�n(�Vx}����RxLo=�2�C{�G�w�t��*a�Z��ȳ�t��k�=���ƞ�a�ו��.�lq�������A�pLn4�O�j�ȃ�R>#�6���+����� �����$��>�P@��ʒ<.�9guG+�4��9Dh��P7Lu;�2ɐ��t�0d�2I��{�CD�U��a�y}z�?��),zS�ߦ�	H2e��і�����7�!��rj���mz�iB$���Y#XT�6���歸���P�V�-�#�c��%�i=p��:��U���k�||�I�ȈIzr.\��G_̱�o:���7
��77q��,-36��n�G#P�@���MU�i�jS�^�$@>B�C�X��l-�JZw�=�=~.Gq�P�4�`���+%,��vGЙ5*�+dzs��`�X��S"�c��uyk2p���U��h���)���ɒ�%_"}�&��L�/�l�x�{��C� 2L��ƽ�B��=`$ݯ�g��K���!o����bc8��j��P�0)<+�rrz)%Knl�ġ�2����f�駽�^^�0)�� #)�bv��"�/19�Z��8�@
��S�6��i���?8N4u;@�,��K�A6�7gA-�_���c���Oo4�?�.뒙�8��H�H�.U9�wM�4%��L���d�gt��V�r��7�h	�Ѯs�9ҧse����/Β>#��΍�$�����?\d�ʝ�	w�w��FɩnA��d���&��5�xP}h����?�v��@���):R�{J����1]��߂hd��S4"x��Ws[��^������]����O�Q$[�ϩ ��0�M�s����ǦR�A��z��D-��[��>��A�Cm��u��R��'� �L�@����u�ލ�^bC.E�.~0Y�V=S��v��מ.D��=d�7�����m�!^h�@��MT�=��e�p���eįQ��(C	�ʈ���7�OvŰ�h��(v��
藇"Ǆ	c�-�,�9��u����SЏ�C9^QKy���6=���<nj��3�Y�%y��.@yՀ�b]1��� �rXf�TT��SpB P��"��1���y�Lᚐl���V�r,�P��R�"{��#2(�[�R�cv�- ���`�LǮ�R-�L��٧^��?�88�� ��k���)i��Y�@Ԃ	r=�ea0�9�H���b
���h��{�y�6�������a�b��zf.��a-�(G�R\�T��L�p:W��xeO@���J�-�~]�g���|y������$����l�w�𽩌���7�լ��Y3��Q������4���L��"�2�`�w����#���fN!`�)�,��ؕ6��kω��9+�+|�0�B[cP󞯭A��a��gji� ��V>�g�wvu����q��[[�u�A��N�g�Ɯ#��k.��tcV%��P�r�mga�@��gwN�BF�Q�t�9����ɝ��}�<�}wމCR�tFԔ<z�~nt�9��� I�U��r߾��W��+�+tK���ǂ�IUw�8I��>#���q�,?I����q�c.�ϦO7m����$�������T�,�aq��2�"�؅�C���(�a;pQܷk��岞���6�?B%�r��b)���W��{��ӑ/�k��s�f+M��(o�}�E	��3b�#�*�����T��J������Q�{��I��
���*%7݉'�'��)�m�.�q7�Z;�5k!�Qs�8��r˰J�L��S�/�E�TB��J�>�i�~���XI̘�v���-�Sa�����Xt��z^�Nm�_T��*���_ӕ��\�\-g	��"�9!��I���������䨘�E`��_z�9�������@c��Fi�eQ>��#�r��=���v
�����q�[�Vh)"h0�S��2��:݋���c|��>G_��0O}����D�0�=�`mѠ��X��#�iD۷k��c���}�m�R	�ҽ�����ƹYc�z�I�sa�-v����b�Y��E��Jv�]�H��T�Kr ���l6M�3��z��c5	�%�dx����(���+n�}`�WᔾZU����@�ҳI�>�<=�y�E=\��(�'�8a�'��7L'3���^
��!�C���ɕi�tՁNG�����uxh(C��_�m��ٖ+Qzp���A�ҙ�T��V�M��X}�T��|�����lOn3�#�#7#��Oӏe�[�n(E#�����"L�{chK�E@�����A��!�����#(2	Ħ�u ��E�tZ�� W���W��C7�$�����)�Gq{N6ʀ<')�q�����s�������Sɝ�FƼ����陠���XlG蜵����s8���[��F�z�<`$��+���#���Ƞy/$�d�&Sv͖'��"����
� �p7��C��L؜_ l� m����iP�̱��k�]be�����XP�z�Øi|l���bB`.�|�7{ݫ;�ś���&��؄��u��U��֏$��7���^3Dc���Υ�O�׃��[���].�����:��=���KJ���y��",�)��djr3�N��yݒ��i�u���F���O�}��ׇA(�έ��h��"��+�T*m��8�a���[AU��X�R�B�E���Nn�E��h+�pa$H5�I��F�ͧ�t��G�	�>�+�n��
6.%q[��x)!!�'��m�ŊТ�C�^Wu&W�5c�������՗� ��Rdpd�7q��T� �!�@�Tu|��Do��_眛R+�?D��{��[
����D���a����)���έ���˥8Ft�+V���H�A\s���ULӤ�Zk��aO�N��&���z�M��u6m��	�/8:#ya���"��8��H+�h"b�QF8aT:�����4���\�R1{��w�L �c�L��j��+ɤ��p���_>�Q7��\��.�Sw���|�FMf����_�,}Z`��	L�e1[S�5��5�
٭��nɱСuy6}4�ܰ�ryv���7�o�%��)��l E�h���H���+�v"�S޷�0ݾ��!Jo��ނ;��&�&���X`9��#�ƅ��O0c�x\%c�|n�{��u�-�E#F��|��S��ZN��q�К"�
��T촹'f��7#�@����!�[�%@�����/�9��R�Ӊ�GZj�L�RF�͟1��ˁ�.�Ɔ�s��T�3��B�-���V��'���Ɏ��	�%��ɷ"�fϝCC���%	����0�ypY}���yFP���Y鏺5c�>�H��;kc�TS���d��ɖ\6�<E�ٶ�N���w�0n ��11*�-�[܅^i�O��V5��H_�f4/k8��Q�_��>}<XM��Y���v=AA���jy%� M��^�����hlF7�R��hxZ6KV�"�d7���s��a���"+��>�C��w��^�N��j�[0U�+��$t|q���,)���眽�Z�ջ}��qҹ��eG����&�]�1RW˟L:
�N23�LJl
[=�C�F�4Ch���#v^Yi'A�hr���K��](e�_��yu� wް��)�<�Ez!Z bM#�
F���+��?��_,b9!J����×p�`*���z^`zI��"�����:Wo���ju���n#�B�1R�{�n�J�ƅ�6�oF�^�>=2sݷ��.�sD\��h���{`ĉ9AC�o7��&�
ϴ��I�������3��m�/Pt7���<�V�@�YO�'���K��`ض�S���)�1�����=����{辝?���(�J����>�:o�>E8