��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�����"WYj����i� �N�7A!�@<e�]N��?�jj�����W���a�q���#����MP�F�pdoF.8��+:���h1�ԭL��L��[j�1���߀/AP�0,r�F��x�N��>�RziB�M�\�P�ua��B�MɥBe�U�����v��+�R��|BC�:6u��8�B�����趟���*���I�lklry�.T����b��`m��O���r�k-
��P�&��3�����vF�w��X���1���Pr�򮰵Vl'��9�D�j��g�Ǚ�ѧ�|�	)����uZ���(ƶ�_��Ę�-yݼ�ܗ	l�u% ��h�ʦ��Syp�Q�K���쉗3f�Ɏ �Ĳ���]��j;����G�%�l_-I���0����O�FC����T����p�؏8�/�J�+��(�'�Py"cYd�b�{�ޅ�솜8]��յ�5�BL	PTT��<U	Tqt����|(ʘ7Q4��Y�L	{7`�VҴ�����r8��]�Hl)�����u"�<i�_�$N@!�v�}#��<C仙�;�A��d �Z_�
/ieR`�>��`.#�k�¦ "�~a�U�$9Iѥ���(1��67PH7/��sݰ;|�T_~�d�>�- oçIm-f˝�*�D�b#����vjR5-7%Е��'�d�j��dgѬ��RK�,�t��g	�ȫ�jp73�,]ޖ.��V"\ttw8���c\*.��$��c��x�f��M�i�04���w
hZ8V�'�)=BXbθ������Li�]c�Ѝ+�_�A������kp�LW,v�3����. ��`�Ɲ` #�BnF�n��4�(n5v��m��,O7F���:�T%�(����Q�H�WƄ�n��?������q��`�ss\n���V�]�|�,)�ŉ�]��ox�W@�:�n5P�Mֻ��o��q�� �;�3�p�㪋��9ʬd|Ό(&H(�{���=p��;܆ �~�ݒ�ko�K�e|���.H�oL8��y��baWX^)�(���
�1�V�ްH,>�4��v�V̳�Y@�u#���vk�YR6� eL��3����'<c�ոI�l0x=!�S��E]���]�(� 
��O;_.�=⇤�E쨨�#�5l�N!�kr�T���`1���/e׮OYO��4	@�D��"�Bj3"׋Y/BȂ��� g�d�p��Rvh=O���QL���9��,>o����n���pkyY�oy㛴�@�N�.��j%j�9�-�R�*ծInP��]�W�n/@�'�f����H�UO���:�.HU�i�rz�O����Ę�26���Hx�zo��urz���S;k�ugY��#X�:��u�6��!���JTړI$'2M�ȿy4�R�>�m�KOT�S4���H]>�c��!�Pr`2<�I�D�܂���=	�/�?;�s��ao�d)��+'��Ԅ�A��nv
cIŝE�k���1TiCg��63�H57v<�\þ��G��B���)�1_����O��!��=e�>���؝�QG񥒛I㒻��޿��,OhY]%.�@�޸�C������m�w�E��h�^��d�U�}m�˹�7ܬ���#S� ��:���*�[��i�SlsD�qN���׬&ܨ����]1d���[��
8��Ce�ޠ��6��ꑜ�q�}SkZ! �[ L�j��Y.��c��8��y�,�q]�1�Ю�@� Лk>���7����௟��Ơ�<�麂�<v8@���������}�,{�>��z��J'�Z���o2��Տ���� <�v�ڱ>(�@�%��3V;�0�`��yϡ�ۂӱ�Z~�{�X����Q&���L'�)�r��#�Q�9	#�uj��)7m��ggX�I[�[Q^?�|��UI����6�/4�=���s�_�e#��x�k��r}܎�dL���q���0���;�Qa�����3�P�xÐ�%ܚ�ˋ�j��R��\�:t��9D��(��)�캞D?��٧��-�"9��d�xK-�%@͎q#��F���L�>��$h:�b1;泄(^�_@�I�t�3m�a���ˤ�%9�4�)F������J1 �հfeS�vY
 ��B�L����v�ʿve����&�f���Fҵ@V'Ѥ\�������#�� JP�w������I��� ���n?O�y�;����Ⱥ�@������6�OR1�	������)T�j��Z+~�k���;页�Q�Ϧ0�+�X�ZWeZ<s��lF��WE�(��e��9��t�3(��.�ofI@lc�=,�U?�W��(�c=�l���I�n�L�)�F�����X��Lcpub�ۮP���R�ȏ_Ɏ�hM�I5�o��Uc�{L�} �{�Aw�Dhd��+ ];ぞX��1D�_�:ZC�G��S'�tǡ�("ክ�0��T�ԩ ���D��\����ߐJ��ı�Z�Ѫk���̟����Mi��DAZ�x�k�a>��=;�l� K����u]əf9đ�e��ų-:p}j0��]�U��(�	̓V�ſ���iwvA�����L�K��~M`�EfB���Ԍ��D?ܫ�n�n��S&��gQYgC��ݟ@���Z�5���̏$;c'��X�S�
�(3�ȼb2ed�����L��dWg�p�&a��� d�+S�P�,��ĤFi���8��B_�$�^����1�/��R��G$#ƾ:hxTE�J}'ݸV��F�Y)u�m����)��o>O2��/)�S<W �ne�{9��A���]'��}�q����Íܐ W]~-�;h*��%o�;���<t,>���k8H@�y���j�s������g���2b�[��6j}���Cx�I�{O E��/@� 뉔oǀ�]۰o��f�vu���,�gdFIխ�e�����L��G��(uOfS/�[C$Y����}_&͒�W4�vA���+�S�v �k{@�"b�YS1z�Y�g]��~D�ƴ�$%d��(w��6�}]���N�������Ҥ�\"�P؈���Z*݊_6[��lvƭ�����Z��0W�Po�O��1��4�UC��ٚ^	|bbʸ���s���e�&`D9�_�@\d�W$DD�c�`��Uݚ@�_{+:k�?ES�g��#:�%p���0F�y�s���%�[�E�rф?ǟ`���EyE�}o���4v#56/����XSEQ� �vW�n���g�)Lr����W�}�%1�̧�l�J�����I$�9�D��6s���]��h����s�:��u��K�Bu)L�D����Ld�M=ٯq�	�X��W��zF+)����3��C�"U�*����"�a�%�����G��5����|�@8�ԥ�1��t��N�!�5P�%L��fu�Ԝ-\�q	�1���L�8���l�J��g���%T������$�u$�ټ�f�Q�;��OXdN!�j���N{	����57��1���X#�Lm�Y9j!gçnN�:z�PZ:ݏYaӡ;�~�&zq�(	��ޮ�h�5&fDf?�@���0��ԬK^+�ӆ5r'J}a�ʅ��x�0�b�UY�!O�g�R�gm�e�2k���v7�1�6LV��7"�h�:��t.e�:�)�JZ[���fU`�G҃+kz�9`G�EA ���J��D
�i���7pW�K��nZR���4���UD��fV�=ܧ04��R�/8���*�]݋,;�8P��݀�C$�7/�qG�OT&k%�i�pM��+��l�64*+]����l��1r�x~g3�+Bb#�?z�2���NC����y���&-�����u	pԎ�g|n��^|�wے�6�y�z����u��π����UүAV3[��|C�3'UO�>�������y2'�<�.'�/R<I�J?R���N�xD ��&qii��x5�� �-�km�h��i-�cS{��m�ב������/�C`�(�.�z�q�c��XWwip	轢���>�;Q�����ξ��{p��T�J��Zg��0Ml-��$w�Z����$=v<��1���{7�81���T������e�~��C���Ъ𗈅������E�� c�
��[w��#�$��+��7�a��'N���#.ԓVp����x���2
l�ci
��D�WGu&kbX�r��ر���K#*6k�k��Un�(O�Y�|p�Ӹ��(G��F�Z�҆����'jI��`���11EZO2�_^�sN�c�|�JY� ����Z(Ǣݥ����iO�<J�z�س� �(:W�;��>aR:w�w:����i֝���}�/x8���仓=��%�i0h�6y��ԫ���I�Jԩ�P�
�N���:�n�+%7-���7����;�C��Ը�/3���/OiH����q_G�}�8�$��a׶�jϹ"�!1�3���)��̟_Z���%�~�I�Zԉ[�D}�����Yה3���B�S��]��P$�²��`�V)Ƌ�e���ݕ������h�EA�!W�2F�����݅4m��V����Te=�Idz��Xj��n�@OeU�ȿ�H	vK�_4ͷ8ځ0���[9E}ޝ�4�N�Ӫh�՜i*�<��,L��n���m&�R0� �{�j�n���t�����5L��KJ�~M���$�S: ��\���ÂO,ODL�r��H�1 ��%��)5ٶ;������Q�d�BH"+�,�a�~�A���J�*�!���0��8�̦U��;hid��lU6���)�N��ۭU�������G�ek�'-l�)%��\R($"���o��QO*P1����(�
JU�j�6�9��]ǟa�:��$�T��:r_�Xb]���
1Z_H+G�X�_!+��sDLD�@�a/ 4�wVX�%}f�x�>��C��Y: Pׁ�� �eM3U���3�b��w�
�����ƌ� bk�.�SR�4�Ib��zR��G"eH[nhսR��g���yM����|�Ϟn�^���?K��߭z2r����n�������AP=0H�	>�fE����V(�Du�O���;��)|��6��ٻ��~sA{�|=ۧ�rI�6��>ϙ,�y)��(;{uM.���?�?�㛱ݾ�ĥd3#$�^���{*~[6"ܷ�n�s� t���(��Xw/	�D�� /ǉV������m����s|�Ȭ�C_e��qʩ3ߊ6�M*���7V)��; �އX� �o�'=��	*��|��S������eItt�р!�����3��[K7%P�=Ib�a"�׿F��33�*K�U.%/�Bw�UI�tLf�&�!��^n^= �݂���7T⸆�`^��p�ƫ�h��Y�|��t��ED��_���_J󮗪�J�?�:yS��r�w}g��\W�o;K;�a
>��{Hآ��)�7c�FLc#3� ������o�veF�UTJ�ߖ'�����kL@���X3f2]����3���B�������Q
h�JmG z��yS��p0�2{OC�/졿�gr�FO��e�������B�������ZMQPe�J�؋AI���t�J�+���0���sD�Rm�͔�?p�&?7�sj@m��ˊ`���"��?1����ez2���ߦ.c��p�O�NS�)��ѓ<?z���ٱ~��9��_H˵;�.�l�_���$�Q3�Z^�8��C�G)=�n����Mh�	7�[�V���do��HiZ�bq ��o�uu�U%�\�NÒV"�m�QF�K���U��ֱH7�RxaL����flz�6ZN�#��'?�݉<�T�EN7�-Ġ����ǻQak��鴯��Z
s����w!��u<^�!D��S���*��G�k���}\./
��U���K0K�o�%я����k��15��~;`?�w��t
'�}vz(�$*G�E�לi�R5F?�ۗ����q��n��e���)�,�d
�k���a~�;4g��A���,��>j4((���Մ� ��� �cD!�Vt�N��`��������ƫ��+Fm��^��(��'n�{�ϯ>)�(��k��<H�#�P�92�m���n�~�^A&*b��F�����!������l��g=�Ju �����0�s�b3�[$Т�"$i�\��NҰG��"O�ؘ֗$G#e� �K���H�
���g�`�_�z�Z�L�U��&vg݁�\9�tk���l$��Y=�v�
܇��&S�4Ni��e���_������̷IC�mT�;��9n]�_�Fb�-H j`Lh�������jЏ��XȈ�>ڧ?��G�Tɰ\����Ե�ׅCX.=���8\O��=�!�mI��'�v�EZ�ߑ���'UD�'F�)��N�ķ_[�ƚ;���� �a�LK��j腄/��K-�߆�9.8$���/v k��ǜ�i �*]z��	�:;���>���]I,�+�a�� 
+ox�q�}�\e�ɷ^$�K�R1�_����
vB�\��'�U:]c��]��v�� ���s�E���z�RE{KC�8NFs�A�δ{�����g��Cps� ����YO��8�,x��`��/}x_$���fF>��>둵XP��%*��Y�F��1&���H�i��6r�'��Y/��{��*3ۧ3�N�j��ŗSm<��gJ�_	Ve��[�a��u��T�"Ω���S��)"$!:�7������f�5Rr��s��*PPh^.;��g>��.���7�7)�(�'*����MG^�ͧ��$i,￢����&�앏����g�섄f`��E�_½u����Q�ٝ�m����/��o�:�q�|U�U��߿q��k�C��_ĘQ �8��w9����-�`[�r:���m�᚜c���-�O�婨��`[A	�����e�2kg��Y�:�ʺ��J
�� E�A�\�xL�~Ӻ�E��m��_و0�lF=[��l��Rv����S�D�
練��!4�s��wiB�h���gV,�^nV�%i�m�
����Z$1����Zh��=���F~�j�6�a2��xP����)�B��o`�����b<�h~N�r���.v�O��tх,�Rn�����/��)�suV$Lnb��2R���k��p1�L��o� � 2-Ν��`p�4��=ú近%�U���3�YK�8��`�B)~T�^�[�W|qT�h�"\���ޜ��st�S�&�<8d�0	2t���W���j�Q6q_}�Dd�e4�|M~��KP/�n����5����nk���x�N7:�wB?u*�U���WA0��?3"/=MH�p�(�/͕;[S�5��ܹ=�#{��)rlB�����\]���`�}Ǻ�T�{�>I]tB0i��fVJ%����8O�u#K���n���W����/�H֙��[Dj���%wh����׊�v���Q��)��dOY5�[����^��b4~Y��9���\N�x*4�� �G369��������T���C�,ƿ �(�����J��`��$U}���M_�\$ۿd�|�%Ce4up�fL��%�,D�{�,����jYK$���A�q���^2�ۃ+�?��n�FA���sm�1��[*�� ��2���T����ZE;��")��d_��f�o�W�I�(�8:�;4�ıd�:]iƜ�(���U��s��8	��x���� (H���%��I��J�F����Y<G�0o�5}��A-��=%]��G�M�J�R鴹�¬�~vc���x3p���̥�����օ���p{�`��D��?��T�i�����A��1���"6�� �Ӥ����疴+^����aL,*o$����S�tخH�˖�U��4�^U���B�G,�>*>փla�D"��נ4S���e�C����i���⿤xw\�����ۨ�/k^��Gu^x���G�O�8�z0(V໖�5��q�ְ��Ҋ�Φ���Wh�v�%D)�|��@
���U��:j�4S�0�2Q�
�O�}�E�w�~���RD�=� 4CǖSH𺣌P݇M|B6���BuFxkf�]ȷ�V!�*A2*�F�nE,B�z��e
�q���/Xd��j�s78b�H���ǡ!�c�� �:FB�� �sKc���Yv��,�N�d�
=��q7��Kr���+V�G(%=	�jlY.�p�19����4@VL�B�
oF�X˻k����'b�0l�~ ��$��<� �
2E4�`f<Wǩs���\8P�e��IS�f6p�Y8FZ����]��s�_[�_3~�*���GG^Ŝ@���7bl��^� �*9^�$k['�D��A ?�*�L��lE����Dz�Z�]o���4���gMVa��s_��Ŵ�˖��l���I�RV�[a�L�WǙ~���/г�{t�m�\���|�1ei~��C����߳h��̦�AUo��$��V�7�
:^��<_2Ȍ�4?��m��?��^d%��T����`S����JES��Ս�D���	���j*�����Ab7�@�,V��0��W8����Kϊ��7�e%�ނ�����~��4�Dx1� Y�̏z����w�?ݬ�����`.�S|�f����|�u���&;
�bY�G������4��p��|X�bp�^�s�8-7���W�z�~���?<���s�4���a����0b��Qi<��.��!���GO3>t���2D�H9�4�ε�jf��@��+�V=�ް������,Hn*8y����w*��^¸U(.
Grlo}���TƦzx�y�� �4E���=�h2#�:�a@'�@�軀���@��V��x��l��K������p�wc�g���T���x��B:�����m��a�&v�&��t`�!� ��1����QG��{��dՐ_n��4�A����������(R�'M!�L4��.YVZpn��A��a�5!�«R��s�rٜkhr\���5ɐ���*��;W�J2�U��h4�rG��r���OǗC<)�:r~F��_E�����
�.�������I�$�I#2j��K�M]M�S�<c'����GF�"N�����/!/���-֠,Y���$AIˏ�x���G�n3q."h�����	BPS!-����Fy�M�t0�玻d�`��A��A�}�7�d����zW��d�B�l�d4�-.[���	OƊTW?�P���	���f�z*�_�~<=�
I���W�����L�pt����(�/G�d�"�y�lD
0|(?94���u��|G'�OF�ӕ�_�5���L��r�:�J�A��M2()>�?�?f:���F
�R���j� ~��[]h[n��:��dWk�G��L,�]#Ǐ(��%�O��9��>]NR7�5�J��ϕS(sutkbu*�L���p��8�Lk>X� �B�xu����d��l��-������w����)��s2΋�����b�8���q��)��=���
��
U�=/�,L7�ۑ�����ؿט��2���P�П�
l�ɫ�nBDդRp�l�m�ryuM_�X��<),��
[a�5��2��a�K��kw�42�X+�0n����Q���,FUX7��V�3�'�#�S6�Y֓��AP�먘�f�a A����'9֧�$�T8s�c��/0?� �w[w]�9u*WN��%���*�p"��a� 5٠gF���_	�� ���3>݈��5�ƃ��
�ⰛN����ًh��Ĩ?���/:S��i���3 �d�7���?څ�x��$��ƽ)����^1���{s)b�V`��F-EY%�;�lr���� ���zQ]��9R�u��Pަ�U5�)5�J������-cQ��nfʌyjf���`W6�ӮZg*�����.��Q�I����j���K	c�'�otO�~���]��o��x�&�K�^� ��7l���4�_>�&��GF��K`��������;�P]\4O,��٦ /�����2��,�񽦤g)�����V�e�����=� ����|�?��kv=͜ڴ�Ġ�'(�k�f��U�seʢkSD����fG�m�R����1�C��˺���u٪y�+8��L�I��[a'�$U?� #|�D��"~F�E�4�y٢D7�?�Z�7���G������kt��ݷ9A�į6���{
���/�f�k��b9�a�hx��PR!�<�W��2SMɊ��ث~�o,%����=Ϗa��7q@^kѿ�b���$ �B_,�Gu*_'#�3��6q�<h�;��<��N�}���7y��ib5�@�eE���D҆�����o�>HtĤNJ��Ye���/��IYJi��w�R@acX���
64�G��DhѶ׃!�}��eՇ��*$��gG$^S0�D
"xĂ�1����RK���]e���ھ:�ȣ*��8������j���҄�q 5|�%]}����j)��a57:Q�;�-�(���6�A���g�1��y��0�ʚ�'�h����Г4a���4��B!�>$<�dU�r�5ܚ7}��Q흓RSQld���~v|e�6��bݦ���V��%��+4b���@_M���{��	�{�Ӓ>�CK>���:�d��ϳ�H����=���B4�%W}�[<����s���s�����DC�����t���J���t+����r/������|0]x,	S��*�wD������&�U��$����t�������*B9�X��\\�,H-\����Eg����j�?I`��H�����Kv�b�}ڌ��˥8��*����;�i]ݯ�����D�6a�I�u9fƫz�1|t�z��<�C���%�c8k|������
~1���.�fA띯`�yv�s���ܸJ�� �̀�1��t�q3[u�m��hT�Ȉ{`'
��Q|�>x�+�a��qXK�4 �����҄No�=��^V (L4�;F�P��O�5�6��˭�%^��v6
��z}h��\�R2:~��֭OS���ˎ{�u#G��u��#~�]z4�ƉzyP�k$�lpJ�*%�}���ْ�R���.[y2��)���?̃g�)�k�G��7�]jeK�ѳs:�z��W�)8~>w2"̙�5����?�p0B�c��#)�bd�t�����Rq�U�K!H���P�vY���Y텸�XMbP2��$���u��T?
̆�����F}16ն�9�i}���\'mu�`���g�h25�v�����Gc\�,���U�������;�����o��SO�ىQ|��6z�^�:73i��!;ʲ栜�|��'�n��oc; ;r=�n�ס�ӡ�"RGu)%�|�}r����U�gnz����Z$W&{�>9[�V�"��-{w�B�T�������� jrIo�������*/�:��)���E8����H���������!���跈�	<H�,��7�,�MZ�EA���Iˇ�p��Tl��%$�y(��'�W�ME�_g��	�]�"���f�*b#(l�B�^��U�)��ո�!�1괠{?�9ٶ��cC��щ�]����CY�N�YQ�ZV��"��s��HqX"�|oO�/����K��:{;=��߀t���ll��hw�9aj�����:����͡�h��,�4m�_���ƻeL��8��)J�T&_��A_��[�7��o��ġ��'��S�����z��T0��%��"���+�޻��+~=�pe8&����Z�㢘0l��B�o��N�HAr̫��/i/�-���l��>��� �h�AUf�(%[n{A+v!��̻��D��Ҍ.�iZX)l���R���i�W�|��PLi�??���Ai&{�q4]C�� 6\ϝNtMD<��g�ap~���]��\є��ɻ�fh#B~���W:; ��(D2*n���(_6e�O/ي��a�s�J�a{�����^g+����R���.���l>7�,f�i��?.�֪슿/�@�[�v�ύG����z����#�;����d)�S��Os��>�ʗ��������Y��h{�C���� �	�F�/yه��(Fip��A�:�.��?������U �0'�<I:f	/eK�2��Q�'�s^�/X aV�����kY'��?�W_!
��gneyW�| B@6U�ov�c-L$}	��Do��s ��[H�'�v���g���[�ԭvmvj�������\6�C`�*�W�[P���&�d�.T�σsP��J��i���Tܡ����c�B6�r���U�G'�P��
4�/)*re}�l�B{:��4$�b�0󶻧o���qV���r�~T��|�+	"�(��KHu����Ђ��9���Dv܋�6h!ҸCLm�!�ؘg���Dd��
�ج���V�_��w�M\�g��Rm�����,��w�-�yOB9�$�+�1`��)nb��lݖ�<hʔ���~��<�@-�J��g���u�@����m~|��z�oxQ���Kl���C/U���
Yݸ3CPa5�>u��o��мa�C�o�g-���QuK�6$������=�( 4b�$��y�"�5�oև�- ({����C`I�t��PdV�y�����E��w�ª���e���qj�ݐ�N�w�˰����T�����k��*!ۿa����*���A��ZlkB��ړIn�y&�ǐFP�2�a���3�64�]�����E���Eݐ,0%�3�ֱؐ�|<݅25G�n��G���2�X�6���7��4K:�Z
`����0t�v��(!��Ό�����*�_�
Z|-�K{�����xr`��goa>^�|�����o�&2`���,/e��E�9C n����]��e�:�<Sg� ���Q�8���W-��V#a*S�1	�e����[�ۙ��T��Н��������&>9�T4���(�uR�_�1�ta�=�t_&c�(����|�oAJ�_%7fTJ߁��N��ND@s��N(%z! \L��堥��U�����b?&�����}���yMI��~h�=(�$���5�	M�(�{��1�֦�!o�[D	^g�[�oK���&�~?�1�oe�Z������c� �'C1��:���.Z#�A�Q6[j��ע�G'�U�`Qgp�a�v[�Q#ݾ��+�V��������P�J{�X�����مq�����;B`)8��TDQ��:1r�"�;��YV;@�K����D�j����ΦhE`�
�S�5W1n�$��Tx�V 5ϵ��ӤV+�jM��WⱾ��M{� ��.ʸ�E�1I��D�OK�s2�-a���.��\�p�-eSki�0��8��3��_�󊊘נ;H��X�
�P{L�4MQ@<C
�a;}}��W�lς���,�ԋ�Jz�0��=۰$F3�HZ�(Ѡ���������=�d��x��p@8��#M�z4 ��!$�1���w��|D�;3}�PW?��a�4�3뵣�(��[6�^Ȧv�"$���*fk�??IZ���G)�����S�7��L�W��[��Ѿ�ʛ{I#�R��t�U�VGt�N��l;s)�� j��W���ǿ6�<ۅ�}0:�kpgL��V ���g<�؛���U��xꄅoWF�ڭ�}��4;";;O��J�3���-�d�n.vOS�e{�ʶ�3��]�þ�2�
yR~�T��u��s��Q0S�)O���#m�r͏FV�+ c^Hd;�q_�ģ�V%O����F@_�4z,|{���;#+��4 D>��X�dT�rǡ�Ґ��I� ����]���t٤���I5ᦄͰs�oJ�캥j�z����q7��ɐ��+��{�yUB%�{U���1uY	N'��hW*䕹T PAh�ڬػ��Dsm�X,C2� �U�%p���%�j�j��^�:�z��4�-�����ƴ9}��.)wLb���Y9p�=��0�)
<�+�áρ��8���,Vpn?ڱ�D$C&�ޫ8�)���AGq���&⣾�/"�l�>�=ȿ,L`f#��=<�#A��WG]���i&M[o岴GȐm��
��3E�Z)�^N�
��Ey�r��-@t��b�"���J�OK���5���v���jfC��tq��D�����$�L��LH�a�!91���p]\-8Ri�����z���6i7Qf� ����f ��|�q�)���Q8=
�]��;��s���E��c��<Y�NS��)6�{wV�^v,S5�-�~��*Dsx)A�LS#��m;.�8G�'��3��5t{��m>?�0ؼ�"�l��������� �P|�h-�Rfݳ�A��*��}w����*������!4WF
m8J�0y��i=�v֒w]���`�8jt����Gͦ�Zs|�`�8����Ġ�i��@�,LV�I�j>��/�j�2 E���A���w�_;M� �|9�~������2�-�]�ק�c,od���r=��Ϛ�z:-�22��LL�}�1z�'����m��˗��fߒ���A*MÚ�d	�ƀ�=�$�y{�h4hPσy"2�c������
CƆ��vv���JUF�ک����C�1��h��qϸ�M�����y�u5��W��?mJ���=Ra�0�$,������e��\_)��x���t�3.)̠d<����]���|�����=�����8��0f(w�)�h��hMR�Ta��b�V8���2v������h�+��S�$�Y!G���}��B;$�("��}�ޣ]�|'C�Z�IR�!�3z����Ŵ���
Z��`���-Ɋ~\QX��fU�׉�H�=JL�τ[���ym}��	g��T���-r�e�2Y� (��'^�������v�����z�Uc�\��ԍ��xL�"��6�,���h��ÂL
�Y����N��"���~F����DٜΫR�z�K)?I�Jx�=��7h=�%�O��;z������N��6�Kab��> ɝ?
5�KyV����X�;]4N��5U�@�����A(���B캙pL�t}�����c<���7Rp{	j
wz��F~C	a,��u:FVCᗇ�� jl/i/�_?�|���&栁K�6�^�3~\$�PE��w���:�蘙g�
ثo���(܏�0s�W��uK�!�dK��O18�aR�V��2չ*G�����.i
m
M4�a�
%�d����v8Zk���[��=�va�����U�]�(�7 ���6�����.�����]l=�3	p�D6�2�X;���K:�*B,>�`��`�5���0)�#|����~����@�m�x��	![l+�KV��M>�~|�<��� ��6�`���e���8�ԯ��g�}X�(,�j��$:؍�n��Ho	9���0{G�N�n�����;݆��_Q5�Ds�������߰�y&�,�Ћ���ɇ��b�X�����R7��"�f��;��"�	�x(&%�LL�Uh&Wt^޼$�HT^�^��� 's��t�Bj��
��Sd��d��s�.2��_ZI���_���:R� ��d%�K;��oX���^1��A>����;�ESJ"yP�/�ђ=�Φ$	-OBq�'t��f���]�3����%�hq�RT��,�0��TK[��U?o��R(�M�藍�A���[�F��űą��&m��J;Dov�bE��׷[\��ŜIv��,�ZYc!{=���h�H��W�7|�0cm��f����Bk��0����j�= 6��,���j�|�ݷ�ϭ�1��5K7�	P�ի����c�n�{�O����<�!Ԥ����M(U��AN<���$(�R�Q(�����r��HH�a��k���*9i1�ۇ׆4�c��r-:N�ߤ(�yV���h}�&�1v�+��As�0w��鼥Ni��%���򛒜1*CDz��&����m5T��/h_uW�IWD�{\����/9�V��hw�%�:�FR�~�D��N���~�/�t�	RSM��&{ÇOr��F0X�F���S��n��I�����-�����l&$�G�v�uA�"wP��LX��hjH�uO����-��m�ZHɯ$a�'����I4W��*>��
}�m'�bT)���g��}�9ۻ)�7 ��ґ-�?���^��j�;�Ã��|P�th�*]�gQ){U5-AT�"-���5
���P�hWĨ�pC��uZ�_�c��41��K��'�@�����AA�(�N�n��ϒ|�p�J�]��~������X��i�DqtQ�L|Az�q���-3
ɨ�qN��g��s�
c9�.#�h���sq{]�yb}fֶ��(�p�E�&AKa�N����r3�"�c�pvŤ�f2y���i����>L8��/���{�O�i�Z���8rƿU�m,�e����Ղ���:��15B�?���\�k��	¡�+���!V��lX���Dm�U�Q~`�w�rѷ1��(k����:EǈV�
��g��~��.�����`�	.�/;yb]�*qΩL�<����j��F�]5��A<{.�(��|���	��	r�
�*�a��B�I��V{J�ek�Y��(�27Z�6���>?]���్��C��`^��L�&;O"'!�M_��Jp-K�Q��3s)>��|��w��,�P��,B��!n3m���\����pCT����'��1Fټ7#����_U��W��m�y�O=#i(Q�N���2�X�&j�1 �g�U�P��N������F���6�$Я�� ����͘��a����������OG\Dᰋ�ڇ�J�k�uR�ܧC�/�<"(��0}��7�ë�ɢ;��( ���z�[�pv���M�� ��k��˝��c#�&���]qIxS|x���J.~<#��{T�-��Rob��9�"����	�Q$
�R�	�fD��5���&t�IT��jd�<���nQ�����@���dk�]���ͯ���?}�B��s#���o4"���_#@~6ސqj��u�,�&�""��+�w˵���F	�=�%PõJ����mpJ�٧*U8]1W����H����b���7-�+�������آ�kp�bh���M�����Z�_rմ�#���e���h�	�c٬�S�W�n\ޡ`�h�����~�\B����x�x>ͨ��j�3�X7?e��$�Y58���D���m����S_��u>dx��m��0`�>�Ze���'<#�B�۲�Xl�;��»�;2��x����%�=d2�a#���:��1���ܝ�Օab\��:�Hs��O~�U8ZH�hG�R�'7	����ѐߔA27�#],��<�#�}n���L)~�`n2ȋ��#��� s^E'cB Z����į�����.7�9ǥ/%�n$+�o"q�6I�ر�`*,������]��"����t~�?<�9!H��Ԍ=QM`���g��h �A�H��Akf�e��j�<��8�N�F}����I�V;T�e.�o��{´��#=���U;[UdlT��<OH�$I�?d�TĿ\��a��Oڍ�����\� >��쌈��d/gɤL��w�W�ᗄک�8��s˔����JS"0�MkJ��-���!2� -At��h��?��g�K��b�n��­�����8.��G�(��S�K�e��-�[����hd��CCD�|dr�ɢ쟓�S���zK�����f��ۤP���N.w��F��Td��EW��8%��	�Ld�X �ץ�[N�CK�s�n�����Z�%x̮�b�E!9�j�u�R��N�Q����o�6��U�J����Z�)A�&�TԌϤ\��q$遁���ī%��(S��W�p����nG�~�)i�SK�����cw+����2��ԗ�b��ݹ��Q���s��Z���r�v$$��U*fn�Yi�Dmh����N���h`�A5J~�vN�=ߚ|�9�_e��F�7T�#��јjzR������Eo9�4i���ā�Z^���OK�М����ى���vl�j��t-+@���j�@�d~!G�
�����ƍ"�@̉���t�@�����w?����?�����ez_�ȉ :�A�Ju��5��Oz^����
��e�6s�C�ܕK�C��_U�U2����'w��Y�y����W9�e�����;l�����3�����z��K=.ñ��:a�M���L� �����5h�s�-H-up4�iA?�<C/�(| �!����ط��4��
��%�����	�d��Or�;	�}��]�R��l���%F�d�wUF�f�)��q�Rt���ELcw�@��m��F�u_n�cCm�� Id#����z����#���`h�r��)���	��*�c�3�꟪�H��8�j߸���6hۖ9��.:��_ݴBN}�(}��7��qE|$Do�g�h��O���$�l	������t*zu�=�6���������98͏P�'m}���>�9�#y<0��(��ډ�q��nރ�w�M�N�h��0k�{Bzr��W�7�:35ͦ�(� �=z����ߠ��������R����^X:��� /s>h'�>�c�*�|脽Mm�PW��-�乢[�՚�����ɴ=�ۖa�E|���h��_W>
�aap!?i�[|d�x6��L����{��+kw� �b�lB�L���и��>�ѕ��O�����'8cE��6>�t��aϟ�S�79�f�׏��(JR~mk9���@����M+]�7&8Q���{�����闘��U��2h�/ѝoy�5��KB�~T�n�"��*E��vI�H���Wt��O!j��@Vz3��$���P`���2�yH'ܕ_TVrt�X��o
���u�<��~�`��OQ�Xෑ�؅��LE{���c\XsQ�?B�a@c
9̨�ǔ| Ы<�h�Eۏ�jf������F����q��L��I��;�� E?�t5\�e�F=�Ѫ�-r�F�ƅ�WLY:�f���_Qh��T$i�ig��7k�A���&*f����
�Zm��(��~I0Q{dG��q��'5n�T�����#��sr����y��o�FP��h[j���M��xi%��8i)!��e2�[1t���Ҹ΅��gψ�QPz6~pHT�-lO!8�}���ps���";�������.�Ox�|��E=!��I�@��:z�/�/r^����.c>E�8�'��1�A5�3MoB��8�G=�N��X�(H)-Ml���(���Xl��t���LKQ��[���`~��lW�h����)�����b�����&�X�iT:��9$����P_�6`�ON��`K�	����ut���U��?���\�fck�)�s��z���-�&7��nI�x(�����/���a���cw!k������BÒ�ڨ-��j�g>>��k��XL�2���V� 3�`��:o��0�*�ʎ��s���#����j*>��e@>�e�qp�o+���?խ�!>�%�.\��v���=���ob�)s}_'����@�(�P��x���C��C����EG��ZA���{&Mn@�S�M�� )J�7�Yw�1? Wm/X&��Pă�H�(��>6�ë�[�nn�A���ZE��";�#kJ�y��7��Q��-u�cc;��:u�Kؼ�Xu���8��r�驤ُ	�c�G�r��afTQUఝ��c��"��z*�C/�Y�|�EĿ�"+�!�v����*��4tO�� D`|���&m1��O���Ĺ^�C՛�G���чr���h� ��_��]�F��Z�#��<���ѳ�I9\ǃW "l����{�ΐ���^�h,����j�?-����_1Gt�&�_��'�Xژ��'������Q��
�
1՚�,3�t�H�S1uY|�'�N\��U��>�9��5���uT]���8��!��_� ��-Jo{e}������r�@�u�7z����6RK8��{g����ǀn�
-^E<��o	���_z��{qfС�v���?AE8*-�u�@8�("�5���=� ̛X��8'�4q���i�#�W,��MLx�è
��d�Iqx(D���^�����S	�
�+i6��fp�ZYO��:v?��&&<�sS���<��vB��a��`A��xB�'�
�t3�^qH���pU:�ؓ�~���� �%Lk�x �>�
-�<����(v��o��UR9A8BILҁ��mݣS�+��̍�<��I�j �ץ�vm�n�(�"�Ry��.����a1?�o�G����N|�.ePH�gH�]�S(�6��p�<�&A_��Z���]�9L�{��K�goH�9>!]��S��V�{�8���AKFY�PQ��|t�_�b����ݗu��D��њ��ےE4�冖�1��(ΡV��jr�� �F9C��/G���J	*�h�j�fx.��ރ�J�%	�I0\�Z�Ǥ0�QZN��s=�'�:}4?���}ݽ���Ӳ~�������#�ɴ���BR7O}z+�3m��c�LÁR(6���?w�5ަ��+qC�0`%*�8U O`'����v�<�`P��:2�_��x!`A�;�:�GfY��u8�b��2���������yL�3���rP��ؠx������b���A[`2��"X!9�RgMv����%�:#�e�g����W �Z:����ŧ��JIe�J�.�I~?ϝ��R���,�����mz�Yn$`��m
̓S�x@@�K���b���w)�bt�#�kL[�h�^�=|����=}�]�̯�1���Fʂ�]�{�%6��n�����a�N�n��J9Z##oR�Lu���#�z���hy}z�]���UVF���{�z�^dO9[cB�l1Iݑ}�G��=����Iz%�T�OW$4�qi��� �l8_M-z{�ο�튉ϛw�6A�9G}]���A#�ϣw����c�!.7���K[$�C˽���h�ų�����OCo'���F��V�P�+��3: X��'�C�m��?"�{P���l�ymuW�Z��j�	�I�M���yh5�dh���׹������3������������dXh/�U�zj���y���s}��B��L��ì*ꐼ��OЎN;�;�4�`�-�dB������Bp���5��.6�����	D��+��N�/��&LA~�/�oA���| �,i�u����XipIv�5��:�ϰT[f���	�'�\ �#�Kx>��s\��ZW�0�E�1l,#E�DD�a�G�Q>�?�����Ƴc.[��.�d�e��0����FTJ�C	�^J��7��L��5}
�� Ib�%E���N��%w7��>t�Z�Qҭ:��=A�~c�0�A��\ϧ0K?_��J�J-�DV����E����t�Qƾͦz}(��MN��bx-�[��
�a��dAJ$07��=rY/�# �`�17���n�P�D��J\�cL��G�Y�SYS��y��h2���q�@�1w��Y��p����ʋ��i���>�B�OQ�!��u��@?�L۽�PW��B�/A1�����j�r��9�QuQ DُF��K�5����7��ߚ�c�hB��$�@���r�����̡�Z����&�^\�ְ�f��=e�����V�v�����K�eJ�@�脀O�S��}'8W7��n���A�N���p�FM?+��?޼��ieA�� V�T`n,b>���;K%���҄�!��g&i$~P)�B#�ǚ��yq�f\~��/�����F��?�GL�mKQ����E���h%Hb��>�X�(V	��Һm�Q��M�1�E��o��$����vE��$!	������v�K:���ئ��?~��*>vY�q!��:Ӕ��n��!�;ɭ��灯l�g5|���4ʁ�41��A�9q#O���$���C�ƭ{��U��[�Q�<F��M�僴�=f@��U��_d/���;�3��}��F���:L.�#��O�ۂ.�����T�I��Bu7u?�Oi
V$�hkkD�(�G��S8�ﱖ[U��<���Aó���� k#��?I/��i�ֽ�zձ���t�}�"�?���X]pa탣��Y�"e��)�%�����tλ8�!���r���Ѫ����Z�E�2������C��ՙ}��ٲ�_s��Դ@�ӌ��|*��.1�&���TE	OF
���AT9$��$e������<��g�y�`E��k�?d؉T�L]��ZUe����lS��.���^X*�,U|Z�O($��؍
mpF��Dֿ�!8�w�u���N |p�i;���rF_��{�n��/*�`��@����aKLUi����{4,@&�ܿ�Ρ��$����w���A�U��}�3��D��+��',}k���Mx��&���烉{p��៸��/n�D���VP�$td� y;�����]qK��ޔ���_�q�E,�޲EL�3�Þa$~t�Xo����:G1X�8�C_rh�$y��>�%jަlS=`?i�%�og���ۧ��#p�vT�9�:`&��Z�8�^6�v���A~�&�(P���l�lC[H�y�?�Bh�ޱ��d�=ڪ]�:�q:� ��GW�(F�Iё�w xh�A�_.f��Cg-��>2�������ތ~z�"(�h�ע�>�Ѥ�"r�ѡ�����q*���q?��b��d��/�vj��*B��P�4ƶ���#��n���i�+�y�'���m�&&�aMRA|��C[����&�"�Ad�� ^�EW� ��r���y.���OU*M�ǗG��ɟLɒ#	���}�1�rj�8�*(Q��G_J��q���eJ8[��D����eM��Ʌ�Q�
�o��C��������K���ڋ��H��pF숽A��?�,��-� 1D���9����k"B"N��?����ؽ<�*ʼ�!�Wq%eM(p|�����T%��� =u����e҆����.?b����Aᨚy�����3t�,��ΛQ��1�8{�� �s6�5�X�
5Ч������*���W��Rɳ��vi�X�2�_e�Ȝ�(X"D ���3�NĿ�c�����n�c�x�9�/���܄��Po�@���i�b����-�Kg�*Wf�'���tCУ`'����zc)�L�5�!!������K���{��%|�T�-�!+����~	�@>t�(�k�(>���"���;@��6��&D(�d���(4������ti��U���S�,�(1v��%�B�-2%�F@YUZ�c�W�q�'7��[A�-�)��n�~�U���I��q`���ׁ��_�Q�+�3a�9���O�] �����FLZ/� �����Q��8L!�F���m5���U`�6����P�R��WK�����(0�Zp�n���w(�E������?2��&��y/Y�;����@V������,�<��mu?Z�Z�S Y��p��z�!�]M��E/d�Piu�^�)�4�!w:���e�2 ��r��{�SWT� ��������ktK9�h���5}$6��`��z����	b�A� #/�-8����і�������8l�}%\������Y�݊'�({��.�<���( 
�Z����k���0���@��3����|��ዡ?v��>a�����X~��ɗL����Y3D��&LZlY^�ݽ�Pq��@h6^�������Gv~������4���*)����~�E�ˮ�(W(7u�NL�{��0��K^��?8���ko�!�����ƴc� _U�M)'�y����E�C��^�9<@!�������*X8�%p�<"�P �ہ��Ϋ�s�	QLMA�'+��QZ�K[a��F��"��h���x�(��d�ƪ����xݎb(iie�ږ=�x�bl[_�-���9�]KN�.��I�*�t��⁺��-��bIn�,}����UJN�L<�V�p1�W%4���,�Jm���P����>�t:�e��+9w��2	�	@>��&[���/W]�&&5�Fs US�cm�&�BD��nS���*�uFkb��p'��ũ�[��I��5�������Kg|�晼��@]�U������1�f0�d!���_�-�H�e��=7��ߝ�2r%?�?��gH7� <�&�ُ�]:�~�&�|�*,7,��(.gꕫ�"�$���R`���dTF���r��GHCF"�#"�S���D��Z%mO��_K� �t�q��4��n;b�xʺ���l�3B�?�g�Y�X��d!�TΗX�Ok�r��Bși
���,
����@%��C�_�l�-�~o3=@�+M+g&͟�a��l�N�8��D���W�M�q�����n�9�/�[���o��a@ZHmN\��06�;R�9b`���m�>�	QFL!�Z"Iu�t��,B�B�t��R�O�%K��,�!dΈ�kİ���V��t��5�>�֠�sМ&��z�c��\RCy����"�V�'�	��_gǸuLµd0� E��?�\᠁S>2�x�)���<Jᥥ�T{�W0�U�X�6��i-���� T1~��/rY�Ҕ��U�-���u���k?n��v@S������g�t1����9���"k��^�G��I��C2���t��N����\���9�[�����嚯��(�L� �[BE>��@�x���SP��z^�� ۗ"M
��_�-	�A:�x!����~�)��Dطb���F�m��� u�0��e�t�>�;�hm0Rx��iSU����Lsi3�V~�Vz,����7��8��3��r�1��Ihp��:�Y��)!4����;�=jK*�)}��$�bО���@tWk��2ځ)s5�u�;��ۇ� C���[�~$����{�L����1
W�z��e��l��̴�Gq���v�Q��˒@�庲e,6�x�Z�mz��c�+�]l����r�7��@�����.�h���"ﮥ��ـJ���74p��}�T�E��F>y�T���M�M����)����4��P%����y�]���h �ρ7ϸC;ނ魺*���vP��A�T�ܫ��>Y���R^�v�����&�X|┍��r�F���b����=/tE���-�k(V\�V�g�	���$꺱�*�F�T�'���Hewv]&��r���,��OZ�6>F�.�cc-�|���<��^yյ��ȆY�!��#�G��N��i�����@C�	�Z�f�M�����&�9�D�u���"�P�oR�k;���2č	��My���ms�b���?�N$\� �t[!�އ�7�v^����uT�{���#����A�A�B��N�T�y��[���eoq�O�kh��a����QΥ��N@ѕq�j��Z��9�b
�m��,�k��8+����?r�-?�����iă"1\��9��*mMi*���"|8\>Ƌq|�t��)���o_�^�ASbc����VvTHk��н���}����FdD)��E�n(��!��0������z�t�z�akĽQ�P'���B���+6O����T&*�14���XϽcn�%e|�v|o��Ĕ���ԈN�?et�������{Omm���7�<*M3��}��2k�������Q����:F��`,@���O���I$2W�#����K�ow"�)��)�TQ*U�'�2�dj@V)���8���Ǉ�p_�'߹�O���T����خ�($�8`*或��D��^�gi���H� ��+���D�%���H�-Ҽ��n7��3�04>������Ř��2��B��r�m��n����g(�rD^��.�U���n��5�X�=�zu�<<x�s��G1��.�2Do=�!�.�� ��9! "�c�#���%.�G��}Wc�*�f4�լ?������5d�Q(\	�M�ǁ�M�{Oi���E�z�d�I<t�lJ"Rn��?,���>��5���G�ff��X���q���A��K[�Q��?rX����I�o��ƥ2s�@��s�� U�V&�^�D�j4��$b^=�"n�E�$:u��KWJ�^���%�}�L��fl$�)zI��o��x�� ޛ��R�wM ��B�o�n�k�I���q�#I�I����$�l.����6��\�"`W|�����^�jk�^P� Hm0�IPe��<j�N�??9j�OuM���,�+�.p�����}θi`F�������c�O���|�;�,�o'JZ�����Mͽa����d���7���`D���4}��('6$��%/���i]b,(;�X�NcǡJ�"�e�{�1����hQ?j�u#?��y=5d^�TVXJ��1��0���ئ�]�Aw�Y���?&6�a�^���v��H�������E�	�H��R��:�#Pj��Dvrq��4Z�yc:mS8J�ړ��R^��_��l�*�F�۲wO5���+\/�c���� 7�>�x��Z*x�6���V$j��TP�� K���Ig�J�@i��Ϛ��
)*��ѣ��`i���!]�ϠD]9j�u��|_�(���Ţ�Ǿ�ڃBl�p����������h���]}���`8-C�R�&�1Jk�������iqK:P�D�G�П�C��V�_��ѯl�֐|�3�	�I�\��S�٤`������f-�I(����gL6��w��I\�W���fV�%�p׌w��"95�}؞^��P���8D�o���pهg���R,�#?~��'ǈqٶ��*2�x��b�`���K�-DQ	�|9s D�6��cx����V�9��{�fAL�h�w���Q�ڥ�%�#i�8[���O퍉S��{�*I�૛@b��y�D����AJ���Gw:�fď�j���D5��#߫�J<ېN��B*|�P8��l��ďg.X9�p����*�Q��	�Z�����=�f�cv�����W��&�J��X��_H�#�E�Zm��󵈽b�-�*��"EH�Y�n_f_�Zc<k(���H���$��Lb��}�!��[���}�Y�?�6U8�iv�g�yj�� �}�'��D���
Sb��L���+�yS7`A���W#M�c�=��Kcn����[�}�Ro��ٌm���������E"�%�}h�?�m��D[��38<��NG�9��?9$�R�*D�7�=�`܁�����+���ⷷ�63?����>������t����7;��:VjȭJ掴�"����6�Ԅ}�Y����|����^,m�q:K����LǷ����4괢sz5�ܦz_��>3Z�"�7��r��k�9:�a޸RU�,ݑk-y�x��[*/�x�?���J�S��E�)uѓ�=�u�NҨ��	;�&���ʄ6��i��ds����Z�>�C;������mЂMW*�ԩ�:Ξ�c&B���V����	��4�і���HG%,)���yyz-2���5�d�L;�	YZ�e'Yx��}$,��k
t����"��1���Ok7���X����j[68��ד@9b��|I���I@���W�f@��>/�ȉ㦺8+�w�5l|R��K~Z������)�.�һlc|e��c���9�,w7���,O�FH(9 ��K'w��UA�D2jl^:��u���D�t]|�P��_��|
n�*��3%���Bb�C�R��d�ַ�?�%+{�.��MY�>r3����G�V� �RM	���SP��+�@4�*l��Qq�ǒ]_{�r�]�'��}����ө�;���	�b9�7�d��î%���>i��*ti�Z��_��`�&���#�L��[
�a��p�h����;�p$��xFN0�^�~s� =T]<B��O`��<�G	|��.�?>�ЇS�?�YV#Miq̚$`V��:�B�	,Ov�