��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ḱ	I*�n���}וLM��!lА�(��p�&q�;y%�(���)��_��>�>�l}cp�o�6��NO�3�r'{��?�u�>n�� ��<[[0�¿!�csY��[i̺'� %Z���٣X�gG������v��VW5a-��玀��[F=V�o���H��Y�X���L���`��|m�-��a݋>=�+��TGZ��.N��Ľ�Ĵ��Sj���׶��\dr}A��==������Y�6N�
�;�*v^��rz����7�#&Md\'�Ŗ���A�<]-<:�,�y�}_�u��o���=�0'�bH{�z���Q�W�c�ع-ukN7��c��	��Zl�������9i������l����m\>(���<�ŉ�{��׮ �] ���	P2��jK��4J�] �F�wz������$��ܩ�����IZO���2jE�p0J�:��(�4Ͱ���*{�9���K�^�h9Ec�p���t�����STo���F_�C�f�������|핓�0嶔��#�4c\�v���1�+f�:RF��2�%�04��6����A���k�@9�DE�hA:t@JZ�H���[ӟR&>$��,�M�1�]�TM���)}�K�g��h��/�s߃ m;y���z��YXڜZ���9>'$7�x�+���_��fW,�������OB�_�4�ȏڟNI�MU�fhؒ�E{p.��0�'��|�ݗ��1^��B��xۀ*l�K�̵�4���m�5����W��=|*�c���̲��X#�c4p��V�2C�w�	���]���B�(�抠�D����Z;B��N���F��׃m���y��(Re�����Oj�8�8���Z�Y������.f���C��y��=rŅ`�O�d�O�޹S�9\:i\�0"ITpce��M��U��z�"<&���8jN���w��de:O�3"�g����^6߆��ᡐކ�� [���J�+��p��q����s5A$�3�@O�^~heD��[�L��*��z�ԩ��P���_�˿"��ɖ����SN̥+A�>u��>ߖ���Y�e/�����s��L�J�H�����+l�c͐&$� b 3C�R^A^@��1�l�t�lM�qc��=�%�0�¯��?L��`�P)�@,���]7qͅ�@�����p��+���
p�ԗ$B�F ���l'��E�»x~����#U�Y��R]E�7�D�l�)7�v�G�2��O�w%�Xұ~�5��il�>��~hj���P)w�/�|E1�j[���[&<���V[h.\*Y�
7��.u����C�>�^�'zY,�1$��{����,B������ƣ�$�9&Its�~�f���-f�nvhت�),�"O[�Dqc�����~�b�*$r�t���i��A�����F!���^�K �=h��z?�C8=�+��!�!�����
�/�^6L�Q_��IIT�n�#-"#	1��Y\�A���g�Iu�K�@�$<J���2����m��n)cf�\�f�B���μ��c���No��̎��5�4r�76���T���[v'݇n�=�gLϴ_�Z|�k�g?��dO�إ#�Y��1��u��K,d�O�u6�_�t�L'�L=�f����	@ �?s��Da|��D�0X����OR�U��&i�&CH�m(�%�6�v�\&��|�n߻�Z��oG��\���Q[�`D����@r}'�͍.��Ieg.�H�ZW?*Y���[%nitbj�@3mб6�2�;S� m:ܱ�]�u��t��T����k�]�/K8�����s[��M�Y�\8v���D�P�p�c�3����lb��a��l4��[ZP����V&�7L�z_�(���o�F�O��~�:iT��w��g�C۹�X�㬷$S��d�s���,���[`�*��u%�P`e�K����"mЋ_�N�:�3
k]�����j@�����Zl=���%��L���EP�d8ϷWd*9rKP%I,��b49��.���o��<�b0��*���NA�1�-���C��
�����؎ֆ�_F*=]~�wFa�k�@g���6li���d�+��1�钶mC��[���d�a-��"�e/�eG�|~�7�r4ey!�U�I*ً�2�Z���[儵�߂DQ��}4K�-�~�dq����*p�2o>:�W̴[YdZ~m��jS��8b�LF��|�::[]3�I�R�c�d̳}p��+�듈����=[�����'P��o��),U���\�?�
]���^Á�	��a!�(�p�-��u��&����]�~��\ }���3�������2�d���/M#��R����M�v��CLW�[�P+�֫�.�^��?f��r����[8V��߹�8�D6ې}1�VՒ�z�[
�+yM�_n����=�0��2� A�EH�`�������ا�1%��o���^O�gN��J�~�s�h�][�_?{t=sK�%�Q���2�'�� į�67����w�0�����gi&O��
m�EAo��8��piͼ�D������vO���y�m̩����G��e�R�)���WfgQʴv6d��#e��ul۝��JY�����4�"�_<
B[����-�oio$$��9�gt
\@����=�b@04vgM;��,ʹ�d��lBD�Ӫ>p���|C�!�춖&ֈ8l�Fy���i�bb�] �y(/Tp5Q)X��V6�$�Aǀص�Z�S\>�wfZ��au��57�	Q�J�1��T�\E͞Z��{<��q��g)������d���v�}/n?3�Z��U3��tp?�������%�6إj�;�r���d;��@:� �"��Y`���I��Mp|u0d`�s�^SL��j�AQ��Wɐ�t���I�������V��Iy���'u�cT���&��"�f{>jE�N&���9`�߱Y>wo����U�F-;�����_��B���?�Exc�E��nh��%����������l˰��L�ֽfY�)�����E�xR�o�	�N��޵��M���.ަ�wx;;�.��?�D���f�#���)�:�|�������.��(Gո���_�hz�c���"���4"�4~����h}L&q�d�g@=��$8�CS�DR���2��1�r�4�������jԈ�QMN�L�q'�D%1��L����gq��\m}���H'ġva%��ռ?��y�%]��ޱ�4K�Y�
�qM�2]����gg)�G������)�;�+�d�z�H
�kfu�E�3{SК�Qg��a3V�oǎ��X��Em�U�\Ω=�r�t�5���n����9Y�]I��Sͨ�.�6
K�ܑ�)Oj��}�c.h_�d�ez犼���k�N�^���ۭ`d��o�<Ѳ��I�Gt D%��^W�5k��_d/�HRZ�,�J<JE"����>�t�a�4�W!O�E��������o�;\�����{&�X���&�׉ =��NChc��~wt�L�s�g��NS����/�! >�I:��ns�Y��W[ʶq�>�k�V���\7�@��ᱳ^���v֓���. ����<g2�/���B��j>��3*ϝ�y����	l�8j�AT�b(w�u}p�e�t>�G\�֬����k�	vL��@s�+�G�	!�g�O� &l���ǯQ5�J�Mm�WÓ�k��Īr��cc�،Q$�5�Y�%x
���f�w07�M�,�#:�>�p�Q���]�d]�l�{��0���x`qaa����Ǫ�*���d:�}
�&�����9�����b���&m{�vN�m�]�D�q��f�n�=�+��I�gD�2?��ayOQ�X��aV�yɮ@��[��������\=�"F�������
r8c�V�)�K��Kn�ѧ�q��֙�s	`h���EPh�m	'�;2Y���K8�p����o�ӥ���igyz�}���}k�- E����(O��8\��Ue�ڇ�Ϻ*��A�Ҕ����v������ܲ~�!���߮�J�֙<�� �9�p���i8lN�1K�*�Hw$e�xKe���y��"?R�5����N�F�F���8[�nR��rք�u�D琠1�5Tn����I�,��<�-bsΧNU'����ߴ=�d�E	�>�������:!Fr!j�ނ�c�֞��k�;N�4�)���||#H*��H*�p����<T�(�OU+��ď&��Q�Wn%�(m�q D�Y-��z`Cl���{�]�f��h�tc�������-k��H�x�yr��Eo@]*칯U�:�J���t�v�""-p��V�yD����S�c�M���Jj�*W
4�Em�0t��{� ��̡�pm�40�K/S��"��,�֢�x-��~��Y!~��# b W�������������R| N�Fވ�aP>��i�1�R0I�v�r �2~�r�,���n��9T]���K�˹?����H
gN���4���hڥz��-R%+فE��cH�~xC7�	�z�O}���Q� �����_H�4H��`�g�'*��� 3�;��%�_����� 7D�<�[��+�N�;�9��{F��Z��7C�ې�ۜ�s~�k��f��E�s��Ύ��L��;5�6�'r�l�@n#���Ӹ�B��EL�g�/, �╟�~�z�I�,ѫ�1Xө�����"9tws�û�_H�4O^�m�N�`���{<T���r�����a�* j����x�Si�Wy��a]���C�{~���Q�/���P����A���mDa��i�½����)8��+26����񘆐'�C�Y���v�*����:�g�n�������3W�r��{�;P���٫�˻	���V~������*6���q�9�Y]��^���j�9�ݶ;�tL��G�n�Z�m�5%����~BxA�],��	E'+��J�S���0��X��������mހ|�(�K���VC�	MC�maz�,]�ֶ�YP�q��g䤹�J�h}�^�I�Mσ�~�B���D������&�+te�M��	IQ�~܍�N�?J�+5�g\�@P�� �2J�����ۛ1�����*�/�� �>�AP�ڔ`��K�R즙A�1ww2Q��OE�d�߳Sl�f$G��m�1t �������W11bul�p���+K�l�k���PZ3�E��c�&9o�P����b㦺��4?��K���%�绫x���W7�����=
 cM�Si�JOt:? .�p��hv=�L�W�隰�
�	�]�
�~O��5�,E��U%�!�m�k�o��QÙ�Mu�OX\�+�+V��hj��۫�lYE(�щ4ȶ�����_C�_"MR<8�������=�:�\�R*��J�b��G�71�bjH��X�ũ>-�ī�×�4W�h�3S�5�/�z_���JKto����>oj�5�@�߄$i����\}�H�X�]�т{�!����i�s����y:rSPڄ�[���&f\Z�k��)�q"x�=��jqv�ti-S�r9�a��&O��ݠ��WJ�� �N:W}A%�.J���*G�3Y���0ሗS#�8[V�3\)o��ɴ�����ڸ��&[
Z� ��� �pp�调Ȼ��uǳa,<��L���
cnY����Ҭ��pո�ԓW��N�#��j����=�~\Q����t��Y~� �3�,h�\���$�b�{�~V9q��1�J ���ƴ�LRF�Xc���(L�B�\Bqe�GZ1n����?��l�KBY�'��?S�w�N��`p�Q�K8W����j��$���H0C/���C"b�����l7��"���rH��>N|�5�iO����9}@駧v�{���\Ů@�'_�#�*�HR�JZL2�����n�=�Z�6��?�s��h`�;s�� ��m.6���]�n���äL;�߳Úq���W�\�:��b[��@���
�X�Q�˶��b��'o�Ra(L�C��*�GU���|[h�c�J<�M�í�M>���%<o�T����n_V;� �7yN�^�Z������]�Wp�	�>�+~f���Uq��������J�:xW���r;d�p_-�yNJd��46dՏ���_C�s��|�L�������!�1~ ���<�ͧ`/�uC���;]:�Y�	P��C���37C�և���e�Oݧ90�:���� 3�$�]\�ԭ�g��A-�!� �EY�pE���<����H���9��>G��H�l��?1�LoP���H�Ȁ�\�<P~⢊4}��|~�@
�	N�7��n��-�0
�3ݲ\خ<4"i���Z�f]���f�
!� �z�Qg���������P6��04����ަ�Ux��K�(��]s⿱=o�3@��U.Kz�R��v, ٶ��I�/�4-�r-��<���m���ͽ}��0�%]��A5� ��IG�И�m-�8f��ht$�?�"��_?��:�<
�wh㢎�������Ԕ��`����J�+���o�?�*�E��G#G���-h�6�m�ХE�{�����]��\E�-%�߿�����
��lS�E������kn��c�zĒ�2_��?;���nc��Ч��.�+>���$}�	 $�ZR�~Y�����k-�ŻMU�r�\��O/�I��N'p1�x���60U�dhP��4��Y<����Ŗ@���6b�}/��t���ܸ�f'�o6�ް��{\�T`*0B2�+��	��9�Z�n��_�p�ѣ3��K�wX��6�62�q�p���ݜǞ�濺KIL��tw\�7>���R0f}��v�̩h�`Mk�L�2r�u�*��jiƘ/J�n/�CB0>��fK��q"�jd�!��$$�FJ&���_2B�U��V麼Sef�2��xD�Q�򓆓�.f$	�e�;|EU'qd�T�A�&/K�xvx��>ɰ`�R��h�thy�w,$5]#��炏��^�e	!U����30���������q��t޲5!��qh���6��^�6�R2,U=�'ИCyM5<���j�,��IX+Z�Xu�j�`��Wŝ��}�O\]�#���2�S��ᴒZ�E��x��r�%���(��|t�O"!�G����d��[Aă�)Vƒ�R����22b����Ӽ���� ���B�:�(^3��8ŕ��șF@�{�r��J�����g�o^@��U%�{�E�4�4�?a3=֡��/�*��H�� �0�Wڋ�':�G����/F@C/��0N�w|�ɔN�`���u|^O���
��~����!>���d�>���@M%�y�����EnA��'��=AJKxM���2 ��ULf���1�w�o���o�@�&"���,�b�>�SW���p3�@�P��\ۍ}���i�u�e7���'^��ݽ@$,^�YH_Hfob*?n�&1�'�CO7�.B�E��:5��g��,�j�����������^����w�â�A�f�Q�mE _���� |�F.(x�a��b���4�e�w2!e��1������������.�����ٛ�!�1���L+ߕ����pu�����Y���L.﹍&�u2�)���K�[5�1%���F�����B
-�Q4sz{�k�8Di��O{���5�$��a���ɌV�碄ř<������dx��%�]��}H��٫�J�˞Pҏ��!S�u$)m�W���,�t������ŕ���w�o�ɺ�n'����E|_I5�@���d �~%��A"`M-�iNa���:Ǡ�h�������k��P�//�H��KE��?�		�5�Ԙ��x&d�m���#�X�w������,	��zL�Jn?��=ҽ=�����ו�� �YP������L6�-5�$l�{Y��:�V��R����%}@����K�C_�)5+<oX����"ϛ�	���\pԎ�g�Ef.c��8o�L;t�fS��G��4�^m��&(�#�xXb�����`a�vڬ�����A[]D��u�
xW�k,-��0E�<h"ѲO���h�wWƮ�\���Gφ�T ����h0>X~�e�����	�Uf�^^p��뙥�j���Y݉��ې��D�o�]IkK�4I�	����s�H�щ�򕢙��Lz�!��&J$������'�����Dm*F�����l@�����-�\�'��r��̴�Ѫ6���^�(G�Or�l�n�g��$��/r��/�0?�ڐ�ƑVm�8\�0w��DnÆ�t'M�qFC�7�'^r�jQo��8E>�u��eoP��t�+mg��C�E�����<�!w�_W�7�Lƍi]dg���W:4�ꚦ?��)mu����^Hv�|\��/.�:sF��M���h�bbu�K�c����� �Fw��f�Hܼσ~4�*"���Z��|?�^[ �6�RMLA��Ub��G�����D$�i��G�ȹ���v�{`G�c��������
�f�����z���_rZ�wܴ�����F�<^,J?b�Ks'�[���5�["�����H2�,���㘓�?ܱd.��4�>��)=��ǲF�̃�I�\���|�b�2�r�q��Z"H
h#?@
\�0(��{>��v�n\v��Q��dE��!� �s�wTG�Rٚ�R���&(l�Rm}l����yt3~�f6Z���uR�t14EAقz�-�j���du�d7���'-�?]�(����\a�Bd/@��Z~���r�yJ���"TX[��d,�}y��b���b?�2�����+~+w�m�Ue�c�|H�O�p���췒Ԣ�R�U����T8�0���"�ܽN�촑:&��o��ݎ���U/�.�C���<��L�D����?�i/�ËԳ�����S-QVJ<�3�mQ�O3"�|�v m܍�!�'��2����j����o���ʮU�k�f����.�8�Ղ}h7K���x���Um�պ���)��e,�!��(�)Oq����y�:۽>����ѐ����E&����/��G:]�����O�]Y�f}�e:R�b���i��ViaHżX��j� i(�*�ܹE��w����X	��1��9��s�iJn�:�?D3�˞�C �:7��ʩ~��\���h���0"��)���	���1��9mX�O�� eP�rwĔ4	�HX�w��?f�Z]�{�%�S�H.��I��D����j���9^Ar���\5Ȏ�>��\������K��Z�����C&��ީ������Ň��Pa��	�^�YӦ��A�5�ƌ�_8,v�^*�q��,I�Ҁ`�̃���D��<W�<�_�y����i��0R�DwiX����ɠ,/�-�k�+�o�z���S\߇tGwe����x�7@���"ዛ�Ԓ����$;�M�4�� �h����7��Nw�o� �(�F,@�<ծR�ψ>d	d���I?=`:����I�� ְ�h��O�>�
`*��6�21���ÿ��j�}��r�PS�M�v��4�!��G���m��嶏�S���ʢ�ZHX��k��V�%ҧ.����&����;_���g��p�Y�������7���H��,Ro<���MQY60"�r���s���-fZ�䉤E�<�q�&]����$*l��T��X�C�a�q��jyZ�Hj���Խ��%.~���W��٢CA��Ŧ�YR���%@����� � �����-+��������qRI����u�=� � �ё<����s��'�hO�~U�?Sګm�2�#�
3�*�(+)��.#-qD��A`�E��_�E<X�O�ɣ���&A1"{�����z�X�@��~�^=�=�����k�<+x��mE��؊��8�������Pz���<���<p��^�d66���@��^)G[�A��1�+M~�U	�N�N��>�2ݘF��+�IU�ϙ�����rjђ�h?J+�`�l�	uf�J�-��g��Ҩ�G�26:�H�X*3݁ʎ�2fk�t
�IT�CITj�R2���4�=!n
C��|�F/�^G\0���짚6���7=�9I\V:-�הe2�&���^r&�)�(��>z^�!ڑQ��2� �<��_,d(��E�C?���r��}:ҾJ���B�[���x�f�(ͪe�[Q��X����.�I���mS;�`�5��z��÷����P�y�Ƴ!���n�����12�k;U\��+���9ʅ��6�����u��LޑB)L��U����n�������><�_3��E���u�bolA��9C�mn�6�]�pq��P-)юn	�E����f����'���(���P\�~��ɽ_Ǆii0v�����Q�)hu�J�S_+�g���v����@�| Ũ������s������ݬ�����jm米k�3����p\�
ytP�F)������'�n���ѱh);����g����W=�f��O���l��\�瞩	֢&� �:&�}�ճ�����$�u^$"+�Z�x;4��5�����3�x#}��Ve��z�&P��#�;@�<�rB�8R��� S���G)�"��u�k6p��z�##�2�_~�ί����vP�]���A��3n�^�شM���ڸ���{����-(׬*��չM�7��I���܇v���d�@��E�<e�! �0�(4a��l������5�c�{����;N����̾���W�O��R�蕃�-C��]y�y�[q��3�"����	�IQ��gK�&�Q�N��Zy��"a st�'�փN��Ȭ��K7�:��YfN�i�ld=�O %a��O<:��nK�����.5u����p�Q���ʦ����H*����?`�D_�<F���[V�X`��~%'R!,��h�E���2�)�����a�֏t}����5�t��`&��F��yQm���vĊ�
�Hj��]F)BE:Œ0
�*�]��j�� ��ϖ&����w�Y���mc9zn��f��L���k����}Y�񰰞��}�B�|%��Y���'��M�G �&�H��Ο�:"q���-ƿ@�ޮS���*�/#>*�L~�/O��d-\�m�������ɸ��$���ً:�M�/,�������-i�t"�&�͗�����`�F@�ACʨ�zǎ�}�/,7���~�/�������l*"����.��}�~2_>[j�w3D����.|$,�뒧��/	�W<a°��{d�ɧCwK�޴^E���Ii�s{�Ï).o5���i_E\滤�������z��c}=]����O#a��W���e]�b���3'�J��iJIk+3�x7�¸�{E�:�b㎐���,8w�}��q�2MU,?���Z���G���uw�yߥ��_�[�Hڶ$�XE�Y����[��Uy(����5�%�h�h|�1
�6�������D�G1}��鞻�6�}dzd8g�iז��� ���(�����n|�đ��BMH��}��}��*L
*�V��v�}]�Tq����K�"ט�6�n�>ʛ��"����t�r��1���޺Ƽ@�ø�C�ښIK�.|�<��D9孲qKlX%��e�ؔ��:��Z$��d$`��W���S ��)U���S�;������Z�l`�5 7�`�5�.H�l���^�=��<f"9�H��N��?`����d���S[�������1(w�'��,tH�e���7핢 �n? ��8Z�'Oul[F�<�����#?�ܺ�.f[P)�U\���&�-�n�c�33�}������<?�I�#;FocDw�K��~=�X�E�_�=7��:����i�jE���NI��H�?K�$��R#� )���a)8��#����j-\�+��\�*a��^aDtP��t%���pM��� ���<p���ڍ�|1ܵ�Hb�r �����э�H\�;O� ��aӕ�(0�7-�`�>X�:Q�u�e>�����n���+*7��#l�U͉��Q��sl��i��/�k~�UhV���h-�*8@�kz/��Db���^��P1��؉�{xm�g�7��<�i�!���n����ʰ���j�\.�~�h���1�Am?qW��������v��
v-���fj/�U�C�}d��x�vx�h��/d�nI�qO���j�e��!�B�s,���vƗ7q�<���i�����Hc�f2��$}����Qk\h��U��n͓Q�*�y�42~�8g�������p�����큼� ���Κ��jl�K�Q�0p���)ؐ}�@k0�|}gk�8I�[����qU��l��lLhg��_�,?��O]��&�55P�T����O9��	��p�Xj	&�&?H�uF�䟌�9��ު��/�V�+�@��W����}�"O���/�P(G�U�_$U	x8�m���G���H�_��-�2���lhK���� �W��mow]6��C,�y��Δ�Z@��,�Rp�0%A��!_���{�	?'��=H�.s7��~�⍶�_t,�N��J�#^����b�U��VB#�(V_���Eo��*_���i�X���Q�w�<���a�e�Z��@����|�Y����b ���_�c�I�dJ&�B�/�7�����U�D���Bq��d,�4��I�������/�¶��c6O�v�?Ss]S�~�P�16�k�����L����1d�`��`�z*�<�A�l�yı�����"uPp�:�HF`���w�f����(t�2�G괲��ܿ�Y�4^�������`��7�긹�_*2�˭6���?��$?���Jhw1�O%Q������W�i`��0��.=���m� w�>����{�XF�S�l�`z�����)��j���2�s�����R�������}�@��v"�+��\�?U�4 ��Q1�V�B�����h�T����n�[ �l��ɜ,�w���*�h�,��0z灏 ��J,+ť�R�#�q?dZ�^����e��
y7�����q�7������%֐��ȏ�$i��X��O~��>QQ�0z{|cC�y�M�	��K�e=E3
θ�y��s���e�bia��a3}]�0�rwI�ms����hC�s����`���?�x˯�pz�6?��
/q��븫���/�;�;+�'��\�Red�\V�dGZq6W��.����p��	�$1Q{�)#J�"��O�)�|��{?��Uc,�
��D[H��s0���?
\ ڻ|=O�6��F[��H0	��qK�)5��Tt�c���ˈ�d�n ]�\�T%U�߰B@^x-��;����$�SL:I���	n�dĈb�}�����}Kg��ar4�:21��Y=�O��%��	�G ��f��8�Zw��v�\��[(yM~=}�!F��ɻ@L��5讇�&��Y>	#VR��5�sV���	u�F�G�M=$*T�Ϛ2�����LJ�S�����*"In��{�*��!��bI9����
/��J|�:�aV� ݍ��!�̈Y��B�P0��r�&�o��� ���D�&�M�U�s��I��Y�PV�pG�m����V�%].(�3�g8D�����/u��3���B�Ǟ;R�M�o\��aB��*?�$�?��xj�m����=g�Uvy��Je�ATE1E%�&e"�Sxb���U�h�%|�L}�jY�AQ��ۤ3{�<7Ƚ}������j���N����p�ї�C3�m��m�DJ���&Tt�kӀ�*5���#^@�s�k�ۚ-FN��J&F��,��Sg��`W�ԁ��x�ţ�7}O�yM���)��Bs��F�:`xʵ�"5�(+�+�$�Vda��3���P���'���[�Q�Ʒ�x�f�+�^��>W���̿]�������Ҏ��x"WL����!����3��vR&��h���h�d�s�{�=�{`��S&�_���99���;\�OM
�A�˳��+s5� P�����o���eacc�f���$��kq'Z[d���?����klX�9�B��g��6PhC���ȶz��b��M������>��cc�t�Q@����Eu�趧��{]�;��'����Cs�ȃS���-s���z���hBr���EL��oG����Z��l�����ٴ��|�b_{xp�V���M�ը���	4��Qi^G����\Xq�Q]:_�V�ee)?Q6��^�n��8MQD�q�hZy���^ k�<�_t���s�p��?��%�/�ą��m�(�<�� �
��
�[���R��cXEك��=r
J�1���ƂfqowҽC�"���r�}ʙړE���~�ak�����E�x=�2�{������D+��� �
	�"�����r�/�k3	�F��J����f�
$.�� �M!�4��㱯�/���N���+�~�uɖ���y��P�-	@CE�b�Bc=�q`��,r���_DgD���&!}j���О�`�k�+�?(�pL*P�]�P�S9�r�=�M���(Mr�'ʲ
��b�{+�8JzN�Z�2@���aE��k@���|����[3`�;0�"��H�'o8P~�����M�䠋�q6�@�z�9��8�7u�#�NI{
3xlSV�!�炁�a R?�6,�X�Π	��S�$���Ť>�"��hz����0ɔ5�ujw&,��wo�~�:A��+l���G6�`�)�)W�N��z+�'�o[ �w��'�;�1�'lL�;�1%��x�t��T��%���8O�)�q�*@VPdۯ��Aj���"�!�Y�	g�k囀� ��=P;JCS�^D���X�s�ir��e6}�c^�d�G|���8�/Bȧa�k��BO7��T���.�V�6�$��: �?h�!�s�{MV ���'o�g��+����j,��׊�� Y.��B|�J (���M��h^�%]ۯT"E<jt�fe�.�� �G�?�	�K�&�a�+�%1�+Q����ըu��1�����ĢkUr8�]�U�8��w�~+�L��V������[.����q�j�>�oF�����F�:�c� %yo�B;آy�f�$�d���A���&�55�j*ऱ�P��u�%��#n���,s�w�WQc�>`���g�^�by7��WS� W?�] hN\eV��*���5D��y �e��K"�ڜuE��� �- �ͺ����L�%b��m�.|�3el��V��F���Q��!g�lU��1�!��x�'�1wgc�Ǜ��"�ʾ,,iy~���T-cfY4%��KOn��9'�rq���0=���񮵔��C!;���R̙���vp�9o��9�ɇe��n}��y�5*����]T�,J`��<v7Q#t�P�Ʌ��>��|����O�X=��l�4�C@ь]�,j!Q[�W�?�k�3��ɡ��b2������2��^�����?�_?�ZZϑ+s@���9��a����&W�DQ[r�O�H	��-޹���:�Z���	������Py���ܪ%(ŉ֑�s�S�RCx����I�?ʐ�{����0�Y��4��.?��ژ	���'s,���]�cۣ�͉�C��	f̡�	c%��ܩ��dsoz!M��^��w�<����y@��(,�����Vă/�#K��/�N��#G�HS@n��^��w	�i�Q����!�>��Gl��I�Xm�����aI��N$���ؐW�-G"�Z�%V͆K�` sp�͗�d�(��t(�(-ӿ `1��`�%� �|Ho>|;����(�ҾKB?����tw��\�DWj6��wɀe��#�&�X��_Q�:��I��nRYk�F�V87�ڨR&_QR��IMM j�-+�����o	`f�#�oQ-��]l��h,eI$��!,#��y��R%��VH0�{=�>�ł�f�Rh,�Phv �;�K��YB�\}�e��ϐB�°4�2�" Cv�L��hQTfì�m�τ�x|h��N��{���{�c�b��=�$�,!�&���eA�؃\9:�{G��A7�c�Y���P��b�U��u�a�b&�+G���޹E0+�O^��ϛ��~|�(%a��O�h�&q�GK
E�M��0�*;��S��������`Ѥ(�Uo��S�A��Yi�q�V��9�q``�r�:`z�"���=�xYi��%n�$��4��B$��9-'I�����OBق ���ё�U��5b��ALXfFͮ!����x&e�?���(t��
5������Ȏ��/�EߖZ�J0V*1l�H�`&/P��x��p��}=�-�U�{.d?�땮��5)�C��7��rvvZMGXax+�E�e���kCJ�Q��V����z�R$N�����_K�?7�Ú�<�~����2E��`b�a����ߦ��7>vS�����V߻��F{C���x�,�l`S�l4����U��Ok�h�ae�|�l% ����h���>��Tr/��!��a����xqxw6q͖4�e:��'�F�>P��Iqm�����������v\��3����a��j3;�υ�������Hgy�'*�8��;�[z����r����"�֡���[���<�x
�@���G}>()O���g��&o���ۣ���hU?0�_��V4<�Y:�b�H������� �Txn�@��T>^Y�|�rժ��*?C��n����R9�O�����P����(���|uC.-��e�#ڀ������ ��+��tOs
�l��5�wʸ�Dv�J�qn������T��X��Ϸ�s݉B�߾"ր�d�T��z`�"w�ܩ���+����&�B���Ur`FxUX�V�f��u*OF��V�-���(b�����c �;ϼF�����\g�*��MM�3����3
ճ"��ߍ���"J�͆����	!:iӡ���{&��e��S����j�X�ג[܅54����?�5��`Wa�#n�ޗ:I�:���/�����'A�C����j��9>g��;A��َ�b�|�q�I�`��Ǔ�����)��$���ͬ2ԋq�*��^�)�.�z�w1h'�e�:�Mli!$���[|�˗\\�Grìq'\L4�Y����u�/��0�O'Z��z�ȥ���6���8�jY�qǢF�&`T�n��,�9�EzR�+p�T���X�X�_~~����l��QϾ�*���G�N���aP��|BL�6�w�x}`;�24�!=K;�ޓ�|��9�B����7{�;����y}w�)�(���j	𸇦�8g �A�Z�\hEAw�jw� � I
��M�)�?��I%˙�6�$|�� ���n�!ɀE�W�kI��_���A8�@}17��s��8Ej���b�`���csR����M8��!B���ʙ$�Pǒ���%�TZ��	�A�����|h5*�_��UC}��_X��p��'��T�8h��5�Dk��ՙi�(1��1�i^�c���DV�C�-�W���6�dΫ���~�߾���4�Ϡ�J�pg�cٽ#�E⁤X"T�"r$O&��F��w���F+��`�wJ���{GO��bD�Y�i�~R�+ �P�U����4��޵���*�)5�����)gd
����J�+�'eb	���5��E��%�jg'��`-�g=��d֥P;v���G�B��������;��[K��O��ڪ�n�o�Z��z��m��R�]wQH�󯹎�����+�f�o ��E�Ao��X�j~DD���:K��������C��|W�������V��3pC9ԋǎ�:0ev��ٱU��U�<F�Xڅn���6���͛�w�6��d�.{A�춇�&��G֫��X�d�\b:uD��*wn��o��]MG�l���
>��,2���#�(����C��S*p�5)#_�1,N�öc��wi�z-��ڳ4	�#拡x)��r��E�YIxs��_Xl�Z�3[�CÁi�ڒ���&a�i䙤_���!��s� ��E�@O:f�E��4�(�;'B�8�8�m��4ʵ%�*m`��J����x�:�� H��ʲ� ���T��K�~�����,�[L��H���B+���cV��B��9��9x�]x�!�\��:�ƚ�[�-��ܘ~Up[3�%a)�d��tI��P���) 5�X���
֙�.�h��p5**��&�(a�;ns�R����=��Xk�=�>��o�}��?N1�~�� �U�V��n4t���*��q�<r�D��pZ�ޞ���!�7�2Q�g44,���v��ʒ�#�t����3uO����4�Lr�o�M0��~�zr�S�(�o6H-�$�-}l7T6%�&,��m��/h�����QN��s\C�U�����%��v�0�!�� I: �U�x�@q�
��
+
�zH��-��(�D<��B�Z���_i�''{�^�atbQA�5�L�5I�)>��eU���l�C/�nmhηFmŊ�)n#o����H5�����o$�Â�!�;��j�@�V�`�q�����  	+�_,ɿ�z;����1eʚ�V�V�A,���f?>�{ K�����fwOH��_!���o� ���1��;)��	'z����e#��*�dX=��"�%������K����=�b�}$F�M�����C���C���U�j)���J0��{_W�p}��(r,y��W��&�ҿR�+j&�`F9ղ��S�g_R �c4����<�O�K�����ș�5���C�)]J�z4�����5��9����g�InɃ���Wj�4\�;�����#��q�ͮ��R�ੵ,b6�F����gT�	kt�=�c�v�Z1,;�a0��a8xH��g�/1U�k$�����LŚD1�s����[�4�1�D|�й'2�x��4/<�D�iʵ3�2P�ؿd�w��"W�-�<R����t6}<{�!'�[��R_��9?��*y���a��8V�H��<*�
��<f��ǭ�yTj�]P��St�ݍ��J@���}��8���D��^���6ƀBV`ꣁ$#�_z܈��83�:N%�kn5������S�8t����xZ�������O -�6u��2��d����'�d�L��OX�Ч���}K�)Jvn�,����<�4� ��r�6��_mVh�Ij��s&/:�W<��
��D���"B�GA�\�U�U}��`�B��1��S����L]�Աs���&�|ԏ�̧�8�O+��Ј�K��7�������4d�kՋ�܏�w�oZ����}O����13����^mn\^\I����j�Fb�<�b M([o%����Ȋ�T8k�E,sS�Ҏզ��������6���ЧU����ǁJ��Q��6!D޸��G��B��;V��[H����|d��J��S7��I�4>K{Ĕ����#F�#w����>���eEs����b�1�k؈9����FvmF@79&WYv��c}���@KN�^��Ae_Ҕ)�߯����Vf&z�K�z��*�Y+w�>��o��y����3w�Ⱥ�}&�����0�Gz�U9��O�H����P�F�{J�đ��,v��]��&�]��6�a5�x݌;ѪIR`7��!_���!����]q�����ѩ��d�M�ou��`,���� �a�L|d�����E��c�KZc0��!&���&z�pS�|���*�#�2+�N�#|o�5)c�m/��%r{�l�:���Qյ�K]}��>�z���r���&�́8��р���c�
��B�GѦ�V!���C-��3�IYB��t��T�/��#��Sȁw-��7�#�A͒"�8�%�F 9�VUb�=��3~>�O�l^W�E�ԥ@��][7H��r6@��dnQo%�䛘�TMM-��ңυ�+�~[L��o��? ������3��]�m~���?��>l�=+9{y��I?��e̟
��>I�|�}�FG���~U8�?�y{�C��M�% yf���y�����1��/�(�̀���+B���>�'6&��b�D��I���25p0d	����.���qk�1z4�����W8�?��Gx6-��J��ix�����52Vt�y�S9� x�{�H`s�Av�u!}��),<�X�XV�T ppC� |���<c�jQ���=۟���ǐVA[;6���h�֗*�����He����>�{Xu��G Ayw��N�=�:x�dj�=0a>��M������@�R �r��M7�2��K3��?�652Id�ՠA ��Kv|����q���w����7���?=�Wq�S�Yĝ+�7�̾�v^�����xNBR�8c��)]��ʀ�B�����s��{�/�xzSv���Ri��'z״u�r�����M�����K+��H�df݈G���?���n՜(9d�u&���M��Q�"�Ͽq��c�[���Q|�x�+�k=�
ݕVL��ц)��@����pCm�s���� l�E(�%k\�5��v>�1����H��<��cR0CQDwOHw�/~�:�V����6�ؼ J��)D��	�eIJ��8}��V��o�ZQ�NA��։VZdK9�ˋ��N?)J˅��cc����$O@�ܨ����G𸊳��!�'�jO� �g[��uG��*��p���;x�n�v�bn��6-�b��?���H�bJy��|>|ŏ��	L�v*�h�be.�w?eH]�eZ�M;c� ij��V��w���$U�,��g[�^5��]
Ш���UL���*��o]�UcuU���d'I���b<���t�N�Ab;%�{�Q&���a��;��g&�k�r��z7��W��_V#=�Yh��>'f���~$}��#����O7��_�������۾�xM�N���b1��BJ@�����`�A�hA->?i�v����l���^KT}���)��
:` ��X��î_��轷* �G��葇�Oҙ?�:�Ǳ�6��K۾U� ҉��)-2|B�O'�;�k ��b�M�"D{� j6%*�IdC*�Q�8�/x����A�r�b����SDN�
����ȥ�Ƙi��ˆ(%� ~i�}�wgY���U~����_���������H�%ә.s���p5=Ʈb]��-I�Z���}z��/��{����+����?# ����B�wJ9X��ܼ��h29�4�{yw�^��E*�J9�k���eԓ f�tL�A.R4�J󦦬.�����V�W���u8��4+=�1ڸƼ�l6����PMv�O,儹Q�����D��i\�>����N?�����V8�m�)}O�aK�����7G�'�+9�D�&>�({p�G����B ��,#�D�i`���q�]|c������F��Y�k�ׁ��f6���^�TO�?�.�l�\�u����Oh���R�[L>͐��0e�����xu�0ͤ�Z�5�+I� �.�ʰ$P�0@Y}"@���ź�B��tK\R�]����g�ya�Q�����/�86{{��,�IJ|m4z�m�v�y�r��c�^�l ���H�����?�������p�Ƿ�@��([�ġ�^����ǘ}�y6��2xҸ��?#�J��a���~w_�K�r���d嵼3�W���|�ۧ�+K�#�*4@�
�9�e"�t���7��!@L�̰�T���fD}7C�z��(�Ӝ#�-��3���p�3�8�?���e0�$� $G�x�!��.���~v��Ў-�������n���{@�F|>	 ��s�W�w\�OThI�m�����>C�Gx�[u,i�^���m�oմ)SY�]~��ڣ��BKJᾫ+�.W�o��*p��M��n�&^L{@=���ё~��+L��V �� cxn��OK{��<����*�fۀ �٭��������ۧǫ���l*�cgX��y��CSi�;&������N��k�J����.�ƤL��H^X�NM������Ƥ�(22�K�iV %�D�RC{��ȉ#�оnfB�=T(�X����5���Q�TH��9D��")�:�Я�{ث� �懨�p:�J��Q暕
p��KO�(��~���6_�t��R�8��4}zL�Xb7Jq?_p;|��>"	�|�%re$O����)(h<R���tN��CA�������9N������\f�T�q��8�^���}��5CH�ȵ5d��F���yRq���=�_�x�<����]?�ԥ�d�x��%��Z�q8[��a]q���E3zJ���O��됹�}Z�����r|T���%ܕ�����3Cu�]��i����g����rc �Ym
�8{� -�0:�b&�-�