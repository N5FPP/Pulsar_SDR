��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY�y��[��Hm�Ȼ|O:N!�W������w��5o!�N� ��7�Ѧ�9X?��E�ȏ��S�nI��F�@C��j�W��	�i���q� ��`��������c�Rp�T�N`u��/�#��<��#v�,�.��.�~6���ţrI1��"���R}׉d8�����gX��}ɡ�{��S~Z�Թ�f<u  ����tO���D�h��_Ձ�R*^�>V�	2������"��"��<@��\������� "1*�� ��U�s��/��.����`f%����:�A_H:�C�k��JC��f���
�׸��
�)���n:�uѮ�$��;w��l����s��v8\Ð�F�"@�e���$�L�^H�+H�����I�*�཭U°�7=l�H��Fl)�v�k��i�!q�No"�.s���`��wr~-O�"| R��m͝f�A���R~m�8#���]�_�V�W�,g�BaFA��^�j�� JwR��$�\�`��'h*�Ȋʽb���%rn��a!�@����{���ʑ�h?H��&Y�e����W6��gV����� �)�w$;c�kV V�|���X1��~�=�{���hƍ�}Ȳ�}D��0,��{��""k<�Y�����]�#!`y�~"T�����=�э�l,���α��Æ�9U��Ỽ�kk�\�En��5�"��l��Z��1�������9�H6���97(X����ɋ���8�-n�L�kG�@5�~��g�g�|�ѥ�%�c�ո˥�Ev�h6d�z�K�|;?�{I(2�AL��AQP�q��rOC
���<��M�e�t���
���˘@�R�}F2�<�Pd
OO4%<R�a���Fg�M�>�ſ��X$"�<�셢S��I�8E1�^��5�U�Ñ$���u�u~J�`�rF�C�����[�l�u�I��xv�S>w�y4g��T�>O��I�����<n��P�����p���lOH?U4�d��UL$��5��?��0��J�v�r]� ��L�vP�B�3*1�>����D�ʷ��{�Q�n9\��U@6��3�e���'Xk��|�&2��Ļ!���Ky��0�Ն䧏��Y�>9): ��{'޹k�v�Z���*�/yIc���1�$��������>[hI�
~'�Zm��α}�?+nx�̌����i�z��j�ܛܯB���̗c
�#���j9J�g(��/�#��_�Q�P��Fr��ێR �;�r�1G�ì?�倽L <G��,聰�Hj�g���R���A���H��:�1̳�/�(Ua}[����{��(�"�d�Â�>����^8�Y0�T��;��nN6z��uv�B�����Ɣ3��6�&T��3-m��|���L})��˭ӿ�1�Y+\�?3�@��m)�8����|�PO�����1��|��
Z�A8���T�8�̩�?_��d�'�;�̳�
�оi�G�0��F���4�b �.TG�@_\h%�'�'�kM���f-��`�4��s&�4��T�͙}�z�RնI��z�Ek쥦Z`&^5�Co]��)M#r�e�TpxTA�#��|d37Xr��*v�VSӖ TX�J�9�g�uz��3����+<�k��_�_��}_�;7��k�&��~޷��J_���ۚ��R�8\:v�m�Q�h긎��*p�7*�"�{(��*��2kfd�񿆨N�&�6\f��> @aq<H!�b��r��K���3�2���a�A�/KG��"|%zJuω�m����j�e�"T��㒒,D�䁀r��}�q�����̅������m�s� ?�{���gZu5���R��4 �-Y3F^n���*�/��CDs�.=�7���Ң]&�:%
.�nh�W�G �Y ��`cއ�;U�g��f��)�oAmq.+���rZ��?�~��(;�R��������_��ԗ��[7J��@P���\�vR���ҭnG}G\�D�f#�o����>�ﯴqr-#��2��F���9��.��F����]�GFΘ8���ZM̃���汾��!�?��)"��7��W
�
ZH4����V�bR��o�����#��K�0<��� ����b��͡w˲vI�ٛq$PC�5
kV�����&�Zm�O?�>����3�#�H��)F�A�������&�a�w4gE',4��y~��b�� b�(��>-���>��V(/�J�i��Ng�)oCȼ���}�h⯾�&�R�7BDg�f�x����3����*<
����~a���۫ o,DV����g�=5r/��6둢�m,��OL�|cg��;��N�F��@��0Vj[������t��Z��(�,���w��D�F�7Gӊ�&����.�oGcy�i��	��P�c
 '���}�;<����׈�Lf����~_8Ƅ�㳅������g�G&���%AzH<5��FcC�"�qr�0Á����_(Q4��v�q�-�h�@�}{��+F��Y߼2��ޥ��?b��� W�~��X�ߢ0�^<ٮcy7�DC�`��ϴ�fU>¢T�+~la-n![�p�~�,��/�4�� �Bgg࿼q��Y��1~�Ќ����PQ���>���]�a�w�dqg`V�\�R	�(t��8��B�;�10~"�� @���Wu4M��[$h���y��K6�g~z��T7�M=i��l��f�<�=t�����!�`Z��U�k.�#����M�E�02��q�0^���{Eؐԯ@�0�<��5�%�	��A�5Bej&���E&��s�	�%k��Z�U�t���%t`�"5(��Ϋ<N�Ȑf�EӆاB�ol�6��fїYsc���b%�;3%���8�W�~F_(�Ϗ��O7�ХJ���� H}��XV�ѻ;e�@B.l�̾��@��&��/��E3�85�:�o��!�R��Sm}�{(�׻8Z�<�;E�J;�čy�'��~���'��5�A8�1yL�$�ԯϧ���s��oTk>�HE�QĘ��R��� ��1d��>x�RV�T�T
�@�Xϡ#�o�M���BH��MDǛ�)������`�X��\�+�N�������/D&��U�,��ˬr�f�)�sF_ܹ�j�p�-/C����)��bX�ܕi�a�DH�Zl�̔�Wò�7�E���E�%�}T�a�&��Ռ��]������:;-���UiN���N���b�D���7Ik��G*�L�(UfO�6]g��׽:�,�y�Q� nn�:�ʕ�T	`u�٥U]�|��0�wY��u��pO�C�^�*X��G��I����q�����:��YW=�1(;3��ߛj��i�~%�.��wС�u�/��W��*;�#cH�}l�{?ըaŤ�\k����`Q���[��� �|��H<H�h����[
���8�^LP�O�|� �DA������xb	��g��Y���*��"B���|v�{&#�<&q:��%]�i�Ͻ>jIV�f��ː��q.�`��v�bC���)�.�O�u�X�����^�Y-y�]��,�ŜM�V��&�d0��N�yę�0t[�\�ja�����k�K.]���
��&b40����������< Ա/��ߞI4��j�Ӡ`V,�b{��*�_Dƞ�o�qT�ԍ��ȳf�LQ 	�Wq#�&}O��ү���nxqV�x�+dN9yf�&�lÌ��R�iG�Ѻ9Kϰ�Kw:ْw�7�S?k���(^�׮�����Q-�.��s��$�`g�6Ҵ�DJ���P�����qM=TyZVh��ПGv�[�!�"�"�-���|m��mp�H��J�����^��-p������Z(0�H��{B����`����͡0�q��N��������i1�H�iW�!�p��!�Z���b�;:����"iַ��f���d�ٯ&���z�L�-C;k*�{�i���߹v:�~��R��D) B�#��>+�~`�3����b]OKZ<�X|���5
� %��A�=ߦ�d��f2��8��&�8n����;�	�͈��UÔ<��Ԯ�ء\Ů_[���0�)�L[-������u�wQ�����f�K����p�5:�}/7 ��H�&���Qz��e�?s*�M�s���1�����mW	����_��QՆT�A7� Ya�L��g��8QG|��2ľt�ff�й�ĸ�;�� ~�Շ���/�%�^Z���YyK�����!O�ВfS�8�Q�es*�{TIϮ�U��:\�4�% K�
�~�gV������3�u����� �>@A�%�Rli��`�%��XLi#���%����R1ܧ�`i�%�
��ߊ9��Ɨ�t�Pd(1g�R��)�
q�:�I����е�?\T��b	�@���F� ���}�̫���\M�;�v�?���e�Ҕ}������Jd�7��w�]�+8R�@KY�%On�CD� ���rj������#d�Ȯ�m+8���p܎�t�f��J��R�xR�T�"��.��h�L�^y��|�PU�c�ڝ��?̋G���F��c�Bm�V)�0h�-�����3�x��X�],�z�8��`~�r�^[z�UȆ�����#�L����Д�CL�?O�$�7I4t�/F��}zr$a3�
�;&� ץ�7�:�!����@�������<\	~Ԅ�?;��H�s(���ʄ嗕=F�C��?��]
%ϐ����M��Bʰ�1s��G#>�"^쿕�α�����$�rg�-�rO4y���9c�0�a���+B�E'��6؉��]L����5jTIy�9�����%�둂���t���VBN�= p��.�Z��x�w���ۨ:�'5~=[y�K%
��$�⸼���)`��d����i�wl��(P�@�"]�\�\���5�c	�06&��������X���CK���u��~D@��o�����hͰ�.��|��\����EAG�kɧ�|b�<���p��s�>Gc�,�ށ�5�΄�{g[,��"������,C;�QZ}o]^�8L�$b�dM� \q
���$w�6/�lHEu�����;�p �X�ː���8N\�,��P�;��{K
��PN�����������ޱ�l��iJ����顄���l��˞�����d`[�Z��a��������?��$�1��C�V/��R2����	���Z�RV��$q?6�kŵ[H�����em
Cp2�s��v�Î)R~mR����WL�c�㩵zkr�!�2cZA��iq}�C=���/<�	���^39AD4h-��z�)��HO[��rȆ;����1d{�c�(�U�)�cZU�Rz��@���h������k��C�9O��QωK&�
��m>�̰�]|59�BfD����xKӰץ|��L�����Ǝn:m�Ҙ`7��NjY�Zԩ��D����֥�� w�N��Y��W�?Px���4 ��Z�@�|*��{� a��)=n7��e���SmV�y;:�`���)�NZ��ګ~�[���������]6��8~cM����Q��b�<c�l��-���}���2��/�Z0v�S>� o�,_zIA��`���\T`"����Б�Q��.CHY�M.y!;�;�20��D�A�m,� :��)d��᭵ �|�͉Q�#�qd����V����ikO;���e��-V��>��a�w;Âw��Ӥ��v����^��E��z�n�_F���3n�O�����wQ�������8��@����
m?���u�Rr�؛�&�"�x(� d`oAG��w�`��mM$�����x�'�0�b�j���Ul#l?fQ��}�HK�/�ų�-MC<fz�s':T�P�E�Aԯ�_uH��r�}7Fǡh$+�}O��C��2��x��%����|�4st���"ʬ�
�ea�C��)�H^�u�3Cl�5������
�����I</j_�Ә��,����q���#p��o3���(�fjQ�ͤ���)_��Q�QJ�X��y	mHT.�I�s�������������e2KzS���mF'������� ȫ��{�c<�#p'���I�oaI�&u��;����Zp�UJe�k�����y=�������U������v%r
�F��Dl5,�z�
��:�*�ONT�Hx��_��~D�;���ǫ4y���9���7�,uT_� �`�FȪ�J��7�^��#��w��Lx4[|cX�С��`\�-y��t�HB6R��R	��{�_Α��؄��=�V���כ���9��hј����{ɫ�o���-���Ǟ���R\�/�Vi݇$��߅��?����
�y�^;�����a�I�lxu�:3�`��+�������QE��}�ݠ�����ʼ9���Uǜ?��\�M_�F���Ʈ� Q�8!�����s%P&���"zP%�@C��O�V�Hv~m
���y��=��cX
j���S[�` *�o���� �}x�,�=�q4h�Cq/�|�"/U�c�c�1��c�6�v'�3��` wn$O�)B�W
>�17�����C{�=��$���IR��FL.T�;O���>�ߎ:N���P�!��F~�?h��e�1��Tԍ��|�(�0�jlN�s����WM�&�
�W��G�����g�į2�0��qM1��M/���"G��AdqC���ZL*��:Q���J@?~�o����	�7�hx�w�:|tp���t�k]gW��)e�<�����=eҺ�rf��f���#0�����Bsb)"����fU3k(�2��e���u�ۏ ��.��E�!���Q���"�9[,�b���T�xBn8�U�����+����H�!a80�;��1�h�����,~��b��q�<����)"<���������?��'� @�}-_'7����6�:���V�S䦲����sK�<�ꈦ?�̅�o���K���^��P�e� �b�9w�z�P���1(r�w���<��t/�>-�9e0�����s �ʀW���"��Q!��������=�S�)���y��}��)R�Ǆ/'[7ͮ�M�(�#�æ�H���U;+l�ud����\Eb��	0��v`�Y|q�4�GT�}B��a���<��U>�o����N�� ���v��V��|�X�?�k���Չ�,񜛓�b��-q�c�b�gW��|��6ZP���k\���e��*e�K�n�nE�6�E���Z�5�3�N��R ��&��;k��[+��P)(�~]���j�+�-�G�ж���؇�|�(���P*��{7�e�f4U����9+��]�����m�X�J36c�/����>�^8�8��*�ƫ�$PdE+����(�W ����Iٟ�wTI�Y����:��eM!>��E��1��`�7]���Mѻk�_�(��jƙ�H��d�WH=ұwf��A����4HP���x���0�����l`!G*.��B�(�سoz���aE�sȽ��.e����H�L����-I)A���ONG�)�����h�W��~C���{�����mU:�[-D8=fo�S?k=�M&8+ӵ����t�������ɂ���EBhӻI��A ��7Uv��o�v+�fJ� ���k\����D�S�������H������zK��UMU��Sq|k�9���7�\X������(�1i�bm�x��i���GH�`0�a�n�O�v��Jݎ+߭;�y�<d���2׬��/+^j�/ՃQ}�U�����qn��8(�{Ah_�S����ҍ���Q��H�lQ���}5�ą�V1�?�5�U�M}��y�s�[�%L�q�����H�?���i>?�ҳ��]'���{|'||��taa��?FA�/�"�v}r�d+���R�Oͥ�`�ڿ�:���b�\0(7C�<�G2������n$�swgT����'�
��J�I��`N!8x�N�����r_ܤ+�RӪ��l�6�������-q��3�;繹��aO��m�cx	���ӯ���G2�2�����"}�c��)>�7�S�Ƃ�E��U�	����O#�J�����&,+��t�L�����e7If���G���PQ����PJ|�abE�*%Pca�_2$��O�Z������8��3.�A�<K`D�򇸌����*�C�j�q�D�iV�S��=�e�˵$�/iV]�A��r�+�D��6-a�盶���ju�Rf�4��w	�'ț���Ȩ�A���r1���N[Z�U�I���� �����Q=���&̀͝���T��}���TW?��?� h=l�5�?�������r�DKZ�
�����!�[�ݝDV
K��>��fu�ul����>ʾ�CFC�W���-��v����	�,ޡ�����FɚS��(ya�5Fx���4���=7R7&�7��)�%�~nM� \<�h)����7�+�܃���败$���_ش0�Izhܴ���S�@�/�uROƆ��>���LI*��~�Wm% K�Ք�8&�p}�0DZ� �lF��GM�g
L�1� XO���C�y�]2�3"]�,t��^-%"4i��s��TK�eAԠً�����q�N��}�V��&�IX�"���qR���)D\uN�Hj�f���s�&|��E O���|�
)Q{B��>,��d����֚����k���s
tg?|_nr�U>XP���x�*�܌��Vm��]�M�;�V��}j2��<\�0wN�\0�������y�D�TJ�ɕ�,���\2��;Xz ��Ϭ&��f��"t���N��Gٴ��(��=�#u�0)<r��'C��̢�qO����������H�$��#����%�x��u";�d�J�0����6���
{����jj��7LO������D����{ő�@�&��Ƈ�(Pz������JCmp⑂#�#�$5�M�̯#Jc���.�}Z�^c�� �F)����+~~4���^���[h�&h��U�#��V��0��b�-"3����LaG6�"hÆ ���$�\�d� �K�)315ҴQ�B�#�68
:<��n
�T�_�Zip�d�Z#��Ǳ}�$�qWD"ϧ���7��,r��	F��-_z�kI�E&ڥ�ό�5����c,y��L�B��5|h�-L�5���������)��c��L�T�=6�@�`6TN4���gv�*��|En� Z�v\4Pz%��=.D��똫��b�M�|V�1�B�	�>��dn:���-�n
���d���w�r6�&���E�IL�X�F�4��'�'�'ZU�8G��k xX�}Z`�e�~�q,Pmэa[#RMG涼�� We� nȞ����CN)��f��%u�t�ON?�WO��K�L���j�[�ʀ�0���=I����s��U���x�_,��Wj~�������  �ho=�Ѝ�^�>R�n_�S.�is,�% _/˞9Y8|$�s�r�dm'Vw���.��z\�
By~���%� (�Ӂ�uд����t��C%�Ua/�$���O�̊���9e�o����:��ٽ�J�F�ֶ\�߈^t���%]���%�u��n��sW=����]8�a;}��Y�����hN$�w�u¯E�� �BN.���3R�Y�+@)��.$iR˕��o}���T&ݶqa��+ا0��6$:J1f�Ql�Hi��o����i�w5__��(��y*���_�%4�� Ӿ�E��51����7���S�;��K��G|ya�MF|�R�ck;5���ЄѷY��L��'y��q�1��`@KY��f��݌����v�e��w�2����\ؤQӉ�u;w��(��?bW����;�TT��GUx�@���Q�K�8�2R��rH�|�qu.3R[y"^V�Q�q4�t44�|?!}3İx�����6ƍ��뮴�"�*�@>�P�'N�)�-�fXA�����4����a\�a�؛l
����j׏��~z��S.hH��[����QE�(�Uvk��R�64X2��X�O���dO���׏x��x�NF�I�3ҢϠ>��s3SϹ���S��Rf�~A��9R:��چ-	УZ:^��T8��1�Mʼ<f�w�pe_�|Зǉ�1l�b.N달��*$���r����j�X�T-Ͱf/�q���N�x�Y����6�.�C�D{qK��[>wEt��ݴ�c�ggyL�����3
��>�m+�T��̑��~�&BS 5��.�j5G�޵2=l�M�$���;�9��J���֦_��[�2,�箢�He����y�@llvM��'
J��V��KP��:|"ΪS�}�i�^a�z5��\C��Y])'����6��#�g���p��|��1 M�v�;�ؤop�@(d�0�9-V'��?�cƃkL�W7iس[^i�l�>q����,!c���
(b@�|s�+Ƣ�(���?�:R���n_�L��6��2]N�$çB��Nב�W���;/��A+�{s7�t�=<sD�(�<�����Ռ��p`㲟�������x����{!�2�ܸ(���-���_���*>�y�mAU��Cq�.Sc�Gq:�y�-�u��^.h�A-�)�����E�:��A	�Rۙ��E,0=&��qEs���xn.*g�K>�+���ܪҧ��5B��{k��`C�xӆ�2FE7-<5���6�Hf>��b9��]$܌vv�c��`���S��1B��[��d����i8��f�����m�[��?ۯЕ��D�qI�����Wc�!�v��2`�Ti��XB����a1��%���h3�a��v|��8*�6$�-��d��s,�ޖEƧL s�vN�Nz�za�5�@�FS2$ �������e��P�!^A�F���v y�H�������Uj���������q�O��ЏRh�j[Őt?A�{��F[{��|�uqô#j��־�[Z����M�F7T�$�9?7����pu�,�nS42+_�k�S8�[Z 9U������y_���:ל���E���9�Ы~�Y�O��ֆ�e��&�f��S�� ���«�\���"���
�.�5�Q�p
W?)-
�2(�YO�1��H�o�a��<��S~b�̑���_�?�tP��1����f�k8�w�d��2N�A�N�~j�L(K��g���z��*\�[�6�\X�2e�������
n���Ij��]s����ӫS���R��󆖫�W��3����\�L����(�#1��؃�e��!"vL&�-��ł�s�v�Tm�V����n�j>��ݣ��4�M�8YI�b������*�*�.Ă�qf��6��E�LX �]
0Z��r{�{=_������a���+�?���z�v�t���L~RU{�K������h� �%�qbU&+J��J�(��ͩ4�������^ =4_��y~:r��	*�/�ް�J�у�	�N�Ip��FJ�G��9���l9h��	�d'