��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�۫k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α��wԊ�6�a�3� G��λ�:~7 !�v sh��~��P�'|#��x�C�[�~���{-چ��!�:���)�#aE�C�;� ���&�'��c�w|�:�)��$��Sއ�Y�K��N�4uFLN��6n���)G�Kh\��V�A2�� �@ͽ^+ϓ��zm������/]>�b�_=��R(t<��1���M�kt�Z���u�m>�����R~9z�x�N������7���x>��%h�>v� ag w)��X�lv��?�)����������߭�n7�<ü4I��c���V��"�TE��Η��7E4�#��+t��w����G�\΃�&,6�Lzlƽu��i�����#%qwVL����(��d��\�(��E��?�֧Y�՗P.zt=�Lل�C9a��t�!_�n�ŎCi�o�^&ve���P�%�����Qo���$���n� $�zXSQ�.��y�X�C`ә�!>�3W�0"��hx��؋�@ kD���LԴ��)������>���k]��h���di���������3b�g����R�:EP����'�x`��Hn��Ƕ���x�b,��g��>���Q�ꚡJ��� �hA���ˮ0;�Ǝ��(x�PH�wXG.�Jr��oˉ�7�k�u�fC{�22�uneɂ�[N�7
��Y�T��R��>-k���	ٿ|��%V����ƫ����@:�J�F}�7x���ABF��4�� *����.�R��^�C<@ =Ⱦ�Ď0�8�X	4s���a�E'\ٕ/(�M��į�d��3]�8�����={�M�"���[�=6���8��_+�����CZDc���iO�U�`-(h}L��}w�wN,��kx�a�2��b�$���j��Fq$[C/�kv�:ҽ��CTES�i��F��b������_�,L� �7	�r�OC��'x�k�]3�P�P4ei�� �MU�^M�kuࡲ�{�!�)���뙛�9�8�M�ZpHc���PN|��Ȥ/k��3�D$R�)��N���C1te�0��f,G�|%?�F��!X�_���ӗA}��ք�M�:����;��L����ܓ�חUp���Q��$��$�d�Ť)Cd�r$��tyE�kC��x'ǫ�J�y{��q�2ay���ة%y��r�}����U,�mc]!�')�.��uloZг�0� �lW�+Qo�&�8�Z$u�7-j� �����ڄ���<��S�Kׁ=%��n Z��4 ���*i֗�{��/�[�䤲I�%{�XT�X�+,�������H2է�����$��*E4��������Z���}�ޜ��?��#z=	��'fU�(-v�gj��WJ?�0Ce���E���?&�kM�=����mj�tE	�3׈�\�h���+�1z����'L4��W�V���,� ����rWV�v3���f�p���Js�@�$W=��1T#/|d��v!|�$���Ѹ	��,7�|�i��b�LH
E^�U����9��*�릋��~�[��_G�$"1��{7�����H�ϡ�͏{�����[!6��X�8x�e��6K;��+.��z@)='=�c^���W��v8��5o���Ty�!ǩ�i��pD��}y_�0c��c�9�}�;d6׼X���V�Vx����Ā�1pM�,Ú�l@���0:�Ig��_�;���E-�|�>d�f��mlߘ��8а,P��A<ۨe1Y33�$��Z��F�ݰ��a���S)���ȣ�
��)H�̾�EQ��A��$�V��e�����>�}[S��v�]k��f��&�u�KS���~`4qi���*��h>�P�L��{M	Tz�@����=`�B߃�M���B�YZV�(�ǖP��α6Y�B�kTo������9v$Z���i�2B�q��2d�������,_��Vl�D��V��օos���-��x�b`3��AX)�Lb��N��k�L������M�������A�Tw}���E}E0 �{��:T��<q��3,b�VOJ�X�	Ѕu]x��C�{i����
����*`e8h�Dr�q�sG���2�6\��V:��]�Z��V���W�J���=��%�BE�����m@�ZB��2���� ,ۻ6t=dG�(,�[I�P�۝e��:���V�yB"�{�w�\Ƽ�.�����3�4r�b���;�]�`^R>y������Z�~.�}�U�)K��z)���
����dM
6!��[��?��߹���i-�����&��W�1ʇ���`"|�U���I��i(=�jץ`ܧ���*�|�>�8��#Kh�6܊� �����/ݐ���e�P�E_܂�nƠ�3&�ӏ�"��.���ȶ0��𓽭�`���V�w�r��}j@�'~E�3��
h�*��iL[�q�g���h�TG@�
q��H�~�X�|��;������Z��"s�4q�~y�"_��E�g&��*����c�?+zh�Փ~�
�}�8������/DЌ�ߑU,����d[B�z�4T���h�@�\�W���..h��7rn+e�O{`�R�$��4�ZZ�S��}�(� W�H�|2�~�I��E��t���y��\�Mz� �a��YQ��&:�e-who �f��p��)LԨ7S��A���$�1�u�S�f�'�
��dMC/��t	5��`��nn�)��H��ʹKs�O(�7.Х��@������S�!��|)�^FM� �Z�}���S;�쫰 @����v�]���>C�چ�a���cwP�b���L�ՔOy�U��G�UF������of�܇{G�
0ùϦ�bS_7j^�]!�p�dW%�K)����	E�/J@�=�&���n�f������5�����9���F՗@��
�P�j+�,��������Un�(\�XO��k,�q�ɬ �B�]�~�5��@�::b�-�`@�����r|�v{����Vq#��vK&H�p�-U�6���۰No�t��f�O_iJ�]5���e����C����;O	�	��3D �����I�`O�h]�F������ ��W�7P�eǪ