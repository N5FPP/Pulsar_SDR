��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY1�ii=?B���X��� Qj���M�1��w{y�F�	|(36#���mT�L����o������I>9jĎI�8l�i���P!����Sx~����� �k%�v7\�S�~�s���W���Y����a�x��@ ���o�[����?�h�ʏvX#PGL��X��\�9yN��������DM���JpFa$���E9I%
�I����5K���b��5�+� M���(VL�5j^�<��5��"��%��������1�0Z��3܍7�@i����<��q��}߀e�{�8�`ͥyFJ<n�>˱"��Q<,R��fa��3�}�����6(�h�*Om
�| T�Vڜ����A7m����� �����R�sh�߻���9;IM}tCL��w)L�3��m��v`�v����Ya���_��c�->�)DS�<}d��J�3�'���u�+���ٙ`ݪ�!:�y�`�z��i\9��H5��J�t&�dO�f����is=WS�������ű�9?��>�\��uВ�l�����,s����q��4;��$�� ��b&���YSZ�bDq��]��_�~\0��0�$�Z������6O����͸�GƟd%���(�}=b;�6����=zG�)]C�Q�	�Y��X"[�=���u�R��$��%^"Um�`S��̂.XNp�y�t
c�ϲ�u�R�u�ȝK4��E%B�kH���3�
�����j[�& � �'ۍķ�	s�J�bJ���ýy��J!�8Xɩ�\>5�����7V�l�4h�Js��k����@�lQc�������}cJ���}�'�Y�{ҏ� ,�����PI���T�qVp��2x����^��X�猪V��$�O]\UzR�'��x����Cn��%��	��ؘv�M�=�H����F򙔗��Kg��xG���EGO�p�P�����`j�L��;Z�M��6)�M��&���FPL�c�9RYz��s��H�hN�V�I�A��P!!w�J����2���Za4�_���V�/�v|��H�z��?� ����:i���
�Ҹ	&w8jK��
�b]�|��`<��:�2���G��'��W2!#�t��N�J�`�\��f����<8�bL,�R�y!�22��?|Q<O,Z9|no*�5��"���4�b�7���.��[	�I�u��YEK�I x*"�?<�p{�%hh#�&d1]t���%gU�Xu���%�6��3�h*�~;�f�v��
-u �EY���Py��l�	�y�t��S��珺.MUN]�E�W�u�� N���\"�!�R�(&�1#��nM,�è%����X�ـk�nq]��9���˽��@��ohS��2.^�A�x�����;�_�+Q|P�)�����=�ES՟���`x{�ݶ9��2Ґ����4K�� ��/.��_��k����ya��E�F�q ��_�F|�[��2�\P�a����o_������?���0��@�_����wG#0�NFhy�U�*�F.�3:�j�|�[����h�o�e"r�:���Lc6Y����6}4V\$�������M�:B�ּH5@:c�7Q�������>�Ƥ������/�y8!b�cQ:���Dr����Ƙc��ZTg$�]$�����~��͈X��㌾��T<��H�S�%_������E���G�Ja��GJQ����?h�� W��� �����/1������x�`A����]�1�~�wp6���R�w�!\�16 �e�����f]���U��J y� �mI��r������2��a⑇��(\���~a3��pv���я��*��5T��	a;ɔ.^�q *5�xɯ��s����ތ�Zmm��Vhy��m�����A�/�cڂ.@D�}Si�{ ��͍nx���%�d�g�Q������Ĵ �TՏ�\i��
��)��mc8+ $�u�gN�˪Z�N�SǪc{\��1R�u�j!�T�;��;hh���⌤tnoĭ9y���@�>�Z�8��%�g`7M2(1�Xe2�?�|��~PS'�V��B�9�H�:�8P���΂X\���У�\��Q�H;�>�a�@f���� Y>c�;{q�*H�"�譟���8�^��/�,mb��-yz����G�DV�wu=�V����D��Hm����o�����C�	]�.��U���
�� vT*��w�n��#�@�|���$�"�nr���s|���$���f�{Z
�>Ⱦuμ{rʔ�8�#����Y�HcF����c�-W�Zċm(Ɵ�ΔsC7��[alZ���?�U{�Z]��N�J��_A4r\:�r���?���Y�'b��Q�GRm�'G$�R�i~������#�2$�
~��XF,C���}��W5�H��ЅN�觺}*MX�pm����L!�=L����ä��<MH��?�;��G�C�xG_-����F��[ �ǥ!@m��*J�m�g%�"S54�V۪�&�J(f���H@���d?L�5�r.u�[�g>�4�3Z5.���%`Qf�|�Y�W��8C�:�Ψy?5ٮ[��7�C��i$�PY��%E�)��
��rj�/�+��\�.�m�Pr5�p����J+d� �'��"�W�V�����s��k{���t�|��Հ��SɚJ�� �Z׀�+�v��t��[�u�Vy(���҈Z ��I����+��ȗ���J G)�bt#FY�-�6�!�������J+��gZY�ӣ<��~ �����X�t��Z��U4�ݵFؓ�÷�(��~��m�٠m���-7����og0�xCd������}_ͦ�i��/s��<�
	�/,��Q2~I1�A�����/קsT��X+��e���0���a�Ίh���P��yM/�@�'z_X<|L�Y��*)�{��}t4��op�8���V�e�W�*��$�݃7�=��Ph�a�v��s�aP�j�6�ZC/��g���fpa�,&�߅���yr�mL�v�ذ,P<EO�Tl�p��t������i�ݱF��35�{1�#�I��W�^��=5���Q��.*�RJ��=2��;|���h�x�E�P�q�����V��=�7��P�q��V�]�k�G�Q_
q�H7xZZ-���$����?:w���p���)�h"�#�q�y+��*x�j�`,��9��Xm�3��n�D�!cx�	pX��^������gVҶM�|ػ@��DK՘���Ի��������(s�^O����YcV�h`��뤣]9��k�Ժ��]�k�U_T�}ZWs��}_�Ia{+��	|	��_�p��҅��oH�ޑ{Y8^E3��Ҩ=q�p�I��G�"��3�SwJs�~�����B��	M=������W����Я73>Kr��q���AK(4���){�������Y�5f�ï�Gx�W����8;�^�U���Ml)�θ?❤5�4���l�!:����5�c&!<u;���쪛|�( y�?Z����V3Z�a5�52G �����}8�b�2��Aw!�:�O˛���4�k�
����y��@p�^�+j�v�@�F����3��1�W��#��8��j�}E��tq�cqz��A.�H��lJ�f?�u�K��h�<�B�~8�o	��~(Ne��p	�6�a-�jL=�k��i�A���./��{��E��<<�ç�� '#��Ҟ��x��A!�	�����[N��R>"	�p��^���|C��%��fo�2�^H�����j���H�fsz�W��޻�]?���ԡ�X1�����V9p_:�ܗq���I&y�^�����(���;\��`�B!�FjC�9���~'��X�����i�����u^o�Ҩ�jbK����́����-��8`o���PH޳:~׬�K\�
�J�R����(-�|:�(Q�#p���~Ȁ3�BMMh�����Y�a2w�s��qû���ܫ9|u��Inl")����0�D6ȯM��癜\�����i�?<�6��n-��r_�4b?۪<9dQ�90�0n�pL~���X���-4�9������[藬��D�����C�o�QEؙ:�\&� �m�	���y��x`�D/��|/�q��q" t�N8dUʙ�6f����`�<�f]�r�oI��ŉ�k�&y�S�M���T�_eȍPI|KL���ڱe�8��z*x�g} �C��="�[c�-;�SF71Q�Y�o3/F���ߐ/�lUw�0����i��QQ�\�г�	���0���[W5�lH�v��P�:����!c&jk���b������g��ΰ�zS,B5��/�&��" ǁC��&�d�o�$G�Nވo�u�ð�ׁ�[/�i����vNUy��: 5�)8�����{�+���Æ��J���no���Ŷ>a�ƛf�Z��a�5F��]< =�R��ǧ���7&��@��P�bB��k��"V�?�R��x��Z�����O�C�2#�a��}��B��bQ���J��҆���8M��V����R9�n/E�(��i�%1H��y'W2%� �aE}u����&䞞;���pf �beu��耖��GY��c�V����ǾNKyh�g.������=�5' �~{����O�m��@���6�7��mt���D��L��d�f����c�(~���
UG�}��H��7T �Iq����0͙�A���4JE�Q��M0������������l�56��j�7i>C�yG$׏2Zo�V<:+	V$&ݜŪ�#�$�����0g���Sn ��gֶkA}��)�v��������C��8��}�KdE��|��XBQࡣ��z�Є'�Uw�r��G��1-k}������UXs��tw����Ǆ:`���S�Ѫx�G��;?�b7���R#n���-����FD�# �� E��=��ghJO��*-R?��8���i�Kr����|�
�Y��a����o5 =]4T�RKd~�����@@Wvwxv;��2��i/`�"�S�mYX����PA'2�a�!��f \��3mL�D_y���0yo!K�H�62G�U�����҇�K�EҺ�����D���&g��H �_���g��EȢ{���r��:-�Kd7&f�9�
os��+�Ŝ��#h�t�d�kC�	 %�ێ�2n�(J`�V*]��ao߻e���!B�=�}�9�AÛ�����T� ~�3\J�Y'B�.P'qV�i윕��o� �).��(����@:=��� 5�p��}0�:��itr�FqfU��֬�n�&\Llm&�9���_� j[�9����@Yw�e3������^O�˧i7؋�`|M�<w������g�N+pe�Wb��sTޜ4�yI�W���t6�$�0"�����97��;rgO���
��TՊ�^��! D��ߟ'���'a� ����pX�O��!���������n>̧Q"�?�1گ�۵����bӍ���q����+��D���q�,��G�3�J��ihkƵ}��(6���@|�P�dn�,p�wo󣁢H�V�3���g\.	�5IU8��aW����"��)�3�@����v��V�̅h���a
U�##rت!�X?��Sh���o�<�"t?�����>� )'�|�P`䣣:�#�B��m�U,�� Z5�=�3.w���Z�w��rV���t阃�V��	�9��:@������e���Ճ��eo1��\@ƻ��x;�2���Pv������w/��ц�k�$��lw�;v���ES�ɢ����0;'-�	w����8�g��T�A,I$x���%�������ω�XMWh]j|�^R,�۽������^hsj7�ѽ��xo�9�J�]�6+;��yq��Y�Dt,-n�̆Y�L��e]�=�0��"�ާf������`?���������v�ݿ*��u�	��JܔM��ڭ�J�C��a��z��g�"#ۈ�m,���T@�X@�e㙕���6��L��TQ$z�K���&6�Tũ#&~ؤ9}��i��U�b&��B�80j��P'��~��q��Rͳ<Sq.��-p�����!徬+���+�3i����r��wn|F�O���[)-�4�8o���Y�^2���@�%���*���V�[vI:�)�~�O_g�7�=jQ���c��"����Y�{��6ZH�:D$c�3��⨒�NI���OTFc�|�Z����]Z��O?����!�|�d���p�W��`N�kʰ��w��r ��;2~�%.����@��MY��V� �=�1FH .`C�i���:�y���_�9�~w"ekL��/����]֦��J�ת5|�*�ۤ������#s�jU�kB2�%����FH��RV~���7��K�����;�� L����=IvFO�^�ܲM�j�?�bL�C-�x�X���N{� �P2o�q"�.�־.0��Ty��Ea���4i��&_K��a�S4�ϼV��vGo�|yʆ9��BI	�<��6�7l�f�4'�i�A �]���]n
�+E ����S��KJ�V"Te^A\R��{��WV��cZ�|�fw/�7�$�T`�N��o<{$��wYm�d�Ϥ!<W�Z���؍��hϷ�
�	*�)`�'ٞl}�~�:�;�FK�̢��Y�5!���#Y�@u�~9�j���#���q�����k
�&�|@i�L��3֮}D6���t$�:�'�v���M�~�YWr���S��W�s�2����Sv�a��8�c��Ə2�X����5O��сܥo_N��}��z���י��e/���8n�w�SH�Z��|��~����ˉ�^���fh��������i���.�-�=v��|� +�#!b�E�Z��W�8��n�l�ؽ_)"��~ŉ�bB��l�o�z]�rԲOL:S��'��7����7�
�(�X�,�6E��>�";�ڌ�|��7R��Z�j���Y��Q��P:op����1k�2�ϪV��j�$Ѻ��x�]%�AC��G�O���,�=#����M�"�8���H�y�w�@7!V�7���PdY#0�ni�����\S�<}����75�s��J�D��xWk_<���¹� ����A��2ZZ-����+gu��9�����*��ȃ��7q�)�����%�z����\&;��@���CU	��0@VQDQ�C_1ޕs3� -���oh�y��o��٪*�2o6��>�&��F=cs��M~ƪ�|�#���&�T�E'�=w�M��'E�ym�m�fIZ�"��}oۀ�֠z`}	�H�-ЍA�l?����g��W��=��$�N�.Y�ٱ��?�eZ�&\ɷ�j	$�rH��$�#%<�j)�Bf+���kDK��,��/i�tJ�J��U;�cd[��LH9�:m/Lrr�JS�^(i����
s��Ը�-�UD�M�*�M�E4]����]q�2�&9�y�d)���n���^ �>[Y����:(/�T�WzfD=\�:	�E~��yN7�K�enN��/_��O��ń_����=b"�g�B���B�<���I�u���m�#稓�&Er��+o��oNa����[ȸ�|�>���GhE�-�/9qv�	�M9c7����|���� Np��ڈ����:= Z�6B'z��h��[ӮT�pkr���j'V��ev%p
�`�U>��,�ZBuB�����;1chc#��x3ߛ�3��t�H$@[����ߜ���{Q��Äa�͑��q'�?��ζv�D�[���8}�T4:���M�}0#��x�h�(Mc�?�)�zAIpMȀ��'���c�-��!��q�%�G%�ʌ�O�{ ��Ē�+ى�v� _�^��'���J�A#�~�2���E�L�
�+����'���g�n� .T���(BH��Կkf`���i&WY��(�	�_L�|$�6�]cW��4������$��H)ۈ��B=��W�w�gjN+q����"�������.�J5K�[Y�,L�����X:� Ĥ�VFS̃��&�E��:�жOm���_�Nu�P����Ϝ�%E���ɏT��z�U��X�W��쁴:Ū[0Y:�c���dӻyi�̒�i�u-P'��1��1���l�&��c�̜e�U���k�j�w%������0��t�r���r�!�B���z���dr����&��M���9��Mq���5A�����_���^���OP�l��-�Da��.�<w�!/�X�0}}��Xe$��c$��_��dM���e-�*RX��ToRa?�*�\�@y�6Dp=�+ b%���� �-�<A�X�?�f��^�P�3&�8��:�DZ?8s��*���k����4��d����2z)�v�)bT���Y�B|z��`e��T�Z������^��t�R+��5�4�������~��R�	P�m��T��c�a�Ν�Lg�y�Z��|a��i��
�fkZ/�#����K#~�?,L�T��~1���.�U�����ÙA���s	�ӄIz�t�o�&}��2f�r e(8�� �?N�v��c�I�t.Џ��߰�,�$������_E ��Y��D�	hOAE|In����O0 g舐Dh<%ZpY�����D�����I��'�f�����T��e�!��s�p|��E�>;�KB7e�=��Ѽ�ۑ�3cI0�0�^�n/῏C
w�%97���
;�٢��4K�E�6�1�W�v(�;���l�ɡ#���aTA�\8QR��uj�>x"O�2M5��}�W����7}���7K�E�l�J�,=���Q�T�q|�Œvsۡ�PE��˵U�����H���2xQwDүS�d���U�K9x��͎8�6]��*�rJª�q5K�I\$H�3+si=-�x�*(�J�oJ�(�y�F0�yk�o+0�!������� �^�n�m����X�.�A�q�F�[����=\���HnEv��6�𒋮Ct�Tqi�w�D�L�����ꣂ2�n��lfkK�-�T���ξg���<[ƓF�:'ù'N��{5 S�uzLʫ��<�A�2�H-�pC
�
ꡓ��J��A�*v��� �0Җ
���l�)��1Ԩ�ī}�i�{Dd9`ia�1�
9_� L������"�8��>�5�)bϷL �q�Ѱ��4r�MNe�r޳8S,L�ʬ����S�F��Ă�^��F6J�Rɢ{�G�z9t�x�yd`���M�����O }Urv7ii��!h��<�	���1%�&���X�y�҂Y6ymWA�%��p�s�)�,��q�"���7��d�9�Mu��'e�վ��e?�ǵ��׬�� 1��k�ض�DD*�?�� zn���U5��,U�Z95��%&lf��j[%L����1������dt���0,�z*��"���p�'��p�Y��AO�TT�&�tKCa���&�V�������#Y�gq�0�ʁOs�~�%(e�86]���`;s@�����;����oU��_����N�u����/���M�����b2�֙�*�Do�	rl(:���]�0ǉ�b �/����70�~u�M�K������ZD��gµ�1�6�i�Y�*�8�Y�d�Q���~�y��q	��D)��tO����a%�z	��(�P�h��[K}�xa�� �m�6��JGY��U�����Q�02�xtE <��={���_G�x�tV�ۛ�ӳ/k�
O��4	 ;�hp���\k�CKB�4.n޹_�7{�df�i!F2��L����r�ِ��/a�ӷb����nʙs��@w�Hc�V�J6�\������N<j���o�Wm�N���cCA+�ų��#,���'�ml�h���|�|a�ν�}:˜��Xl���s��7��24j����]�2�3��dp!Nt�����
����E���4�Xĥ����s�}������{�3����3M��Ɩ��_l��E�p#�*?�[p�q�vɻ��p�[���ڄ�Co�&��!��- �M!;6L	&�1a�6���TV�'���¡�/���?\���b`���&չ7��?Ʌ�1�w���*J2�V�'��I*�'T������$��z��n�X���Vo�O-���Un�}T]��r�������,����� ����f $by�-F�Q�1%��r�kytb�8,o���\F'��w�����%Z�����ND�z����/�Y{pGz��5?ti24jf�*�@����Be�u`�G��2�5���b��N�8pR'��>A#Vx��a˱�~@v�ÁL�f�7SLƛ�D��s�>��/��Q����B3�竵����՞3�������	cf��� �N�>@����Y0�]����ɘ������r2�����0u���B	{%.��<���p%�wKiK�lǊQ�X���Ǖ��m�吆��n�S�k���>��vd����}�kj��1h~����s����{e@����!��B�d�O�����M1�� ]P)�4Ͻǔ�ˁü~���=��� ��Gv�檯�&Űɪ�n��$2��:g��6~`��_���z.�Q2@_��}v����/9B�I��6|�6��B=�r�Xɻ��4]b��"_#+�?W�5U���=�������F%�W/��ѿ�ij�X_��zQ}��nݫܬ����Gm�d>E���K|ˠ���^�W��U�K���#"�}땮�[�4UM;���	�4-�rG),���^�Ѧ!��<�E��6��YA��*9�
��Mp�3r&R�m�����t@�K.���G2K�J��yh��j�V�>�ь1Ԋ9�1']��t~y{y�gzuP�ګ���I����*zI/�xʓ�/����n%Z0Ϸ7�=�*������� }�RFO�~{}h`�ZT\W��	��k=�`�� �`e:X�%}���ߤ��ʥ+��b��Q��`�R~X/�k���b�v,=�-�ю��a�~�����\$a�?y����װ퀼b~���(��	�4ٗ�p*�9Qr%����n{X���~P��C�m���PѳԌ,��7�8�����/a�-�V`��m�4y������W�h�T^�C	��Q̋�^�C�A�>����:iG�U."_F�P,��/-�c{\�ؔ�.�����Y!�-�X]��3�7��_�U[�$I7�R>.��1;;_���!7=�M߿�-Sb�J[��c�AU���~�үp���lX�@e�'�#�?�\{ʦ�0�20�S���kb1d� �]{\��X�\���}�P{�_��&�w�7t`��en�/}�	T��+�Q���Xr��P��z!d�_\�.�����B��q��q�~N\�&��mΑ.�8���/��J��82c	z��XT7�0�Q"���y�
$](עl��������N0r���>.��w��qj��mA�_L\g0�,���5�р��o_�/�p�E0�����l�F�QU��85 �d�=��[�����oǝ���σ�����%�<���4H��b5|&$(�w���!)��gշ�̫����te���lB�3�S3����Lk�y����ªBs�j��1b�kğd�����=W�(��Rlg��qe�"x����W�A�=�l�|;����w|/��8y�+��Ȳe��::�}��J�I�Y~f�f,z��!�i[q
+��e�H�[�O�n�y��n_����w.�{B���-�v�DL:�E`n�/$��,SҧH}���kG�W]�Yy���6�3ҞW�a����0��+ ��"N�DV���R���3���c1�4��/k�	��U�2���Q�.Q���J"�Y�7��= Ј=
Q8����CE�G-�uO��sP������רmHX���̆r<e��IX]�^N���X��7h0"�1��c�e�4�<�̑�K�(C��?p#��8]�	O����b�;�3�՗.2�[��rO4��B��:��=p�p�M�l���F�}7�T邈�y�D��/��Ѿ�*�d�E��u���8�����\��+6:�b|�$�@�n���))�n	�0�v���X�U7,��&W��T�L���V��3b�.�G؟G��l�ϤA	?��թ9�J�5�UF����_�����`WQ����v�V���N��{���f�f	g+n�t*9��=���X�b{ڻ~�;������h\��S��:,*�#�	�xhтD���8�]��g���X���*���c$����:�`nf�0:��SP�}�n������'��a5
O:����8�L�Y�F�H-5���F�N��}�^ɄD�a1.(>�Ī�d��t?�ԕl�y� �Q[+ap�xQͶx��k{쏖m�`��)����G���*���n�7�� ��?. nul!������v�9�3n}�*�q�hmz�g���κ��"?�1yέ�f�Yыom'6m��8R�]kH㈎���ޥ~<=t����B{خ(\By���;�.�*Y��Ch���[�Q�n7[�G�]d�A����q�bs�U����"��a�TS�B��˞1ҡGuD�6L�;ּ�P�0�亘yM�cDa{����w��8I00C����gT[��a��ىקg2�(�L�A�J���eaxbC�m���7.��Ղ�)��sPtBQ�4c��?EFϏ�&�hw�k�g�W�ig�tEŋ�h����|�6vվx��:�Q:У�܎.4� ��U�l���ЃO(����4QN2 Qlw���u��> �jZ�7檯��T�`�	�T.�����a�j08�����Ⱥ��R��PN ��yϼ���K$鵳��}���/����N���*��ML�5�!}0��(T��3�2j��
���^lS0���̞��복��R)Jq��2,n�Cڃxl���G_���צ�������T�u���8J���!�L'U�g�X���(~�ʠ�����K"��B�C�q�Y�k἞�`e�]���^���T���7�[TbJ�(F�E�)o�X�/�F�Y�.SD�+ip��Ƣ�E@XԑD�FX��)���a)y��Ex�� ����޺�F�
�ET�_�ț�Wb8)n�h0�9��̣�s�M"H��V)�����E̻'��|�]ҭ`[z��6�sT���(M�	x���))J
)�P��L����լ�bw���0�[���
�c���g�%R�wa�� V���F�(��bU��)�əW��4�؍.��s����K4�L���&($ZD'�%�O���2���|�Q��9
8�<�m��4tż���-����Y%31-3�/:�uj�#T2�F���O�	��l��W���0=��x)M�ӄ R;#�Ȕt��U���3&쪮��vT'�T���s.�_�ww���3����&��J`�#�o�M�����j��$8�o�R��������(�LTc�+[{x�_��H��Xz�ۂL.f^G�����~_�ܥ~�m��3if���e����d��i�m7O���RĖ,��ŴvD��v���@��0M�6�N>v:d�7�����+���C�=�?��&�w��Pg�hj�@�]�0dV
��f-,v�\���~)�po�B����z�&��m
,�?rY��
��F��D�pi�Ύ��=�G+H҂��3 ���`+��/��T=\��DK	8�P���;;��萳�o�bH�n�w1�"p��z�OX�ے�"�X������$<2�V��wH[��M=�像gR�*��Ʀ�%���5B��I��k��@�B��}��ݯnZ��K?TC7��p� �d=E�A��^�G�΃\������(X�'*/kO#�6�Z�3�v|F��	83� �����H���4�}_�t�>��g��>�ޝ�V�F4\g��2��[[�&����?�Ab,��=G�L�u��DtS|�-���)$���Y���H�Yrl�^���$q1�u�G���}QYr02g
g�Z�Q+�����8�n3=F�G�}�>�Џ/x�e�M�� ���#U7A-}��pkS
ص~����B�ZaJl��W�E�*7g�m�3����yg�[Cj��`�Wg�lI�?�*�����_`�>,�?%��e�Th�������57�r`I{A��hho��:}f\������b�41��J9��!dߌU�+�Z#��.�/���s��חIE�VEЇ!�eA���g����н��Z�T �M�db&��ܑ���<�P,��ȃ*����ZC#v��=e��d3T��][����a�F`�@�/��MbP�q�^ E�+tl�4G��9�!�Iu�|�9��F75�z�WL�/8R�i���L'�i��jU(�4�3�t�$` ��P<��g���9��苩�U�v��+��up*�r�|���1���~�Uv�7:��V;f&\�y�3���Z�m��H��\B[S��}}+�m����x�;�X��M�1�k����!�������_�\�˂�f��C@F��!�gԴ�D
���(K	�}o`��m�5��(�%�us0�rpGý\q
���yq�&~L!nr����=v������,t_O�,�Q2�I�ϲN�Z�ؽ�8f�qw�4Ɇ�W?q~��#��tLu	�2��
	DN!���%"j'�x.��i��7�nkJ�!a��B�iW|�e�q�Õ�~��0ӏ�L�_�~l��hp�e* "�dȜ(��KHq�Vٳ0%�̲}E�?�sgSG̒�j��