��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��<��T�@d�Gu�!�h�����j~���C��P�Rc���FfxXs�� PC��԰�O����p32iXA�t�"�Q��&?,P#̓�*eA�9T�x��0�8nVHAG8A��J	��c���G܂y��S7AC����&� �?�,�	�B�Ũ��aU�P�̧Θ꾸^�����\�(+��F�I�j�z	�Ϩ��y�g�8!�2���%Q���_�m�$�x���b3,B�6����9�@fZ{�G?֔H���R ���o�;��Hd�����������O��3�m.��]k<�B��I_"Z�L2��:*p:߶����aȈuJ�L�_&�݋�w�����j3�����:6���Ɋ=�����e������0|)
m�N�|[d�)��H���ڵE��Jq�)Tꗓ&�^`kC��O bC������h�j<��+�E�v�)��G�i�SN�p��x��Ǔ,�z1��@��t�ܕ돹S��Iເ��8�^x�)�=��V�fE�s��a�3c�e �ɢ5xE�'�fr&��W`��r�E�m�_R�W�(�|1��hR�%�O��p�ʼvkn��I���T;6�<���d�Gt����d��qkcR��H�5=�E�zD�YX�k���B��&+8�w�}��3V��Cbk�9G��3�����h���7�#���J���j���d�]�O�x�kk�J�1�A_��,�&�:�C����+S+�p�R�^4fN���U81�{^��_!�R�q�Da\��p��{��Ox�o��,ȕ����
J��wܡ�V �p~�P�l�}8���KP��שX���B֬ȼ���_�R_�?Pٷ�x��4TZU
�4E[vS���J(R�v��3��C
�u]���Æh٥��oQ����I��Lm9-��.9��C~im�R�C�_^_f��S|�nL߻�O4�B�W
�r@����mp0�&j�s"��+8���oI���H�r`�Tɗ,��LyP�fi:3eR�~?����9|@Tb�Q�u$�Y��p �
��K�8��&E�_�J$�����!Go���_$"��˭@`���Z%dZ��cd�&ֆ�6V�'z���q �~�� �����:��x#�,qO�J���̱7५�����-�)M�CBk������-w�)z3�!n?i���c��̴��K�QJ�H��;\�;?Y�䣣��L矋�;t5^E�X���Fw��%Օ���H���v.gK�mv�
���?\:Q�����&M]�#����j�\EB'�B�����E@��a�\c��¶ �(@~���6b�P�D<����Msf���#�b�U��r5�z��Q�����7�*@4k}���3�Y[UP��nD0c˵���Iw�Ȓe\�r�a�mߜ����R��ݤ�K���	�=��x�e5��q��H�ƾ��м����ɵ��a4;�H�-��wnj�9gM�E4o��zU��i R�k�d �����O�Ȅ�s(��jϓ�i�w��ϕ�d_�.�������|�Wg�{�;����r�y�|��ff��!��7��*�l��8-�j��,v�}�~v�[�k��FW���g�AgTs/
�1�
�	�ˆw�^*ar�݆�Rkdj�����G���uI�˛k�a-.��ZI�@�]ڹ��Τ�g�wzo��顚���k<��?2w��}_~���๴�^�I(�`�a~��:�_k�E>F.��e��g�k�4 ��cCjMT�A�tv,�"����(���8
��" �^�Yv�K$�į���\e�6�����ᩣd�0E޶ {�+�j�����ķ��K4��&U��J�0�5[�65Y�Vqf�+K/u�G��yP�)~$��)t���8p�PF��m�t�R���p\ ��ֺ�eyˌ#���s�j{��g�E��M�ĉ��||�4���=wX_����@d�z�W.��֡0щӭ��w��G�g�]�Q]���*�z���n� �ۨWWcL����{�U���!�{��'6�y�l�[��:�F������0(���` �
��Aa?A��'�.�Z��/G4�����BC��-yD,�I�$���pE&C��ǓL�"�JߛҖ�����y�h�����ҷ�ϫ�PF�F��8(�8I�_y~1��?,����n����1et�yԡ�Zꍶ��w[�p��[��ip�0����f��K~�w����1��L*�c6f5'a��dT��	�M�Cs+H~�0z	K��ڮe K��q��Ϟ�4��k��6�s�!K?�f��C�26N��\�S�ʣ� ���t�(�b-g���=�_m��g��z���VU�g��[�����^�rNZ�՝���pc��6���K�y�Z1(��@���W��}�LnE�I��譎��l(�ﳛ�˶�����s�$|C�\�n��O��B�}�祐.�l�݋�˷�k$���5�r��3�f����Pߟ[����2�@�=坂r���TJn�IM։�@ӵS��5;&��D�3G�:�6��]c�<x��ꖓ���������vdlv�`�	m"y^��ax>p�O?�5 .h������?'�c�T��>�UV�κ���?��[�&bj�'zb����(WFӗm4�0�&�iD�l��)1nG�ªȕ�X\;��@�ٿ<ۥ����>�r�'��(X
��P�5r ����F󕝬�Q��q��EZ���\��%��]}�f�͛s�__�3z��f}�XB%�wCiQ�� c��R�b�e,�ܣ�Ձ��^�p��&�uh�)`CVg)�4�[D���C��W���ú\԰�\��\��������W�{o�?��6�1폫�z4����^S�F	p�c��=�V����*�|N,	`f����t�=xSL1�$�b�a<)��i��g������ĭ��$��-C1�&����Z�q�TʩE�!~��X�Of��Z����Y�L�SAQQ�D�=�t<&�G����&c���x �/7�s+B��@�h{���1!{<�2r�D��EP�b���5��Cv�^ݣyW�D��27o)3~톜�!�L5.����RI��!�D������G�b��ͱ����7�d��9w?�_���j�!��nx͜�w��`;[Vn��
\�Ȇ���`_n��:�wq��=i��?"�(q��фj�0X-?�X�F��
�ۋF���Π����
2K��A|6��)Cy<�Pu��Іy-/�,��t�h�O]�$��K�,oʈ�$���ܷ9��AbC[�p�����^���X~KbK�
N�N��C�-f>�#�X~�y��}��As��V���2��Y��g��ˈ�3P����B�m)�ǝw��j>̂B�}���F<,��0��9��_{�GqJ��=�h̚$�9R��&�e/>k@0%+��ʹ.yb]�����[�^v$��E�㖪��U[��^�x�j�����> ʅ�|�ī��ɭ�n�a�8��KF�P���a
V7^ ݅=�[�����:�����$f�T�~��L2=�'-V1�c��%��f�ޮ�ޛ��KF���{�����R����� ?�,�X�RƜ�ú�č�e�(���4w��=�j(e5^��ݜ�#EIK�1��z�q�:H�u��L�����c�[�;��!�,% ����ur�tW�\v+V�*���c�]��� Mg��0�<�������N�{چ#�t �Ȍ����9�L;���U[Z��XgEE���U���:g����O�D��U�O���0=@t"O�s�Q��P�"��g�f˄�r�����C�eZ3�\��z��d�X�w �3��L?s���{��13�9��˛!��	�˒�jq�3B����}�mu+y�
vj��&�A1��?��O3��>9���T7�Ä�� ���P�q���a�R��d�G�@�1M��a��w��}���id�/�x_����rb�x���G�$X���� ���H��f ��^Fse�\wE�,sZm2�4�m�\�Y�;���)!�4��6���Kf����z��%uN�}�]*�W����y�(�$q1�Q��l7� �&
��M�d���Ԓ���q$�ˎ���\J��8��|޲�q8��H&Z��HNv��\[�����o`YJ�U$�S�@���z���E4!i��(�U<��͛�iO��ي� �O�0Y.k�7�EjUX?sBɡ�wl��Uɩ	��&�'+=�J�����U�J�8�	ǧ��N���J>�ܪ�n&e ��Mŗs�/�_���):�2�X'�e�Ͻ�|4�(t�≉5o2M{��L�U ������e���K!Kq��١6"DoOj���U:%�:�ڢyN�.����U���#|;v���E�J2��(��5��*>�4ND@���>tл#��`8kr�F��/Z������RIcK2
 �21�[6bʌ%̔��`jE�3�W1S�ڻ�@{2�Ċ}�w5�6��D��~7����@ֈݺo�����N�zUlc�+�m�"����XK$$��<�]RV9�3����>��?�� gF:��>'�Q�&^�_�N�=���]J�b=��a7�!q���&	v���ێP�v3�:�$1���CH8��M0&����������5�*	�RiʹZ��[e�67;Z��#�ߢ�d��βBo��8��V���Q"B�X���P�"4��t��q!��"�:�P��G��	��2�(���;�^�~�����5,��R��ʋ(�Un�	l8�\4��@�_'騦~<_��f�7K��peJ>WA�u�U��񉽹3��B<�y��gO
�jڼV��T����Rϵ܄~w�%��hg@32��W���v��}4��7�e�)v�`,f�a/�x����`ͽ� �3�z�_-	�Z(ϋ�r���Ui��;X1Ym�8@�v� �[P������_t�lq�7P��L3������r%������e�K�e���nx� =�(&�;�N��/sxc�#����r�����0����|�Y�9!����ɏ�Fk�2� ��.Kpd:��\�K��吵�tPFکZS����^H�nc�6s,�MT�r�=7����0���CǸ"�I*1��i�K��Nؿf���.:1��*���r��&�"�
ޅ�U|!��s��,���h;�t�Z1ީ��I���@HZ�� 5_R_)]�T5�F4�/$$(��ћ�6eT2�q;� Ymk����dT�VXh�-��:g�L��UE��\Y6 ��L[��L��pP.5�����;����!�["�2T�|]�m^A��h��hS�\�����D@�����v4*�=�ف�Fu�)���.d��+p������-fڈĠ,"�ѽZk̞0��+�mg�-�à��It�Q�XeL�
��Gg1Tk�RFhz�y$�!�y9V��xR�G�TA\�+��U��t�,��}�����ә�&�ayr�R�%�J���~��ܽ/�@iZ�8�kZ��=X�.
��������wj���CKDe�����0E�P�k�3.ç�h�
��cC_R^v�c��c�-c���Eٰ���}\=	��:�܎Д�=Hx� ����(1�&=���{E`N�\Wr���K����@�^�,*��v^���Q��(�A�3l��*G#��$��]	'?m2��rb�b��Ĵ�?.$x�R���a�5�4
��DE�k��M�����]�&�H
̾ː��Uh�0��~Nxd��Hsg��@/�xE�+���N'���o����z���v�!��$U�M")f,`I&��#�yBi�ȅ�*0!��T@�B���^b�����+!�l^��A������#<�ܜ~�h��V9��-���0p�ڒ���8�]�<��5��f����1GgMRJ�t���F�ER��r(�)¶K�GRa��TCR�q?���)z�$�BU��g�	�X�䝟վ�:6ޝBL����4��r@Rg|{��RƯ�6P1G"��-��^W�`NE�-ʷ}��4��o(��2�"3�b��R1�ܒ�x�����z�K�/�}��pr�^䑙��:E���0L��ؐ�vk�L���*�֝��ձ�_��:���#���p�O�����%��;]�=�����Y�R's]Vj�Y�
-��#�5z>�3hDd9�۲�On�Ioإ�6��R�O1S0[�K}�V�c^���Rzj�$���|N��z:c�Zϫ��H�KE�s�
�6�K3�da�`2�g����I��t�M�.)�)b�|������'���������'�1� �Wi62��\�;�~�,y>��'��i�"���۬y`X�NC�ȞGAL�"=��l�n6v<��ߓ��u�cqt�`w2��V�N�E�ŠA-�Ԕ= k6�
2�`d�E�9�9��0����5$4����6�9�HHa$�	T8���Ӫs�ZM�����\E������*���9Ut���U���N�j۬����췓�t�C�5�ps�ܳBz�# /����Y(����4�F�UpE��_3���>�� ��f>?�>�	��M�}�5�H��e�bT�ݸH3�/���X�Kф���^�;�0��A��t���b����z?��Z��KrAkE��螮[�W�8睯.s��ǞGY����P���� ���͑s���?�F�����.܃9!����6��X��	�u&��rP��2������_1�+M'WEѪ���Gj�߉�U{��ӊq0	��a5����6��w��~6�G���w�V�:� �Z�Y����1H*]��7��L&%�N��g� ��T&���JV�!�����l�����2joP��~:*ɉs�0�Q0�s���8���kf�I~�|c���{��'�b{葫}�Cל��ȠLA���2��'���2��b*ǩ0�$��a��P�\�
Д�V�X�f����@������)�3$٪����b9��#��ʋ�|���w�q��샲�����.�)��F@��g74���)���t����3�i��1��L'7!���Y��]Z�qL~��6q�t�+��O��^��0��(�!])�px.7V�0��E��AdZ�����R~�L��Yn�c���R2A$lH�_�Xs`��f�Z���꨿��&�n����0��n����nO�[�^�{gQW���ݰ���Ar�/��+��W]��4�������I��UOIjk��Ԁ�`����%����^Xc����j����p�R-�7腹�'�1*�p5C��(����p|p;�̬�CK����R�+����)D~@'��
�G��+�2P��[<>
�y�f�E����n��4��==�Q�����p�~r}���c�U����}���y&w`~uﵐ�C���>V�`~8�1f���J�㹎�"���)c*�\����SZ�B��ݐ�Q��?4i)8��Z }<'ěάQ�c��y9PQ8�d��4�1�������|���n�n���%ћ���>,�7'[w��Ӂ]8�ۋ�n��t��$=��9���Xzzz-�C�I��4�BE3ЄӖ/�	�"�(�{��i�ߠ���·�"�
.���?ӥ���?m'K���� _1uN\���[�Ǖ0�KY��q" �ύE��i#.U��@IƝ0O����� \M6j��:�JM2z��q���Pf�2��;���Ș�"Z��(dk�*O	�3���OTL��՞��'K@I��=���Mz�ڶM���C��>B��&lx;Z�9�J���<ʐf��e�ފx>�Y	���[�G�/=�:J
hzF�4UjGǹ��^��!�=>r:i~���`�l`��ś0e?q�gz�� ���Hsg��V�3�Bt	RE��+��[�]��}�a��=��4�q{���	^�OD��un�j?�!B���&�!i����_�k�.�<�zF��WH�i�����F�������7u):��p�wy�7��j�>p��	8P[�$���}|�z��8P^K,D2&5��Zf'�l1:����#An�:'aZ��a���Ke�
0s�KkK�.4=�%����W�D�ߞ�jge`tCƳ 4(Z�cg��a��ߓ��y��RQ�:��v���\U�9�.�g�����ô�5�����J8��r�x9V~8�;,j����xu�@Np9�Ϝ��3Pi�0�o�2�Æg��3Y�C�ןЙ�t3m��k����D�1s_���}�K�Kf6��8���j*��V���5w������V$%��<,�'�UX	�!�ƨ�?����;�!�)��ɲAd8B*��ZD���0#�D*�����01�Lބpw�tz�����ĥ����fj,�ܜ�&H� X���[��}~G#C�+j�]l�
@kh��zC3a�U]e��sF�����ۮW�*u\X`^�t067�X�-�OB��R�1�a>����u�r��!�J��ߛ�`�:sC&�/���լ6�%?������E��L@ cK5p����z^F���#��T��_
��)�4:�ü!	Í\���<�su�!b�F��C����L�6F6�{�K�@?���G�����z�K�gN�3Ӥ�ڑ����j�G_7�Zײ����ۛ8��ϔ����kIW ��
��gV�>NV��@�H��/�eM$�8�	�-ccm{y���Y�D���T>��I��CP����h�f�*$�.�i��lH�mh����ig6��)I�ڊ~m����O����u�gYF�^��32�\�\�G��0��h��%˪T,��A�	��	�؝KU�H,���tr�*�����B�n�e��h�&~�墥���埈8��~ g���\$*�^3�sZ5r��w��&BH��H˟��*��]�C ,\�"F7��(�h���'�R?\��J�m�1���,`���BACe� �(Mar���w�v��G�Qt�_��Q-��qb��'��c̦0��9 �y��۟w��o&\(�cW]�샓�c�_�	jo+�~�q��^ګ�Su4�k� �S�����STRR�
�	�@���R���qƻrtE��`J�/��48�꟱�?���ӠRo����Fth����S��s�fH9;�CG�W!	i)��u	 �r��P�3��GL���,�r'^��l5s���|R�{�F�=�Ws|�ڞ3*����>���_�+v����$-��|E��v�`� �U�v��?n\7V-��O�	��_c�O���ô�t��)�#��aM��&����O.��G#;r����Vy�8SC�D�1�a�(C�U�f���ې�a�޽a�_�~R�O3�
���� \��y��^��n�Dcޛv�l��w�GI�{�Q�T�$;�[���b���oi��S��"��"k�D��cO�\��=#c��%�@2Iaf��d{j�$y�����QX�~Z3e��䭗|��V�gt��'�������q����nL���F��h�������
a@{�]�5�O���D�=&��&yk�g�,c��{��ƥ��R��T��#M��غ�"M��W�ި%��Yzg��-�q�! <���G#6��=܏��%�O���*��Z9ꍈ����W��h���V2,���ݞ,� ��2Pu��?b��$ȫ$�?$���ķ�^�����w�ۥ<%��{��Jv��t$WX�`���_��:�c�r��4i$�6J�Tj7�ܼ���O�tµ�O�%y Rh��\d�3BqE��>�o앓eĥg�k}$T�⨅�@�qG�]v����Έ�O��]`�jhKx�y�T1p�]���{�2ہ��KZ�￵���zf��z�!�>5o�A����\g�1Z
�A��
��w�����R1_��h5*�/���׉į0h�1 �`�k�y���'��HKd�2Rt�<���Ҵ+�m��X̠CNKQ�7��ѳ��3�/��cm;d����3EB�j �9����c��RK־���m�lb]����&�^([�D* ҹ�a=D4��d�	I�c�稔��^��fc�rג��n�����h��b"�9���#k8C/y`�^\X���Y��KC�̎�l����YM�M�-���n�Vq�C��* �ҿ񩅇W���]1M��P(p��Ř��G�؋7I��o�3T*������^h��U�>u���V���K�m�����D9�w|�b��[�x�����s���N��(,�M��������K_4��@t&rR����8v���Ql���Z��EQ���]���KN�:Ԕs��6��]���G׭�P]A|_�t.�B`amL�:�I���3��^)��n��ܡ�dZX��+��I��o[e��A:�9؟�t�)Jz�������h�P���`��0�ӧ�^���/�Ļ�_�
0ۄ��L̡O�@�1�Ļ��Z����<�'�2 A���Ԙ��F����M���eC��-b0��I��Z��9R<� ��My߭Uw�ɸ j0|��+Ɯ*���VO7�6+ ��RF�*��V�*pC0zGX9�!o/{:�nj=�W)�C�j��r�z�,z1�=R͑�n���kk�&�k�����jL|h��L����#�w��ʧI=���I�!1U�*��Bj);O��I.�[I�/fK�4[�xM<��l��Y瑩A�n���H�x�Nț��(�Ӑ��� �6k���g��}|�����U�Q�K�q�	��[zek2[l��"u�J�+{�W��,r����kþ&~D[�����)��|P�q�������Q+O��10���̛&u����-ޟ�+R2�r�C��2MU�9Z�s1�� ^~Sˁ��OA3��+�K�b�A��R�`�-<9,����^~9��f�4�v���7p���4���Eϳ�"n&��T����[�vTv�r�����jb�U]����e���'s��gZo�Tɴ�)���N߻���vM�!/A�l���$h�M�M׊k��~~��A���w�0,Ӧ�E��d'w^��q_�'V���+�����:�h-*��
��9,�먢��]I�A�+�0�\s��K��+-�¢ɷ���`�Y<O�׃��f���fʴ���Z�A��7E��E(��#ӵ�n���A�N�.!��)�|��M������/lb+Uy�}T��dN���������x#�g�њ<.I��F�	�iĭ|-E��i�H��#$ձ�n�
TW;�iB	i�rG�\�n��8��~���;E�p�,꡾����+\֪�s�.i � �X!�{���y7�a�?�
�+ı�_�0V��Ś)U=���3y����y�|�v�@��%4 �&�j��rT>��Pp:y:�O0��QN ��:7|���;��(TKތ�:-���V��>�!��fV�D�ZD��{�-x��7�``2��2#�6�bN�}o��
6�)|�ˈ���\BǴ�SN��2����{�
ނ�ܔQ1@�&�2��Q3ܧ)0 ��*]z3s�O[�M�f�(29����x���K�*"+� �~;?RԆJ�f΄]Ϣ`����B��{Pr����.�{E������Db9��	N8ف"W�s�ݖ�E1�ϐ{y�+�P7��Gy���>$��ս��{\b����xįJV�[4=Pq��<�ݴ�D0�gg��#.���Chg�,E�!����UIN�ª�O�ş�i�aM��C���F��c�d���lL� 7ق>R��"Vb�-��#X'��i �۹2�nl�>{>+U���t���J�f6R�Pm�]�Nǝ����t�R8�-�x�^u����,?��F�ċ���M�}�n1侨�B�ͣE�_�i+JBSc(�`5��]�e�{�Vq�>GiG����i���s��S`�]Ť�M��,��JUDʉ���(v��@0]><+�Z&/�^���P懊���g�$����<𮠆|G�Ņ���<hJjRX� �I� D�v� l�,��S�ߞ=���EE����i~�TD넲��Q`��%�1�c�j���{�쮵0�i� ����x}q�O0_���}�Rj2���{Y.�W�F���=IVȦ���+ߊ͓G.!y}��p�� �Bp癄��6����
��Ǘu�e�@ ��a������s�"�:M�V_[�e��vP�GSH.����B�c�K�7���̧��
����t�R�cˡ�@�Z_cl+ǀp�Q4�) ׾Ͽ���dm�'��X����9�e�WR�Z�G�I%�$2|�CN����'l3�I��G	�4Zr�t�|Խ���ڛ�nE�h�����oخ�z;?xY��Ä��+\�
��	S�5�.U75��!��X��cG�㹍J\�Ӌ�����xq�k7�̟�^w[��CG=�-��9^��0�^bvsj?�����.�2���¢�
k��rN�b�g�0�8=A"�y_�5��U���Ş��n�8��oݽ¿�0xy@�3x��ŷ��M�%%$��&P�x�7Į��?W�1#�p{� 5�� o�zc�aA�Go8�a9��S�J1ݩ�:��ƫ��I5��k&T.$}�= ����h-����p�#e(��9��jV!�B��Fd�lN�lO|�G���J�U��=��r��7��*���|��S#���7.�7\	����1f�/��B��~p�_����oB:���[M�Y�Q�+`����[��d�iC�FZ���I�4 4���b���c�q����M�f̣Īr$"q�`����9��^�<�(�@�Ue�Z�?��Y�bu����,�Ο�#���EG��X����@}�G����s����~����)Z:�z����ޠ��YZՌp����4|�DX�u�
��=����p�s�̙\�1�Q]^��kzS�/
CK��(��i�q"�k�E��)�W�6�`.'�.��0��Bv�������Stؘ]�������O��F�臲��P��<���b-�� )���S
~���,��-�<d�8�=���<��T5�z��=�XJ]0�3~/���/}U��8(�9J�g��l�j���7Ső��Z-JPO�=PdvX�k�O%8�ہ�;�j��a�&��V��K���o�~��݁�t��֤B=K�����:RRX���X��% �W�]��Gk^�(*5Y5b�<MI�߀֫>Ad�H�nh&�1�<=m�����b(�EUz���ҟ����L��& -�<̹b��W��N�^D�k ��ķ���9��K��t���jlw	¶o�O~��v�o���N�s���!�����/It�L�x�^���T3*���[�h�>��U3��fyv�Fo�vc(������iNK�x�]ؘ��x�FP�`�\|X �$�a�Yk���T:K�Z�d�<�{�)1N|��U��\��J	��G4�vbzb�쓡���:q�L��-��/rMC�X��;�A�w5c3|���~�L�h/(�7�y#	�v�l��lB]��'�ϵY,�!�[0�7��������7���*1���[I�P��=t�G%�E9g���t
�`e%"���p� �����/����~L���釶��+:�1������;�Yy>c��~͑�qZl!Zwڮ�v�A5k�?�~�+��$"�C�l�W��rn`՚fP������[G�Q�����$rĒ���n��wM\*kD�����{��A���� ��g܊t���bg�P*��)�Dn�:�p�떪�bƱQ���Թ���u������QjT�]�E�/���mC÷�w~D�m�T��О��|:��g�bPJ�ٿq>���������,��Y����i�^�4�-���l��d�n��")��������ݛ9z�9��@��6��~��ù[ e|^ c�'Tm ��ܴ�t��C�z�\u�7���-�	XlY�%�1����T�y7�3�����XK|��YQq����>9��D ��O`�}ZL�B4 ��Y�l��wh��}.��"�тjk{��[��Їo�~o/6c��X�Q�FlxeZϬ��S�(럩^���.Ȓq�Cv5�z�ƨ5��)���au��o������o���V�W�'	O%H���B�,��V5DB"�?�i���ڣ��zUٱ�*�A�R�C�w1�R>nj����f䀗�o*X�6W��c���m��&V���Db"u�\qKX��TO��8V�t$F?H(�=H���f���c�d8����zꦜS'׷¯�t�g(���^�h�e�/��ew�7���`�w@������U�k��B��L�	Z����C>�	�T�e{|���/��t8��:ܲR�Д�5i�T��јF0�`��!���.�Q]-m~:��'ѭC�n{�K򈝑W�1�����9b�W�D	��kE�w���������kS�n���~�k�=#]�X��Pʾ�5з��nW�,����t�x
[��d�^�I4SWN
����������ޮE�f(/�kn��(��ɼ�L2�<+��OX��G��D��G�X�Ac�k�	J���CO��	��WJ�!��ɒ�s��n�yu���e�籟�T��n����(�S�aw�H#��)���H>zv�/�r�˨O���
�
�e��L1h�ЍbLѧ���!�{���t׼0�Dt��h*H|	c]4�DV]Ȍe��G/����ҡ��:�9]�F �egs�t�S��+kg��Z�v���C���h��`�&��x�%i6r|�A�ƾ��ӭ:�?�N���va�_T���;@�J6,��ߑ�@^]�۶'��m����aV ;��m]{�#�K�@I�`�����#�漢h3�o�&��ny�)T5��S��;��U�w
�T����,ET�W��m�n<2��!��lM�����߭�����].��8���vGƲL-9ft���W�����Z�-\#�MWfC�+LU&G{ ��M�FI�F#T*�#� �o� X��i',b��G��{�N"SP����F;0c%W���tK�}�x@걔|1�Bu��I�OS!���K����3~�5��b����uJ6�����[3�v g4�Ies�E��gH~a�����@�sYl& "ݔ�r}4��؉��~���P <�ݕ�lI�X�;�����z�#�DD�k^}/@��%�kZH�(d'q��5s���T���at�At��|�I�'�2������QR؏�X�r���NO����{��z0U_p�8%N����ӊ���Y� D`�hB�"n+Zx��Tj�]��!��[�E�_�0�BL&��^[��Bb���w1���&/vZݥ�Z+�k�Ewl׽~�s�gwD��M�W��=M��]&�{�g��cA80Z�����J(�%�!5H$<@��,��f��KG{������/D��@嚋O2�C��������o�֊+l���T��@8Hy#�@Ǖ��#��`ШD�׮�d���¥������b�m��01�������k�k��C�T{B$����<�Y��"�Z�ǿRxw�"���gjzp�:sC���7%S>�C��nIl����m �A<�/��A� C�	&�Y쵋��c��2ժ;ӌ�pc���5I$1y���������!�Cppc��ޡUtl>�7W�4���w�]W�q���֢�d{1f�	K�l�ž�{wg>���I�m��
?�[��>�l:vU��Uha2�濕o��N���IV�)��h���0�N8�����L���Rq"�%��I9 �0������lT'�����I�V �"�����u�lB4
��Z`���R����t��<������NϺ]�>�S4d�v\�����h:��G	��P�t���	D}�c�%�!툊�'�+N��A�S����vp�ZCHp{��e�?�OZ�qc����dR� ��
�����#Ä�$�;D(�Z�[��u�BÅ�qTz-z��19��
��lyFz��n%)�z�R1�4ù��J�Za�:�U��=�\>D�>�=X��%�.'3��d��^���@���9��7i���Cb�vK!�~P�.s:�ؠՀ��=rQ��p�R�l1WpK<�&�?�>��a����u�\M����.5<��I��c��8,=��}.?$�T~d�?���!�~��?+�H��p��iҁ��j>��G�M��c�{�7��hol 3"{۶樅�Ҹ
=@��&�Q�L%��&-�盗����n�Z�� çj�(tO��t����D����b�`��E����.J�s&�8�*�	|I%'�>-&V�����u �����`n����lCs��j.�S���ʋU�u7�C�DC�s��Ak��I���=U�0\5�b��[���?2����[o�*/��IKT!�.��ca<�b�V����5�+��� �z/v5Lz6"�+���Y��.�e<��\W��'�-��e����إ��	���{6�o�C&�oI����=Ʌ���r�� ͫd�cK�6j�xd1<,	��⚉D�a�m�a��:F +�d�I Ry���dg�@z@DF�n9L�1�2?�OJ��h�$Td��̞B���U���Y��Xj^�F��"��X������%ƺ�i!J���H�ڻ]��ꀐ{�=U�2H���8�]��O�K��\!�΁��ѯ^	����+ӽ���]Hd�o�e
d�@�+��ps�[������ߙ��-�� ּ�(�;"��3����ɹ{ST�����b�*8HrX'P�P໽z�_������vr)�z��̓�}���eK`�hq���P}DbmT*#㰋{n����-��=�m��&37��t�ȴd�J���G+T���C�_Y*��
F��l]`$�S��I^Z-�Q�
��2�QDW�^׵~����@2K�g1(~�Z�m2�/�6����X�����s"��Mw��	 �%���*�87�s��2G��",�~��|j�c�}�Q��w�w9X�s�[����z��\:�_���h�me	�h(��W���Z�@����*�ʭ��/%���ȃ�(X�.b1ݜ����:[��Fj��B��Q:v��A6?"HqjN4>����P}���@tK�.��D�J��Z��Y
�1[���M�ߠ����?����)D�R_Tǃ�[܁��x�'t'5l\�C�B�e3���y����+?���o��w�+E�����64R��lӸ������Hk��_�U(�d�I�w��g9c&��j0ُ������� z,{%(o�%'�q�M�m��0ŀ�L�P�d��9?����*���3=t��л;�����y��Ĺ�(^�;����8��_�n�,�7w�Rq/�ol��8mu���� y�,��h��
&��{qƽ����UTQ�Ko� b�ݫ�(Ju֣0�@���ӚD��{�e|l�;J�Ў��fʌ�,��z���]&*�W3۶Sdy���ys���t�������Aa�xL�6�8���<�9��6�*����	RZii�-�B�J7vY����x9r�!���ń:�A+��o|� AS���pLGM���
$�Ui���ϒjKatU:�� J������k�$�����`߇4�B�v�.�5�C
[g����`da=�x`go7�(U��!���*E���˺���Pu���O��bgE���e+�=�%�Oj:yI"}���_oH��&1#�y.�;Z���a��
=���/���Cܟ<îw�[Y���|�h�.�,��e�"���D���<�9����&J�ᶫ�t`����t���V!�e��֔P�q ͼ�׭��wN*�sΛ
ɘl��;�ntL��>�t���^�s�ȅn^�viJc}tzdz�OW&�2��Vd��{Rx��R_6��R�=��}.Ob�3��|���zp՝��ƨU���zh�*!u-*�Q���R������CAu@��U:�\d�O=�[б`���V��m^�P�F��*>B�e����_��3`M��A�J�<�r��0���~)��]m	\͝�P#n{ѫ�}�HDh} ,tɱ���[U�ܸ������~�!dO&�ʈ��-�m�_��(�Ul�G�U�6���\�R!E\S<PV��UD$x�fNЇ'�}�1��irޡodk�iBC����kh���ǥ2|(.�L�!=Z�^�cf��U U�Y�;V��+�r��viB��% �9Q~im#�Uث��`uOD[~$�/Sم(���{���:��p����/���^T��U;��d���5k=��XG�j�]'���е)+Έ,��mef=�oN���Sj���!C�v���H ���sN����ui�H�b�*�-���XƷ�ALMv�%��i�x��.X���,��1������#f� �b,��V[�P�5�)M�[�K�d��7P2�=����W0J�;B!��E�D���=` �����d�_9�A�z�"0�JDͯ%HX\GSG�-3N_��gj@�R������nk76��,�'�홺"��C�8-�A��i^�`ޞ�,��b� �j#1�jX�ý���~���:��>��rQ�,�I%ɯ�ujTqV\y�Ѱ	�"H����q_��E�~�i��Z�m�z�A���%�_��-Z. �0���&�S�N�1��9�ڈ��w�Ou��u�0����wb�66�la'PZ�d���H>�Hf�U�f�I�u��p��1���d���쇾6RX\�ضYzEO:�
��5�u�M�� �t���'���=����Tf_Ⱦ��G&I��ll�
�4m��D�xZ�&h�����:�;(�m���c����T�p���h7��i4����H"<��f�&�}����}�ksC��n����~
�-��3�b8�B-�G��[Z��R����ɕ�'Ρ�W�5�T�˞
$D��'�x��7(*B��A�����^�^���:yረ�����t���'b�ܩ���*��B9�8�ѥ�an0���X���m6��PҢ��l���u{R9Qg���G��Al�w�a����I٭ɴ(T�``rdX�}�w��1�e(�Nw���h�)������85-���o�j쒤�p%�J)vvL�iЮ��Fub���5JɬT��>y��Pc�����TS���� el��2C]����f�����ܓ�Ӿ]��+:���Z�ͥ�5�pJ��\���X0�p�ԧ�@�X���<۹�e�4x�i0��b�ȥ�D��-^�`�1丷�D�7�vt�s����1��m�V�8o����xz;}��.Ln�C��š���|�3}�gkNv��YTn��;��5��!t�d�݂�}��с���Q�W�	��
�6��f�RS�u�O:�ѓ}�.^��b��xPd |�l�ȝ/hqJ 847��W��S�G�o�Q�XO��.o%���Ý���-^\�[u�4?�+�:(˕�kI�k]+ޑe��#�&�Q��C���ג���e�\�P-��P�=˪�w������N+n��T��h�Q�hw*�W� bc�T^�'!M��Z���뙎�!0��%�V��'�	�Zv���S0�O��E�R��+��ڢ�q(!ư�&�ܯţ%��,/��ݑ���A�d��=8�g{4Ȁ@�Y�¼@u���à��<������^U�n���Y�2`��yL̯w��"�ݴ5:�`���+$y�c\0Ԇ;�������8=�>�sf��\�r!^�Ha�䱠���