��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����)n �n�NP/x,�Fu��D,�C�)��j�vR�������|�]K�U;���A@A�qY@@բ���e�̍�gF<E�0�z� n��Yaex�1��p�+ [�B��;$ţ!
�_�c�>�Ή4�k-�e�M�}Y.tצ"[^`㻬Kg(5�f��#��D-s�q:�0eP�%����+���ݐ��j\�8��n�p������xo��|�v ��o���o�4,٫'.Kq��$�q��\�6R
4�q0����R�R� :P~�آ@�����Sx,[��0�$���E7ٷP�g����w��Ϗ?\x��%�2Ç�n�Z������eʔ�/�w(¦.o��z�2y�m��#��S�F:�..!U1��#U"�SF��A~S#��?;�
�~&�Ҝ*��N*D��bg�K�JsL�ql���dD���p�1�79F�ryσ��zp�+���W(`$� ���Mk�S�<6����%ү!LxGp�̓\�J7M��d��$ �)�.$JxK��\)�ZU�<!�R������#_�r-q�HJrEѢ�*�C:�&�D~�/���F�������^����S�C[;�Z�5����RŤ�Q�a��ߺ�b����+t��h�]�*Ԑ�;��C#��]�r����2���?]�g��Ϛh�D�;�<��l��W��4hJ>NeH.ř�!?=x,����p��dAdp��}�X�=���y �w�S����0C3U����&;5E�� �����>�ݢo��Vr�����m�4��q�=��Ҧ+$�HIgKp�PB�F}6��GXz���x��b��)~#�_�U#�=4����q�ȣ�&P@ ^\����(L��V�:�������e��`�R�Q*���=W1&�ݳ��C��b�k�,F3��2	]�]^�-��ʯ;fg��GG�7f�.��~i��������Fچ����I$�Y�@�Ӈs�d7h�)~.���0���t�h�:�����8m�Z�"��Oޏ_8��n�B"kk�|�TƢWv�S3y?��ߨ㳦D���2e|
���Z��"ĭt҄�X�����Z�W�Z^~wx]b�[�+i-ja�T/�"(���Ѕ�K<e㹌��N9���Q���G���e<�ˉbbN�ۀp@��1�Z��N��;��G�¹���X���,`����җ��6�N�t�IΚ��	,~GU�"8�h]������q
��KѸH~���p���.�ǟ�.RϚ��pȕ�2���A,jX\���T�b>z6x�X��p���$�J���v�)�]<I-��}�`tڏd��C�%N�E�����C�:��)Cݣ��#�[��7�7�k��΄����)�==�Z��;,n�RRy��))]�|h�A��K,H5��ԯ�e�����2��c��G��U�����`똯�՞n�.v[��BR0O��S�=�]$�G��s�il��������H���^Pi��o�Ŋg Mr�\��F���*���HE�	*�r�\��J�y�P3��U�'��n2#}_��8���/}#-B��(� .�O���X�̍L_G~���i����gHf�F�<���<Km�b���卥��@=�&6�a�,�8�c�t䫄�tN<�N'K�E?�a�^����*닸	�C��'���K��
���x��[\�TQ�69U�7݁a	��qz�0k�pbuT�4	��� �O���9C���g�!���t)�?e��<��#��u��Q&<O�S�Kn.NR���:�@ވ>+c���W��aA��������Hd>*���Bym)\#$>��M�h��M�q���^��6o�'w���a5핆F~v�X�^M�N8��r�ְ'��qݹH�1��],�����E�;����l�Jݧ
�wK�rF���)LA��]mm��O2Q��]~k*-�8ٛ�VG��(w<�m�R0=ޣ�-I�s�U��i��';�VݪK<�u���ܿz��=��l�۶br����"<��� �St?Wjd���s+�x^����@G��4S�ZV�Wl�Mjv���y��@�6����+]3c?rgàP[r���w��E��B[�8�8@^p�z�Tv^�����N���@z�Y���D����Z9ޖ�bO�>�dyy�Pުg����fg$�ݱOǧ�0�_cCD�U8���d��n�e:Df����&���dI�|��"�	E={[�Z�E9���i���@P��Kk*�-��Fd��
�@]� ��m@��;~�W���N�L�t��v@����L��Rb�� ���y�\���g�WoT`�4d�r�`�&c����t�8���`LIH�MW��`0.�D�΢wn�Ě}'����ځG�Hլ�*��۾�Iq��1�ay*E�K���ī���\�'���r�li�v�o���e���u������oK�`qk����ө�j�ƞ;7���aEv:�Z����)UV&D����~����]r��	h�
J
���)��3���Äkq"�5{0�TёSM�P��os ���=|�����C|9�zy\��6�Vv\v��O�?b#t��1��=��o��w˼�2?,tt�)��,��hI_�!�uF�6һV�;�b>KIЈ�	Z�vLޱRu�{8xa��j��o�ߕ�k�9Vb�,���Rzxܐ�l4C�'N�Z��4M$aT�J�\0P!g�x#�R+�j�R^���vᩨv
�dA�l>֫� ,�.�U�c�
k�E��P�L2��-�6!2��wx����|��["Nj2mt����,O/�߹��:O�sݷ)��Ӌ|�tAT�Jm��)MprvJyLXy�#0���[\�W����t#����6u�|���DS���D��8�G� ��~���d�`2�ܭXj��2*�8�������c��l�<0Ke��a�]ᩉ�7CE�\���u���:�cw��O��)����Qg�ou�&m���壃%=yXv ���ۣ)v`g>�!�!J۞���t�����l¬FA�s'< :�?m{�2$Αa���)tV\���O$�c
����;��!)	>w���h���t�����2,U�:�J�_H>��U����~vLX����!
�Z\I%��V�^���r/+����⦒,�	q�T�6!SB3��#�ҕ�tOT��2���I���O4H��i�#&ST��v��b;�Y�TՏ�@Ͳ{S��G,���^�iд�B���n�nk��lٞ�(������z��0�!��Fd3 r�Vy�1 ~����:�8 q�{�e��.����)�Dk��q*�����b��'��Ok����z�R����8dq��~��W���[͒���C����Y�i�x��U�|1��D�d^��B��"ܓ��[�<�lSLj��g�k�}1���,`���\$�HѮ��I�C����7�9�=5�L/ �0'��0ņ���͗�E��������s�
jY�e�f��&���Z�܃�~��t�����"�$%�8]z�៵w����g7��^
kHY�V�S(�0�0�'���2?����/?��=�^��8Mmɝ��W�k��>���m���[�BW����̡��Ys�I�ڭ�j���Y3	�N'�B���s�G�ޯ汒8�7�K��� �)��S>�Ie�Ɋs��zm�G�Dj��դ��R��A�)^C���ӻ7u��)��1<h�<��UX�,:Z9��i�:X����q�&"Z����\T׺��ucHDM��&�{gMG�ˌTv4Y������N0T������6ل�R�]�ewoW��#��A,"j����u<�(�68� E�*b�^r]na��O2\4 zu�����l�
�=V��ĩ��ѠM�!$璫bG�K���q��0,���;��Ċ&XD�7�+��ߒ�t�PDGhוJ}��h+���
�!�&@{W�K�M����|���$����Q'�S#Y4>�[a-��Hߩ�'���v��S��<	m=�C):���rP�YZ>d�U$p�7,֯�3�fg��� ��Ŵ��:+�8eM�ǎ��NP�������nɎ�-.H�.��Ƕ��A��%v	)�9R�Y�"%�Jlۣ"�;4?��&\R:y3�_o]8�z+�n�j
��P`T,#�Ck��|ݘD���a�+$��0~�s���h2?���E+�;�\٫0(��I#$�)��S,<���(�-��:�5�u�!F�J��DBs�$C��BM)��畴�m��	ؠb�	�&Eh�~�e
�������&�MY p�ɦ(��/P��8(x�GS�*������a_�&Q��!�r