��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���tڐ�!��Q�����xZ�H������
��(��B_K;bA|���.-ƍ�B)�wr�q�h1�oDu�j`�3|�?l�d�U�J��%��{�.Q~Ѻ:��E�)�֪�3��g��UvT���F���ћ�2�&�7}C{ ��e�9�W���Z0bnf߽���|g�tɣA/NE�CAP�$�6H�ڊ�>H!bd��=΢b��@�q�:�W�SAq;��ӻtu����¢"�����8J�mw���V�S�Y��X��qk�l+ݫ����t~,�����ޤ�y�2���t6IaN�i�}�K�ZN�5�I̚j��@چj��G#��=�9i�7�߯�a������z��@&����=�,[H���F�	iU����� �wN���d�I�4#�H�J������	@x�yes���g c�JP_�5�P�2�ԃ��PޡmD,�Ӷlǲ�G�>���k��e��+�"�µx��L�����-/�tj~J�ǥ�r��]�${�'j��[i�.�-]�>��r����@�ba8\P<l�1�E�^���*d�8��T(W�3Y��m�0��
>���G�}���U��Zj,g{+����q�S�dPH��U���T��\a��^��8����$�'��1��C4�z2R`�d�2����l:s,N	�w��?X���-�9��� � ������U���}�IU��.gp��Q9Ѱ�%o�B_4OQLἝ���E�gN�f�+k�����wܛ�`b��T~��f���Ul��ޠ�r)S����`��oy�`ȝ�1뫅��Kh�=�B���SA��{��b��-Zf�iv��f̰���?�ʐzq�g��sV�8�q"=�)ܪ���Fڹ�+�ShD�v~��-c{K7�rr.���]q����a��`t�lJ�������N�q�x���Rk��X��FF�P�S�W�T�u)<m����e+�9�cF>GH�.%�����-+�t����>l�ح��Mj����m�����!*¥�8� tP�~�ڸi�G��*�$C�MF��pZF#�Y�6�ফI�L4��򍡏��ϴ�0�f'���J��������L"��� �bx]i6n��+�H����9$^Io��W�_���+H���;�Ҵ��/0��1���+5�P<��P%�:.���M��RK�8a�A��N�TN%'�O˳�=n�g��:;r��H����6+_��~;o\�2��X���|HE���L���kA�N,�d��<q4mc��i �9��5���ϋ��5VHӨ,I��G~S&o��������tCc����"s݊"@�5�Ɩg�� ���
���=Jnr��ߊ�%|�A�d��i�%x��Ru��Z�ܪ����o��TL�Gv��hng�r�JYO6�d6��Q�3�U@90�3�R�q���s�5���1K��jr�#ǈ�H���G�s/,���ڠ�Ec��?���fp�\t=.��7YG�7�<9���iF��G>�(b��%���<�fн\���h������4��M��GB�"�C^���W�* �<,(��U�E?y;'��7��]�~��jJ���?�+��bEJ�x��P;[{�ׂ�����0�@�֦?Ļ;���/�X��=F�}e$����w�&�d�G��YX{`q���obLFt%��Z��*�����ѩJ,^'�~c��̷�.5���˝g�����g���q�7��!-��Ky�R9S�  ����r_W�'N��*/�+.�v�6�;>U3{��Ld���]۲�a�%�ඇc��"<>�����p,����M�\��a��^d'_����*@�/hv��I-�LF\��B�:ҧ�g�_] �[!�ˇ������cdK3",��.�g�<��brY��XUe�I��q� �݅r��|�5��ϛ~s�Qf�+W|�V�vp�H��b��{�|�ӹ�C��TrB�����^���a�ئ�oN�#��;�uJ#��.��+hj]��;!Y�յ�^`�U��2.0cõP�u������ڮ �癃�4��*�O�xyf8�&�;��砭Z����e^T��X~:n�2�7���&5cx��=�=�c�� �@B�,q�{�EH���'!�'�5�(�K���I�nx���V�X���(�-�yE��