��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY� �T�Q.�xC����L�lpuu��
+��5�����N6�
�C��{N~���R���`�ذmAS��k�himTђ�yZC�Jd8o�_�D|-�C<�tʖ)ơ���7���̟�F�We5H�F{��b�]Jc�)n�U����A�6�Pu�e¦�#�co��MlK�����!-�it[�e��u���޿c��@X�a�
�ua�N�!��/�5�*�(r"A��*�\^9e����絨տ�kY��j���*�9��A	n�pP�����z��K?e�L>��ԉH{!����dQR���IV]��[{�D"�g[�6eY'��2o�z���q�yɅ�D��p�s�
���:d�0?-<0S�������*@؈������V�eP��I�@�t�4V�k !�6ǡ�I�)U0�C�ۯO��${��q�\1Z�0?�0$=�D3L�ob����AZ���)Ȕ�g���eQǆ
n9�p�Vϳ-`!Y|%�5KI����3�5�?�3�{��c!'Z�m\jW�:�ޑZ�|�
y?B(��U�Q�8Z�8����)�1dv�(��^İ�~U�.g8M���$��q���}�Mz�^�o�^^4e��d|%�"h!1��w�p��|�+��$�G�e�Y�H�SL���>���o,�K���O�"S��D5Y�iܼ>DB�-���Z3�����h5�&�W�,r�VClxS��̙D�ۯ�[�f:��p�*Ԃ�ܧ�=���^�Jr\�	� ���R��G�Ra��k���n�ln���u�H��`]ݵu1z5�B�;�����t��!����Xn`��-����D4�vx�K�kk��B'�6l��Y��FU .K~��5�5�c��k
�/EP�}+dx�?�!�QQ���-)��h��(�("��􄊛�g��W�����9�w�8�들��3�/G�7��g�"5)Z��@hb����X_M��^Kp,:���:eYy�(��e�)"�^�����1��ϴ6+?Լ�f�8�X�0d�U��ԈH��l�q��f�>�Ƹp����!Z���G�w��80���������*�<� A�<�]�(����}I)����Iٻ�= �-uߑ�;�..���P�=�壴��lT�����6��-R�{�����-w�*_����Q�0P��M'-2� �lD�_�#j4��щb��	�1�?&L9�TwZ�N�H��G�n!*�x�|���4����ђ4C1��	]��H_�M����/^��g*1.��W�!]�RfSgGx���(���m�$��t6���0͗��5���i�Oܑ�F�����&F��h�IurLo�Y:*y�bq�H��3�aR�#���@�|��Y�> �*-H�X!�,����Mջz��m���L��	Y.�M)�!�Ԫ�]tߋF|��t���|*|����x�ڮ$����+f�ҽ�����?�� ��s�C,P�r;DF �%$|{=���JQ�J�r'6�K���Fw���3@KG\��+���iט(�s�s��:Px��q�Z�B��h�DR�,� ���(�bT�8<���9�zl�fFө,�����nt'h�ѯ�/����=z�5�K{V�qQ �ʹE�.y)�?	۽9F��ũ�)Ϳțx�h�q�^Ck��D�5+��k*�s+����ĵ�6�B,a�~��1ɾՃ%��ԄZ
8,���V�^v����GV�£�⑇�'���
X�4׻GD��Q��8	 �̷-9�C�1@��^�?%J��S�$�>��]U���y1*8F8d�J	�Ep^)<	\�ヶT�ݙ��/�"�쇖n~��P��H���Y퐐����R=	�եx��ӹ�H7D�3�c��S@)~�\0�����zub1
(����G�����uֻ2b���h =�}p����I����#�x���nހ�X��A��{�:�/jO?�B�br��O"�ɭOT�JC'���,�G���y;��f�Za�L(�^4�P#�<�	;�����&����pD4~��V^R�M�|�]�t�X�a�e|�T�~��^\���ԑ6aT�R|	h�Q�#��?�N��[F��]�d%�:�n{:�]�-�y.���2^Y��Q�yx�Z���2'��l$?u["G����ncA��hRE���'���I����A)Vmぅd�)/>s��3��TD���;V��+~%�8�:�3���ӳ�Mb��l"h8�|��w,$��A�r�<�%�bIԽ���e��v�җ�v�~/� U7@*L>N��\���mt&9�bLz�0��Ak�e�����p����	�w�)*ݳ�a�A��j)�|&s�Z���u������	ŲgP4��fꢶ;�Q��H�4IbHʎ��@�f��9VJ��۹�C �7�����I{��>�z$�CWdq�����3�R�<+��.�b��*�"���X	�o�U����͵�T��F=.�7����V�FƀӸj.J�C�#�����S��a�_��
�C�lH�*N5(YR-Z�+�#+����nØ�� D���8�F�j�K�o���)x���u�+����t�Y�u�R�&��O����j��ϓv�"I���K�K*�S3Cn}'���G�����z�\Ƹo�4�n��-ٹA0�3M�6kO�&+�ߔ���c�Vz6�?�;̘f�1��&��qv����V���
����R�^��4u��i���{�(�=)���C���#S�r�u=�pݖJ�9'۰zo��P6Ku�t���vzw	V�u�����m��"vr�㼲��	�ra�����g�fkG SC��]�]H�����QXCc`��(8��i�ډ�c�Z����/˂�q�	
�����>f��'.n��[
|(<�������e�f5���t��%y KE���V��G�a�X�8�6}�t�a�C w����\Vx)h�w@�m�D��L�3�C����f�2y��B>���`�q����@l��V��U�g���6J���0{�;'v�(/f���+]�9�+��v��'��C���jn��p
'll��A-:c�,�9��G�c9,{�҆b�"�q�l�Q(M�7�'��Q���mrT�Mj"{�7�ঊ2���a]s2���4M�=;$�p�zq�9��R��Q�LO�Y!:�w	�ˆ��q(�O'n�:t� 7�u�l~��k��j��3�Z���{ҟ��2��Ōט  ��,���P��,튾�si,VF�
�c�'4r5��8�`�qӡ-D��%��*G����|��#�	���%�F;���b�2MW.��r�����J&l�ӓ΢m�c�#=5bP��B�^�'�L�2�P�A��k�-<K��L�C@�rf�i�6��}����4��L��C��	����o���J�����-�x}�,4��3<vD;���q�U�m��9�Ŀ�Քy��Pܺ�%�	�������PzA�	�Nc���Y߻�k��������%>���i�e��u�%G����M��a��Ov�r�]��I՛�Q�n����yW�@h��[���u�����A?jZ��zpǳ��u��A=��uS��	�I�.�i��t���^Y/�]��rQnC�+�v7%�Ǔ�����' W%5�����	SG�cS9�n�����)cԎ�&s=yI]�{ek.@(�ij,#�IT��j	E��

E7�MXuS�?�8�A[W����yq?�7b�O*)'�c�U�Hxd06;�L�p���D�݁G�Ё����s_#v�%~	O̹���U?�꣤*�P����T~��}��<�=����}��[� j��x[�r9�ҤJ")�-i�^�<M�#�>���6�TEj�3�!2[u��]�Ի�m$��K:Zu���S�Vf�;AA�A�����c9�~/L�!S�~����\h�̴�o��K�A��N[�J��l_��8�����&欭��&��]t�l�1��W���؇@9d^ʢ�T�/ɛC��$F�0�Nѥ�X��Tz�̢T�Hc?����u�F}@\%�?V�s>�Ӌ��Ր����t�8��uǙ�]r�n�Ćv&��4�e<���C�,�c�>n�̍�We���"Eyp����E�!�K9��"���.����wUutL;,���ӻ�����%{N(oR��m�#��֣�=�/W�����O�B��s݃�&H�3�u1��\���k*	d�����>y���������-9��yV�<O1��랪I6�^��n!n�Ƙ����$X�Y�L��`��Ƭ�NI�s.���q�;�`m[&�7����?��0�Y����ZC"��#�rgwq�D��Be�8߫}�tV�sI�x�lW��M,���l�U8!ug� ��(\nO�n���rG���ׂ�(6��}#M��y�毤��� �F!��|yϸ�_EM�k�)黢����h���+�uX���6r��2��R�4�� d�6
��3��D�Y�@��l|i�X="E.fa��H=�j;\�=2�;b���\��x��,�����$L6ȝ�2z&�Kp%���1��X��iG4��V�S"��􌍈Ih��d��n�|�����F���u�u}���Iq�s��>����a|t Pq8��IR���!�!P�g����"5����<i2�x������(r	�.�hF��Z�b_��Û����1�rI��j{�˱�[�ja����%�#V�	sĝA,�hr$�d�.��ɛ2f�Z�A�-3E&R�
zc��#.�#��I�V��CE�d�a�$+)�jå�lqN�R�-Հ�'�%�c����s:��ys'w��4k��B7=	Q��VZ�B���oq�����|a13�X��4����	�Zx�D�$Iy�/��}s�E��W������~�2�4׸����2�9�z�VT쁆
��Ñ�� �_��w��ְk~</�/ׁK�葹�q�&'-y��u��~���餱��A�o0ޕ�pWH�@��H(�i�%�m^^΃�׭bǽR�@��]��4(Qu8����+��!z�P��fm�l��g/s�|g嶚�(�w������ ^���Fb�@�	�$Gw=t��Q�&�1�u1�q�°ٛ
w����?��$�K�b�_�����	�s}ɑ���ăƸo�8�N�NB��@��I��$�(C_>ʳ�e�=!�� =�~�>��f���S\9ڦN��-���!���D���gg��l;��|�V)Q��Q_(|�F�����M=�F<tě)�ҕp�L;�>k3�m����(�zLYu"��J�۫Y]#֢m�d�/Dh\��4���횺���K �8nL�G��Ku�Mh�_�J=n�t�pG"m�}�H&Q�^�*��Z�k����.��_.��� =�/�v'V}�_��π�g��#<��_���ݪ4�h]~�6v��P�5^7��˨�蟦X=�Tn�gT��+1�%v@��Dt��F��L��Q��£���} ��U�]�M�(�a�J�ƥd#(ޤA.���(�C����n�.Y޷�L������<���x�����GKL��)��{������Z��f��_�9�5��|3�F��Xǒ�g�*z��Ä�����[�=ۊ�`s)�l@��Uj��n��X��>��LyJ�GǄ���2u���m���+TOz���*.g5/y
�����1��"
�j�t�� ��7^��X��l5����.,��<T����;-͚g ���S�`�s�R�&�5�;0)�Թ:���v--�:*��	w혙�շ���'�gD��YZ�*eU�6����==�$�&�Y�k��m&�B���0�EyL`��(��%�V�a�j��(K2[%C����{�W�	��Q*2�q�]	����OL�+<ή�Е[���T����]�*�~���U�ZPr
 �w���}Xێ�L�ڪr�nxZ����-Ro&���"dT�
��x��#�����O�ס����&�]�)Qpo��$�;�P���f�PM��$�P�!J�Q]�Z�����7ߺ��N�8���6'W�����f	��#a�� f���