��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY�����$�z�4�QT@��+�CR�Ai𨡤I�'�*�A���t.f�~߉�5\c�R��@?�n}#8%f\�n`�W޴`s����#�Bׯ���ų����<"[�����UQL?��X�l�躳P�9���{E ����7�85�[D7����Xٟ�N1>��3xlF���b]7	W[t%��xTplA������zޚ�D7� ���V�ֲ�@���p��Y�@�]"�ɍ|��Em7�>�qy�,��PQܢ��i��P�Ȕ���f,�Oh}�B����߻�Y>z����`X�=�T�$�uh����[�ԼM��� �0�#��|�pM�`�g����U�_���i���N�X~��֑=�ݬ�`u����(~TG��@�k��X��7#Ք����V�+p�N����Z��M'���J{;��/� �
�5��F�+��"��,WX�
oP5A`�����ݓ�S���E?Y��oE#��k���v�V=�]jٵYϵ��l���;�yǻH���ʽ��v�
��p�i�gB�S�p1��/Q}�W(Fݿe��n���dirs��y�׈p���^����z��� B�q���T����� ����ŞQ�=p<;�D�P�4�8B°۲��w�۾΍<�����%`�ʜ�i�Y&:�,tP��<ae;�'�~K�=�����\*���n|ȗk|������ �׊��ږ$AJ8�=����\�ST-2���t����?�.�L�Z$���S��,�^Q�Uyg�ȱ�v*��l�$i���p�1���P�;OI���J8^��,��j�(8*> ������s���^+<����hH�MK��2���@��
"0^�3���, �#��(��B.� .B���^΅�	ب���O-�X�����"D�̽M�;�l��&�#a�PF��K9B%����* �z�}/��[�]��SEN\lG�Ø�N�Ku�W�+����t�	�?�Q<��-�&X���Qc���!d�b��p�S�xk6nn�1ׇ](��F�rٟ�{t��׾{��7�B�Ʉ��"6u���}��x�i��Bc�]�������mq4����}�-�
�^�����"F
�J���߫`��Ƈ�~���������[O�$���Aoj��x5"��[��F�"m�� ȏ�Ek����cR�E&�Ux�֏��*�o�î��x�����	�� =F�!��aj�oPԱ�ѻ[c���.~,���,��f�ZL
�r#W8S�Xz�n>���DU�Lvl:�Yj �� �ɓY�e�*�;�%3�X�73��s.��H���ɲ�2�۷�d��@bo,w8��";L,�O�����ӂHG+�*�Gϥ�	�	���#��d�I���	���.��'�bP��ukp�_�l�ж	���
͘F�E����ւ�'�)|)��7-\�q���[���� j�\kh�.��z{j�kW�z��_/���Th
�?��b�4{i�C�B ��[y�BJ�!�!����<�EJ;�_s����xSG�b ���"[��q`�N�V��5��n&\��z�K����Tj�Z�K`���w�^.8iy�/U���~E�gZQ�ȬY$%/�x�u�'8~u���VS��v{ؓ��E|P��*�#����+�����Z�oɎ�Ԭd���#MF�AJu{ ���@��W��j��*�6���&�A&��@!e���b ��#�Nx��Eź�u��Sm�dv&��!6��-�Z�P����}�fD�3�;��5�F�..��Х����[$��y^4ܶW�t�
>�3捓,��f��zN�ay���kV���n�#p煡e���	X��n#�20&
ĆJ�
�j�jҜc�?�[����,��l�|�3��<דǉ�V�տ�gX�\�������0p�F��s��
��:�<���>�K�����/L^{͹$�\�JQL�䋦�([�|�'NK����s�w�>��Ő�id�t|=���:u!��r���l���l��I^7���/kK�����,�q�s�%����5�
���Q[�R�������{����~��əYn�L�(�BQ�:�#�L����Ӯs4��0���RǄ?�(Da�,l������E���q/	g�
�;�z>���j������g��#C�ѓ��Ba�T��[��u6|:y�u�/��YۻJ+1>�Yr�?D[��Zz�V3#�l��'�斣V�+o����D�V��4�\�a���ń�l����S����"�M��z(0��3�w8�+���>�%E�t2���� �0 w������E�-+w8����}祧f����c�*3�Ɲ�&�|�g�|}d�˫��e�Н�i�X��6�K���=fU�V��!���$�Cѭ�ݔ��c�a����|�ߪA�|��XZO5�ߓ���_�A��X*���$�l�&4�>'e�����v�5릿��u��t ��D@�y�3�� J����N����U�
�}��b�g���(N���{���W��V[F�`��B`oj�M���d�c�+�<U����aQ��8P9D���Y�\rk@���<a'A9 �r���?$
���5g�GX�o]�J!��6[v�gJg�Ys����d=����)#�5�
 �\g<v�?XcyǑ0�EV�T��X�#8���d����8KӚ�sv`����-\���aMy�4_)T9?�F6�4|dX��V��-�	�<����O��Aivfͨ����a�f�96�3�᧣5뛞�j�o��� �̄���K�)�|z��2P-K�(Q�<a��!o�g��x��}Ac��#s^�PV�2����S`�G	�z��3s�w~��(��u$�;^�*Yw���S���LDn� ����_\v�V�W8sP��L�U��O�a���}B�7Īf*�'�u�U�"9
�_��d�Mr9[�� ���|�=��ck���s[6�k�yc+-���Ru�A��Ј��o�Ο�GxBa��!����		��Zi���O��]�<����= 5���7�x�^�Y��1+�2�(	|�
5��0]=��3�;��u�:̙�h�b�A`f�~Y�-yJt*r��ބ��q�\�N�x�j�ο�9Y7�VN�Z[�c<��ނ��Z�e�uњk��޼�=���d�?Q�CKf)��`�A��N�s�W�3`o�v�R$?N�X�x���QM�Ƹ5Q�`�U���x�}��E$2D�ֶ�4�]PS�}��l��.�8�{..�#�u�!�K*�L@��N\�&�6@��S�\�&T�!����f�O�$�Q$捒�2�v��	�k���.Ӏ�Hmþ������%��Y'���r_��w*��(��{�դo�Щ �E�(l��>��X	C�1,~7��C;�j*?�@o%Ӽ���Ϗ=i��yӏ�)A���?�x���u �����#<����ɣ�$�/�vj E�[DG�w��E��/Z>�&�vp�$�����nX��	�lN��
���J3m��k	�⬱���|/��ˆ�����އIP��:@�Ҧ���c���&�|�Eu1�r
���Y�V��f�~��/�BG�H�|�ty��5٩��;��eO�ˠ���CY��e�y9f�֯vM���)��[�>����77�Wo�|U��PY��dL�çFUE�a-��<=���=꒪�Vp|���p�1��,8��R��K%È9�EN���񈏝H]�����[��V��/��U��������J7��z27�p*^mH�z���X�+j,�(�4�4|bE��p�t����~��f�N ��_·�7��H�Ѫ,9��~G��-�x 	++�-�`7�U6�����4����P�w��k����o��5	YhR��(�c�T�݂�6��iyi�[�Ĕ���5Ot���F�6%y�Eǉ�Ub}:Z���-&[�&B��l�X�z��ݼ�ԩ	��K�8�
*�7�]ҵ������J���������{��Ν�$�{5������C+�x�K�/l(6 �[S�hH7�z�x���1����<Z�^��\��1�HOLIh��:`ngsl�(+���E�bW��'�L:'�$�#2u��V�OW|;�X�;�j*!0B�x_�KJMx|M0�����M�c��������#K��w��;�tS�6���26��f�Ћ7�����G7'h���5�N��"����:fd�]H��x��F9��l�e��Р2��A]C��4�p�Q6:(ܡ��g4I�%�A��--�R�� ��hrV04����� `R$����v�O�Q�?�E��gs�N�2o�J+XhR/�IȅJ����Sv��>I,�_L�y��V��n�D���&��$F;�	�K�3��z��T]�h򢷘]�J��>�u�!.��~�j`j�	��y�b+hv��j���9O��8 j������m󧺊��;cB��X�>d�X��y<q�X�Y§��l���`&a�X���MJ��e`5��>|BTJG�(�Jᙠ�V{�.f�ʁ�֖�P��3�����C��@�'r����Lr��)ӯ���N��}r�S,yĂ���nF7NQ ~���xܷ�͈l+��=��+��_>�Z�V�M�Ou_3d�Ix8Ė�7��£�9�Zd�����p�����F,���ř��T���NT��:�I/�����I�lYU����ԶL��0���7�b�AE"��>�՚j^�u�,at-@��J�^�D�g1i6�6�ə\!�x����:��(ɬ#��\���9�f��¦	�v6Ѿ��0:#΋ۤV7޽�Qޜ�.��r�EPwџC��.��tf�q$QpZ�{j3��eD�p*=9�E c�*J4�a��ޣ&��I4�O�4�?4:�]$/u2������!ã|SD�#G�|���J��&"۶ؙf-!/x;:\Bl��[A��<�;@P�Z���9^�R���� z���	�8��W�ωĐ��OG�z��2�6�H���3_��'_#�5 �DȚG�`�Ϳ��wπ�Հ����2�B�{3){�N��Z�m�ێ:mx��ձ�k�G&�\��R�q�U�	���`��Z� ԑx�ͥ�tU��Z&f�V#�"�p����'�w�>��qW&7}m8`�F���}���D�,*'�R|�&�a_�/4E�5�b����vn��8궅�_�t}���a���Fb��5p��*��'�!���e���3� �My>�n��z5�J�<�/��G{x7���qu)|��*�$qyv�/��3��"ny���c�u&Ņz�a���S��$5j�0SԴ�����e�[���LՠpݢD����{֨�9������b�ؽm�4VQ��蓐�qNy��M�`;�n�>���m�s�Jz_�nr�ن���q�,#���a#�j�-���4�p�Q���C��{������7O�ݞ���C�@��ذU\ ����#�؃����ʐ�*3�B�?�@J�|���D˶Z�Bɴ�H��qE.b,k�}�j��L&r+�|��-.iK0X��'_3��$��'��gϛ����]"�h�A�6�-�7mu�L�5�1{�)�Pd?z���]+��p�i�k�g�u��ܟ:��v�a޽�,Ae)��N`eCO��B(c��`}�X �	@�_;��v3:J��+��,�dh�n÷��c�=�`�(�J���iqѩO�Z����<X^@�\qm��T<� c6��`D�������2�Us�}�[yvq�W%�m��*ܳ�*nj �By~9Nfh�ܥ�Yhl�]�b�Qo�m�6��q�l�I���D"��+��>	�W�I�U�Zٵ,xwH�3�,�� t/M����L�Rŷ���/j񮋽��X��)]�<�#�`�-��
���W�Qn/�����ˈ���'gd�Iw-IV��%L��	�fRk��."��,�vi��q��>��&���i�R����5��((V��y�W|��`�;���=+Ma�Շ_C֡�����<�	:��j!�1�-�8Rq�oY���@���15�ƀ�ڽ�������|M��Z��	\�����XɢH���i�l:��Țe���Niqc�J��y��c:�fo�'&d"b�Ю�n�����/#�6F250#�F�L��v*Bԯk��}R8qK�`�SS��qN��� � �O��c��P��"H�)Z%$\������x��*���¬�	0�z�1|�#6�S�:~�	M��`x���JU3�,s�w�K^0ڝ�B�%cOӡ^�c�晨V**�!���؉�g�9�F4�d�|9�"2V� {� 8���e��}h���%���'�<�r�x*��x��21g��J[�u���?{�I�@yF@Y�'kKȭ��$���J�z
}]���̭�H�GF�)Τ|��'�Cqi�e���y�Y����eh9ͧ�/m&�p�&b\�Yp�Q�ysޥw�����u�vR�)%�6�@�ա��.�3���bX�⠀կ	UF��^)"%��PZ���`��� ����!8k|����/�Їmh�fk��>f�A�����7�it�O��2�Jc�*��D;��!8=>�Cæ�&A��hdeP��o��E�$��J4z�fz���v2���ВLc�tJ�
=���]��������b�V���6���LYb�y�'	�ԋ�^���	��^w�0���b��7�K���Ty��K���j���2�U�F�����#���l�N�M�^$h~g��m�)�sY�,z]�&�����}φ��Ǥ��v0QtҰMh�;�I�y����M�a���;����_���%l����%n�l�9}I��& p��u�z�񄧌����U���f�&I���?T�qב��a����#h(C�^��|*�k"u�/o�z����P��i���6���G+y��e�_��bp �T�_�Ȓ{�tz`�x�;�� �o�{S����˺|};�,lTE�$-#��th���4ѾZ��*a}�F�|�H�q��-�i�hK�ur���νXڃ�$����.�C)d��I��dT�Kv��n�L>�Y	~�Z�&|�94H�O�q��19$w���恏���ø�[��J�D�LG��<��a�w��(����>_�ݽ�O�}xk��?�o�*�wvDà��(�W�g�_�C4�lсwt�%[�u0�ޒ�Uo]H��Y��fӰ�<u�ƒ����/�ͬ��jc�Uueg,5�Υx��qC8�#�������[�&0sG�j�i�8㗎�����_�N/�`A�<�(5�� >�)|���!)+��3�d ����G}y�v�~�n�&/������^4��	��2�JzM��� ������I(ac��,r�"��Y�C�4/L���M�re��{~$9/+ ��B~K	Y��!{"�52��_�0KH?3� �+i�C;��yb���OҜ�Fbb_l��?�Ҕ����Xt�.�'桧Ⱦ�=�-��p��r����k�rN��6�@vhf��\�2Ò}:i���[���8�J�@`tb5<��A9�!�ʢ� ����6�}I�
�0~
AF��[�j�L�;�si�����z�j
�)�7xk��d4�r'�����hWR�I��J�`
���,��!Y�����?��/|����T�>���Q�ҝ8�)�aq���=	�����0�l�X��sb�J����G�Z�/b
"��i�!���c��ǭB��HP	ڧ}h�k�:=mu���\�?J@���}������kz"k�i�^�!v�6D�	m�D�J_e����������ęF �.�'��R1��\�e��5p���������HՑM�@;���evE�5s�&5H�Y�Mw��6��v�|-�F��mM�)w� �yB��W�9��Er^%ꬽ�������y8�:��\9��4rBe.��n iZy5\5:g}H�<)*�∟��M�y5���I����3���<ڬ��4qr��e�� �#�� n`��P(����%e�$������nA-�ڕ'�J��#_(�x�(Z�/��Uk���H96R+��w����!��A��2���Ěwov�JH �,Im�1AB���`��@����y hR �ƫ�>�j�F��Լ�;~���EX)�na��V��ٮ�'@�Y&L]�$�F0�C�4�f�&2E����+�O�3NT��]�fxS}.��ͦ�x��Է��'�ݻ�!W�N�`�O����3�h�n�M��Βu���i��/��9�U�'�g|>�70�_�(o�_���.�T��)^���.dz�1��}��>��&g��ı�N�UŔ�S8`���K��F_0���R��5�Y�9
��ݮk޻�޵2��wQgu5������sr̪�o�տezP��>!l�^��I�^� ������_0���#�@Ex��tDKka��8�G��j� M�L�����Gd�.�����)U,�T�q�5raC�Tn�_����z����́�"�zq�d�/�I��R{��4�0�{�? w�#d�G�4�7�'�n_�Z0��5�\�&E�D���e�l*N�!KAΰ��_��T�R�܂�a�Z�jޞp��`����_���ng���7��ؓ�n��L��4��j�X���-�g�=,U /�Þ�m���g���G�5�[q��>4mA�l�Ю��g���NE�Q�M���{]�2�����c�c�$����5�P"m�\���������������˓�<TQ?K��݌f�d�ν�jF���c&Ps
D��h�*ۜ�<=+܏~J4�'p����YԀ����.�ƁM����̇(��0uX�q'����1����p���G�1L�$;�ZMAK�U�MH#i{6��!�u ߛ��t�j�:e�.�Et�!���gz	#�j�ѕ8�E���?ԕYTԑZse��m�W�<���f�L�0wlؕ6�=3�YV�i�Z^��Dy�����qz�� �6��hT�Y