��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY�ً�r"�Q9Ծ�d2tȎYO�P��]iq�L2�>l���vu�5��N�I,~�bQi�3&����4���nPQe�����ܴ֠��ҢiH�9%+�0J�����֡�-���l��`�pIۿ��4���{,��׋�p��e��ȹA[��͠����U�@��2ꢡ4�^@'��=�Ly�刐q�懽P�	Gg�Q��_��t���D�¥SL��~ժ�Ee��fI55(5��|H��
���Mq�9�0�>�Ǿ�n{j�j�f���Rj�>	ԙ�c�/u:�EF���-��0N�4�릤-Y2`7Drn1o�~w�j" H�E&�#?4�3 ���
�\[��'�3���w����� zБ��bCglݹ����x_���?*�X��s'�"������c��n� �ىл� +�e�Tg�2����9�|�h�rjm��ރQ������}������V�
^C$kU8��\��#�c�}��7|Y��B��*��.�pZCb.��ߦ�����^Kh\�>��*�z8��v��<�\Y1���m��|R�4*��4Æ���s@�U��:���6�>)�GA=���)x��:��=S���آ��L#Γ�ά�r�{��	�rU{@8����{kL�\�d��8s6L����.d��C��!@
�F�V�:��#���J�#3
�T�G���6�u�T�^cƎ���FE^ɴ����y%C�{k�����bG�YR��}����$x��=ܹ�1[?S>���v��E���"�5�V��i�k�!(ᭇ5�_��J#jV
 �^r����aV0�T��@���ܸ:B	�@v�Uo���R�.$�mm���&�
�r#.��=b��?�diG��1�N�dΔ��/u�1��$��\����Kȸ�}z�n�N�k;u�>����w6�e���u�E p��w!���VVP��a#c�� we0^�su�|S�¨�Q,��FU�tI%��e���cB/GJI���f�nSU˫]�J�ƓR�� r&~z����f�;��Nre���v��%G<�<pH���6��<�3p�!���P��HĂM�WH�ɼ�]�`b �K�b"��Q������߈F?���
�}K�ܾ�t'Nj�}5�p>d�?S�^���Йqy^r�cž�A�frJ����ј��D=�F"M���j�3\㤐�:��6B����q��I&�0 [<�����/϶�F���hv�B�k�^�a�`ÿ�"�|���<�	�bN�Z������'��3�
��d���O5�M�_[)VAN5�%"x{��h��]�kF3��hW�������K�*�/��?�V}��é:�/�h��=��`�ђ��E�K��Zb_��OM| w�VݙH4�TF�Wk�}�;��li��E���P���K�!|�ܙ�?�6%��#�����~FN����8�����tO=0fJ������I!q��k�96��BI���C8�GQ+�+��@�׈�~�EN�X��,]��%��L�R�
Ĝ�`0���������0җ9�ð0V��9�جa��U=9���Ί`��( �A����B�g9���5s/J�b�pt�(����'�D�R5�qXT�z>�z^D~�V��#�:���RZ��ɧ�s?b�79�lS���JZ������l�JJ٘rh0���֏<�kd�Kn�I�*ia`��n������g�j�?��#���F����Ӣ�x�{��(̻~D}�r���#�U�;��|,F���E���<�+�Hɱ�
ҳ���s�S��M��� �Xh&v*��"��L՚Wv0|�cS@���Aê��ؽ��٤W�$�0n�5ҳ��~h�D�j�����'�&�נdD��2��G��eK�
�:aX?����B��.!����U	�C�G}<-/�"g�7�R=qK�Ɔ��ֳUҖ�є?�5�3m'%3�$�����fs��|��vT��F�Y�6N�ؠ��;�氠[�I�6�'�<ɵ:!���1aK�X;�ZӗL����2��%Ff���&���,�	Ŧ6_�:=F��P�^D NP_ļ����Lg�`�����U�S�UM���~@�\��l���W��Mπ��g6����K<%x���8��$���L=�����͗)G���>�a�����2jg��0.� ��U��,ߙ �l8��v(����sx��W��qb}���qD����>ّ��Oc�.��BH7�l�΂eE��}��N�����t���#����wZ#z3vB"�K��ş�����E��"M`�q��(�P=L�x�u���(Y5?.��+����:mm��M߁�mm�s8���s1�x�H�[���ǋ�=Iۍ7�;�����1H�h+����IW��`]Gr�����S��-a���YP�q-�3��ϗ k˱n�F����z�Hc0+�6H�0�9s<߲%�_�6,9i�o����<;�K���~@Cxg.����=�p�$�+-���@��D��|;�2b�5�*]-!������Ų�%�2��� qQ� �Q��XW��U��JխJn�'�W�5A�Ύm/�5�X���Xr��]�v�"�.��+�_�:O��{���Ø 񝥟bq|�������i�<��<V{�ju�r�nt�=�wmI����7PX"EW���l����$Ҹ�v�ϓB��1mǇ��M0��P�'�۶6Ϙ�I�k���"���p�$�c{�Ub- �zkFٝ҄[W5��b
&��*����!��e+�ώP�״���{I�v��xw�|��+�.%�ue��4Tw�iHHL=7S\�
�_�U�!�`ᑂ>�;l�vi�1���_Q�)C ݠ����E��SA��"����~}�����p�$�.�M�\��_�;B�AP\�E�d�B�TR�5C�t#�uHg�[�e�nk��J������,ظ&c�\�*M�9�IX&G���"^]�=�|�I4�;��]bn�N��&�qY.�_]�{�^�����G-~@۪��&��U�~��)�-N���ƻ�.�kة_�ِUoA����F�B��2�kF�� &=�����%�(B{\�)���T�8=KC!n�6	d�D�Q����A+-����m5˵$qd�s{�����#�"��̝F�
&�=�+�j�Uog\Z��C~���A��3yŞA+�������V�����IŮ���&R��#�Ӽ��Hc�/��q�%��W���V�#��W��NҾ�E��d{�J�d���B�5ϯ�F܅	T��v˻"�,��'����;�h�]�.�;���b�9�e����'h����{4�f��uKO�;�q���A���V��U�`��#�$;���(o�s3'��Yu�5n_� ��/��ʶ��Ed>�]z�[+	y����p�����u�b{r@������j�=�3;���߈�j~8vP��#�������4n*�f3
B۴f%{��2&�)[����)7Fq��W�Âx~��C�R#��Zf�R�XU-����=0��|%C4� K�DEr���^lSÀ�y���c�6bpD$�Fz�x����G�,� ְ>�Uw�+�N�/���-��,�rL[��B1�$(�o�̮���!�Ersa�㤬��)�f�oo��ֲ�X#_��kkKJA&��Xr�z�̢s�%��:��ݫ�Ux2���gy�i[I;I�����-��d��
A6!�F�<O�@����ԩ�mU�]'kD_�1��ԯ��v+�Y��aP�S]m�ܯnP�S�F����@�G C�螳��YP�Ds��y ů���)-_n���
��x��˂>@��&��Ƚ�GkF)g��p��Y�����t�wI̓$�E��p�CϾ �L���).-��@P���]����Y��X"��AV�Ɛ� T�5��;|��N���]/�^��?�f�Q]"�����>�Y�͌N��e2�ol�q��lB�>ra咊8��J�[�澉�a�.��$���v:y.�g�<X��%��&~����Z]࿼�s��m��:�� ���NoJ�RG���V�G�D�<4HS�ht���^;�������e�T�C��2X>��D��N��ġ��0Rz�n(��#�V(��(�8�@�W��������\U-9sq�+�Ft�M����C�/
�V��M�E��{�jն;�GxU���*S�����6 �v�~GP�x�SQU%1���4��Z�qA�F�"��l�:Lc������k�l}�	!T;���ќ{��X&{���q�F5�ͭK�������q~�.⃩�V<�����ު� F�'�"�N�2���vJ��G�e���W&�����h�߈o~����b�v>deȮm�ۺ�)��Ì��zk�w�Z�Z��<��Ք�z�
�M5	B(�<x��VS��G�͎
ڕ�V_$�5�~�B��q���&�RŦ|�G2�(��Q���R��4��Gb��F���!(�����}Wy�k����y�r�$\�4�|� �)�D���႙���0����e�I������i�=���V�+p�E���O�3�آ|���-'ۻ��t]�A��5�d��Y��A�rah	u'�+>��� �q9����,vF���S�6���AgΠ�rYU9m��K�bo+��0��0�Gk׻Yt豏x���#��~���_��B���s����%rV�@���ֺ��⥣�m�"�B�a��6����^	��f�6Q�Q�y��GP*	�Lqe>�_4j^�\��.'�������R���iY�W��h�z���g�è?�4�Gci�ۋ�����Z� 8��Lܰ� A�iKc���\�r/��x7\tC�P�]�|��uk'*��/M�QG u�G�h��/���6mz �匠D��#��NwDAy�nD��n�4���Y`�j�{���0�o�դ]��=��f�q�#�Dd#M�e�<�r��!�&�?_�T��M���;l��k�Fͯ�A�D��� ��FI9�.8v'FFm�,D�2��P����D�j��K�T�]Ä63���6�"�h�֛H��dCL�4�.a]Lm����wYRnN���ܩE5��y���zgEe�=f��a@s$�ܦ�K�QdJ00��.��w�sa�l�!��2���9�̓�\��Q{��?����GJ1�����ٞ����6�z����7�.Ӯ�ڍ�]{�YҌ��=n��e��&gZcV��U�V�Jj��h�a\<F�T"�7\����hԏ�������J	QJ�j�kQ8���N��W����W���0�H5��=��c�U�ɂGg�VX?YQb����μ�\��ۻ?L���Pji���<?��>1�C(OG��N�z�m��a�{tӿ��90��H1S�T0�?֨��x;aƭ劏K�zn��	�i�Y��~�W{�
�G�D��M��_t��"V����V.�Z�;�3pg�������h��ܗ��~Z	�	g�j��y:Q�P5�����^e�S��q��x��#�f��T<?f���/���a�bL>�Խ�	��s0(H46q�����(H'#J6	�)bڈ��8��2���C�̹���R�2)�wэ�e��fg0M�A6*�ZEQ:ug?}���lrJ�ؒ,���@���v�:w�գAG�#(V<b�	�Ӑ�M >�� ����g3�``�����������cj�-�9r7�aL�"kԀ����\��	��c|���˘!V29����1$�Է��Bu��|��g�����0����M_4H�!k�t4�i��yS��d�]���ԑ���P��P�.�/Z@����~�r<�F>�ζ)[�U��}*	[�[�#o��>��We��%l�9�`�ID��)[�$c+�rL(*T�P�6ہ��Q48�q7HRtu��:��d6�/�L�V&yG�f���m{`ii�\�X #0P���}�z�~��l )˂����*F�c10�8W*'i� ��:����U�!+�2(s?�x\�2�c���*ӼK-�l� ��Ʈ�VK �RS��N΀����D�/?9p�0C20.�4Em�:�c����O���5#�y��?G�v�R�0�/eK�W59�Q,�Ӎ�dɼS�[)���?�]���Uf�Yb8K�]����s��r�w��^z}q9��a7.��)�{��z�Mq�&,��nu�[���kB� (�ϵ��&��5�^�Q�ƈ��v�E��R⅀�8�l 2-�7d<˱*��(0��˱��1��6C�ٌ|��@Bٹ/Yˤ�Y��\{L���I��X]ίb�-�&hPf_��8Ǽ�ǎi��#@+y@/9�X��'��4K�x������-`j�ݒ���R���N�)0L�[�q���w�ĄН�#l���?���]���amw�`8���oy���ѵ�a�Iz�k��Q~ֺ%f	{ze���U�:�܍�O1�/�Л��Y���&�쒷�	Bq�?ty�#� (����x���x��N���-�)+_�D\�
�1/��s@��~�٣h&�m^s�-�����(�����@��^2�n(i��益�~�5�d���/?�[K�p!�r`���[|��WN����QS�\�����U!�*��0�Q�S��H�������隇w8E-lJ��+���t����L��~�ٱ�CSj��I�B��Uy�c��^�J�Jy����џܐrl����ߋ��e�S�̃�[����a�p��V�j�F#�RY��qN��}����'�ϓ�����n���!]sko��8Sf�>�$X}���m��W,�bͷ�.?bwM䵶Ғ���g����mF������D��6Zk�V�9�ݵ�����ڵ�Z�_[�����;����9{��d�(;2*Ο9G��f%�����ϸ֔�(��X��&^�������^�4�-������6�²\����Z��py�	����}���z3�~+.��#1zfﰭt �
ADY�k�i�#�h�,0b�	:���ۧ��(��l	�rmo�rX�� G�-oq�F����
�S�ł1O��˜���
���b�<ϡB&�A��L45s*뜪/�ԟ�`7�oꟀ]�>L����k�����Ei�-��]��c�7�etq��P%=�/��C�������N3��v��m	��)D�b�Ŏ����6�D*�*}�{�hb$����X�q����\,�ݴ����C*�~u)�b^,<���`c��1�������6��~��`����������mA��>%��������r�����j]��Re�Z���-@���C���ª4)�b��w�Uj��Ѕ���T0�51����0�\p����E�`F&��zb�/�rӣ��'�8�ް��~��y�)���������[8�ݕ�2J�{ƍ� �$��&ۃ�-�&� �L*{�{;y��r����&�q	�\"X5 ��ci�R#����>��+�Ki�;f�f��%����w�/����9f�/��O��Q=���g�U���[�A��Kзa�@B��8���!x�����`�_=,�ZIr����csl`"j�nZ�z� ���*W�p�����н'��u�^i:�,j�~Y~y	s(�5dؾE�L��Il5��?FZ"zR��z�+[�Ù�wY{\��Z^-+%Ӝ�CâG*�9�FQzivV%���!���h	��9^��n�.^�lt�G�$����F�T۰W����;�l��@H�i켜Za�.!��7J�$!e��4d��}+�w�d��K,Mձ�gˑ1{ŧ)�5�ݪ�3=�aH��ZZPV����y癛����i	��˼����� �c��B��M�G�^�&|��eI#"���f�X=)�J4"$8���l��_?���d-���o�9v�������`��Q�^����z����L�=�F҉f�f7�L�5��z�|@�w���4���G��e�)�i`�&a�K��A<�\"50m�$��q����FNȐ�F���L˶�;���C�R���p�n�ļ���$�C߆���%�ذ���P��K�'rW�P��G�/���ONv�37�&�bs�Սn��Q-���"��N�-y�A���YQ6�uO��Z���k���A�L�"����g�p��:�.�Y��(	=��G/�[�"6��PE�C�>U���v���]�C���P�bBleIQ��q�C��]��ӷ�:��\���E�X^�E�j�P|�(�> ��/FZ�f�a�aH���4kaw��X�6�L����^��3x�V�(���h]3��������pw������F�]�m����
�������;�L�I%ͮ�;[֠I���v�g������v�"�Х�����;���A��ʷ��_�g�7�,Ɨ�7����"떗�=SF�-`�?j���˴�%ߓuƜ{��ykw3P<f�����i�r�b�3����O�#�2�YNkh,�;��$V�T��!���}��ʷ鎺fq}�}����3k]킸���QF#�U������S�[��۰�a�?��Ți{S�Ӎ�4K�*�}�D��W�P�'js}�x�����L��UAL���/�^X.(\)-P��r�:X����N�]�Ew]) ��=%��I�NZ��R����IC��Fz+l��w��H�BR�P�VZB����h�nNy3�	��0�6y��g���P��Ѳ��#m2�)[,i��	��/��E�͠�f�����������[�$)ށ��#��$�=�J�k`�r��0���<5Lϛ���CIK�%u*�bo�
�='��x�J��?�0�p �� ��CT�ңM�9P\�{5�I�v@ʋ�%�I

����c�d�ßd������鴡~\�^$�`����W��s�&w���P�3�I�5�W�8�(��wu���R�T�ע:�}J�h[P�9����m�����*b*��B�0ߜ`j�s�Hu�'�`B�g'���9�˴D#��t���Z����fߎ��z�rEK�>a�'E��v���<8h�q�|�׏��K�8�4�� �/���^ν��]|����P�y�/M*��Mi���;V�����Tj��/@���ۄ��;R��smIц��p����>��}̸!���Uc�F�W��)Au%�DsƐ�> z���ά��@@�{{T�
�����~~Z��������W$/�����g�7�6�Pa
�+1iA�1��R������L�i�M(�����t��b$o��9x}�m�e���ԇr��.���>o�Q��Uئ��������M�\EeF�XRL��⩭{�*���,�xUA8䓒��{	C>�x�q��g�z��WQOH�t���G��� k,��$���C���>��y =�*���0cE��u)my��<V��	��2�n��:;�8Q}��R#��2�Â�	2�������]pST؏�sq%xX��%��!�24`��5K�!7&ݴD�/�kϘ,EFs�d�c�6����:Q���^u��'[�9P]�a8��mL�	ƥE������Ah����nT�T�Y�mr����&��w�~��H�>��sCT�&N)A�e�L4�U���o�s�V E_H���x��n��C,!ٵ�?��o�Z�B��)P�0Ļ���&Q�;jt�y����
e0�D�?t���e�M)Y"n��EY
}��u늜e�a���s�Mᬸ3
b�-Q��{cOl���x�+1�Y�@�Щu��&q*��-F��:��D0tX������ҕ�/w�©��ԺG���T��	nq/(�+��<��GCHZ��ꡃ�I��/�Vl�4��o@D�st-{�*+n�v��#*�)|h��`hǭ貯p�r�)��n��7s�]� h�.�Gl�Mo�9�&O� ����/���@d���B�F�|�%�l��>SS����M�.1z�6*�ǹ��'���gy��l��F2���0�` n$�5��2�2A`�9ޛZM�9 H�;�/>Q����ƚWI\|l�'�1_w9�#Zq#ߣ����ǥ2�7@
�#`�q�j�� �s)?�	h�(��_��K.��1�.o��Rw�a��ߢZ��EH��{�Q����|Z�2��o��{)��		������ �������P����>tv�Ј!�i�f�����GM��p���̇�W'^�����ϼ-��<�!5&�{^.�f!�s7��GFƦ��'g��]��R��z S�?�e8F� �N�;���Տ9n	Ӻ���lXz��/��څ}�U�R+�GR5@�����j�t˸'u!�ב���q6�X\�е$�i�� ��F�h�2Y����+�Ymm׉c�	L].��~�^�'�hc�1��/&^���]=��Q}�A^M�,�qgmb\��uK_{��7^�3$	^���A��fo�����
��(n��(}�zն `�����<i���æ5Y���&��*�@"PC5���=+7S�#��s0�������]�>�Ƒxds����A��UK��q�#[ҧ�����2�d��?�+�w�GV�	,�m^�C��J���c^d�%h#�>��Jؐ�i<b����	!�I$d���m��o���#b"m�Z�t�k�s>�J���R�b�"�>|��d�k�p_�}�B~2���9+]]�(wf�2�F�N��X���4�j9�����C���է�JY����)LF�{?6v����Ob�H���Ģ��?ܸ�(��&�a�`b{�wˑ�I1ģRZOB5鐨�aN� �ɻ����.ֆ G����#+( Q�XY�v�q��Ū0��3� ���<�ᓣ��?C��m�_���&$W�=�&�_X��n~�#D i.�uhC��e�D� 2��o�Q�ce��cT�@ZS��>�q��"u�Q_j"�ǖ'V6�bP o�.	.������5�%�T�(�h1f1�����=�[�!�^�D�m>x��S���K��,u��R�jr��X���p4�]��$�]ÀtL��V��m�8�}��t��?S^&d�,�#J[�.!�sU  AF�#r�PÜ����9g�w�Èmh�H�F3����r�J�v6'+�'Cb �����t7?��+���PQ�����9�����_Z=�-��D����BY9����B���35����Pԏ�|���բ�;�uS3Ϣ�7�$���RA��y�=�-���[�xK	��`��Ǌs���F�?<+�%��c�6� ����j�d��)�:��[9��K�%�-p��E�O�F�Jv>�������I���s�%�@`kX��t����;%&h�a��S	��GP�gX�=�a��l��c�8��y� Ƨ�3���:i|e��j�&S��>B	����#�E��Φ�K>1K�FC�o[;hAg�%:�!����g��LM���.��G8�Jf�ˠ�q�
�uM|f�:����Db��sh��G�N�,���Ƽ��>��S0؟�m(��Pk6C�鏛���Ɩ��p�C����'(�mr�k����j�M&��^�a�Q/�JL�x�ws���u�?�e�8���r�:�2��.��x�Ϧ^����ڒ�K�&��1��������w�V}�c�4�N+zb]�e�M�_��S;����:L��t.<&:�1�{�lͩN)�t��5��&��.BZA��2!"%��<�I��'���<Wŵ���ȇ�]���s��
9�G"L���z�(�v*�ˉj�*ZӃ�� qk�o�(�xZib#��� 5�~�dˋ	���u&
s}�2�H�`$]�t�����KH}G�|�=�z�1"��t������$φ��z-Y�.Q%��|��~ /i�wwnH���9���I�P�@�F�����^ޙc����O�l�
�:j-�߫`IC<�u�,���Ae��gؼ#��>��%�kz��^AP7Z���Ʊl���W��h���*�����^x{���;�f�B����	���(�f��W=W2��zG?uI��,�2x�PL?���ʷ7��ف����B���`F��t%��QMl�����"[�����,s��Hy
-6�ԁB@V�b��sj���/#̦�2�E &������_:�I���X������ݡ
¨-ݜ��E �Pf�3W�_���ؠ����´S⑕�GJR֐[JH��9d[�t� ]�'�k�}<P���:m4ԫn>�&�`2�O��:�R��=VR����e��)�N�r�U�ݯuPΏ���ٓ��)��M��E_�S��C۩��Φ��Qi�o*�v���qr�OΞ�Vs z��b�/Slyv6�6$�a%����%v�����`�C�郟��4=KE�]̀Y��E�Ο�"��{�x�3IU��Z"���H?\w�/�4���0"Z� �p#}�襒�Z��xx� U�Whu�s?��Cd\�~i$k��f����y9��n}$H�=٭0��&�
K]��Ȗ���E�-��y0�`�DQ�>��F��>N�\�m*��_Ҕa�Ԛ��|�N2���C���������l��|U���@ ���F�x��*q��/#�e�V��2��L�!��/9�C�o�!�/,j���(�ռ�V蓵ǅ�&p��\Uj'8]F�����ǃ;3��K ZC��~�!2 �@�QN��iq�H$�p�3ZO��H��_�ڊ����v�G�U�+鄢~�Pa�<���vv��F�)֕rSHg��p�����ħ���m������D��}�{�,ؼ�Yf}�H����r�F�wjѰ���ڛ9$�}����+���?��F�� �y�jW�����w�o3���Ѹ�3��
n�Y�ӡ�qg���H�:MS�o�B�B�N?1���z�DG�x��"yy��k:X�^j��brM�:#4I��"�7����P�8��̉�1AC��t0���Ϟ���C�e�6�촜ج9�f@]s'P��*���
y���"��aH�U"E�Yګ�>�>���# ���+��)��'��H-&�i)����V'V���ؕ+����}vRJ�,�%����@U���gCD\�n�%U����޸ -��mV��I@�a��)�Gy�"�Ņ��˸t�>����Q�k�=눹�n���q�.����+�@�nk�_��w=&� ���#'M	mU^�LO�����t@�l�)n巍����j�((�17e&ei��;q���%s�R��b�V5��T��g��7���z� �����.�e)kD��0�?���	��ԥ�$��]��I� �S+�'H����ۆBl����0RK�);S~jS������bT��~]�����퍸J�)P�`�ʾ�m�E��򅃰�߲e>s�m����\�(�������j�]U
��(3��oKN=B߁4;b�a������+���^ܻ��X`jL@q%Yԩzc��ED�[�<���b�D�H���2���ӿf�ou	�(� �<n+�i��|v��*�ёJ(�1��~�0n*r�L�Go���M������ӥ�*TI�g��}���w7Spj ��+�����rg�ƌ�ƽm�����մ1z`nY�����_�\v½�,�:�i��r f�g�I�=o[.
})0�6��{R[^^�'�3G��wg�QIü�l��y�74��v��ܘN�� �����6Zc���?�S0U�����13��NO�����f��#��+nq��6m����:[7�������{��s7zk'x�>���#���τ}Ԣ��T�٣k�+�.��Z�:�NK7�W=\�ۄ��L��N�ꗜ;�9ta^�����x�/�a��c��p����6֌��m��7][]l�k��Ԫ?ع�0�*���ӂ_!��OM�:�D:s	`�JK��ը���2�
 ���4*�8�C��}��G����է�#���1��m�{�Ot�{�B�]��}�k�<�I�ʇ�j܋	H�~�/R$Q)�Z�A��uS!7�����i�(dQFdp�&�/�L��H�`O㭙���0�JR��牱$�����I��Onq�O�^�����X��^���񚆒۳?vo���q7�4�Goh��/�@�Jfы�nw��Bu�C�C`n�g8�!1ե�ؘ`����)��d��P���J�4�i��!Q_���ΞHm���?	�r��u�a�F�X�%��(�U߽8ܡ����>���뛹�z�uNgS��Bi��PM�e#�ᄴ��4x<FB�m��$���)����\Tl�����Td<'Q������&2i���@-�ɘ(F��ş9�XY���F�W�~w�
�����4g6����s�+���|<���d��N'D1�_���K׀��D�N�'�p_�?c���/>�:F@��(�
�i@��0D��m��m?�`+�#|����7��ʟ.�U�1�����!A�͞��iy�h�ͧ�B����ϳ���M�K����9Q��e��&
���.x,jRypgoϺ<�q-	�Rug�
�
آ���A�E����;��RL	�4��;e�ѐN�@��.�<��a��n�pE<�@a4�$Gݕ�,�`��T�Ej��r�ϛh��w�{�%�TF����B�������Q�[��߼]x��4�����>���6q�l�H�w���?K�%�e�k�\��-w�ώ�e��j��3^�&���.~XÂV�{(7��+Q=�YIq�����\08�R�3a�*����~�&���gQ���"Sb�~K��Q`�蠩�s���z�Nz�2W!^�jVm�V$�� ��l���$pl�%N�H���ܛZ�0r�~"@��5��� �ݨ ���jX���_2�;[��i�s����6W\�6Y�TZT;`���"7
���{��/^LC@�CLI?�:�ShQZyBVߨ883�g�R�F����p���T4���e�������v��2��\/^����)�xT�q�ç��i�_�e����."s}'�3�h�bea�X����a$��+�ʞf���Po�Lpa3��lT���sg�_�R����T�����|,�.��-M � �.k��C�e� �f1�~��s�t�d�a�H�r�Q`���ʇ�o6�0ér��"E����u��
��M�@n��c�~�!�{0m?]Z��0����EP����ǿY������ʕ�#&����qA��:�k�s�Y.�'r���U�<	!H���vHJ�T
d��޾�L	�����9���"2���&?JZ��3�(	�ϞfJ�'���5�+�:w;�Fhݰ�zN��]]��k�gK�pː�HrB�LC@h���ڴ�v��� ��k���`�~pY�MH�%�b2�yF�� ���d�3O�K:E��n�:�V�Z�1uxy7�貁m�����Y������I���vBN�1Z�t�-��{8Qq/� �0Ĥ�f����� �ds_�3Jѽ��}"���`�X;�d�)��y���1e�������-M
*Jβ`r�'�vf252W}��1z^|�}��׉Ugrj�C�~h)s�ma,s�q��9�������;����Ӑ��m��m��:0�7	C����e�;����i�w�-��v���T6Q����7�䁧|�i��76�L��~t�^�̞��e!gȲu�Р10Α�1=@+A��{���F�D���')ɖ�����?�~Y)�F�=(f��k��Ejn�i�F����q3>����~����X�)^b�-n��x#r.i}J��� ��.k�EK����>��ؗ��%�i8��P�Q
�0�:��zu>.�����nR�Rh x��.#�`:�C&����oo��r�X���L�r��M]������4N*�w�S����A��7TA0�f����=L`�ƬW@zo)h��mw�Z7<p;w��a��.���|[w%gr@/���H�YFjy��M�M���`�&�ؗ�p�6�kUߊ��ܖu��:�>
�3H�G2�u�+���O'����K��r	���i�}����.�2`D���t=J�h"JVkJ�%`"��2��9Gנ��L�����ʳ�̅e�X2R�A	ٽk�*��d�CO����W�N2����g���I[� G��k�{ ���)娆�@�t?��1���$���[�P$���A[W71���h�x�b$J[$7S�Z؍���� [rN�R1~Q|u�>ڢ����)��I6+�᝜���O�/|a>\�A*��l2L��Z����C��Vǡ�I&�&/87^�6D��?����f�Q�u>��髮���Lm��׆��l�1�e�����<��-�_������	���l��x��U<�)��?cM�T�S�)�ժQ��|b�Z���*����\8� e�AY��-�]0o)E��r';���!��-A}?2>��SA_��z\������E�.�=tj%~��E�u�պ�y��t�]��M�����Gs:l�A��7L�N�d�h�5A�Э����ҋu����uEf!T�	ϸ�[o�RՍ���'���$�Z����]��>ib�C=��=(	:��c�
����&���l�N��z�E��bz�_x�7-��A}{DafDWK�+����\=w|����d|mp�#���l��{�����R�՚�x�5׬�e�4�"c�>���3��
�Ԫd�ƙ���RG%?�6�g��Rm Ώ,H�L�άm� H�	,�̐�-L!1����I�fu$C�
�>"
ږ-eN����ɭ7��B���X��qB�e�4����ɟ�B���ujRQ�s��U]�X��l�}.�I�Tm��4���mNxH$)#0����Ӎ�����
�ɶ>Q�dG9Z�H�6-������=�^%>��r��C��*��'�W'���ߙ���.�pT��	A!&��*��5_��\�!��˩�-�f�$B�kB]�I�V)r�R�x.�7������]�����QZL����I����1AH[f?i.��������kr��-5�ޣ�T{�3��Lm���qũ���=�s]�N�蓲ǈ��l�Zک+�ڙ�������MY[���_ܸ?����OTR+�W&^�Z�$���d}�'�]u��k��QkT"]���64�Y��}d�ZXDk�ϕ^�0�I�
�IC2J��d�(39��b�J�5�����k��������J�K�yv�*	Ф]1���w�+Lc͗9���F�B}�LMAcmK\�:�-��*���Bd�	� �d�+�F -��*^���tè*x����4] ��{~3)�'<��UH����I�W(�#A;��	���Ѽ��x�hE�qX�#WE���%`�~��y���������H+C^gKe�<��(]oT(B�-����b�����#�b��h(�TR101zt~ߜ;w�����*m�ڂ��S�h��W<&��7(�y��p���Uv�S��S������P�w�ήa$8$0��d���l2�[\��B�xASIm7�x����g\7�v�;;�oR"B}��-XxX`|Dĳ-�z㢗� er5�����p-8�.��?8�+��Y'�/��R=����T>�(6����m�<Q�SZ_	3�.�"�o��b��~�̡��0͑5]TEa���K�|x�WhОg2\��� �W{�Z>D�[�-l37R�$���B"	�FM���S�-��/��������1���	���ҳ���n����s�&#�9�k5�D�	C�M$�
Z|
�4DS�JS�BF���%�B��K��qfL���e�A�lu������S�++z ��>����UZc�iD��a
o�EBAuZ9&b܄��XAXK<:Aٴ�Psg6�C�c����G�l��j�I�+ㇳO�eҾg4�����yW���]���_��2���$ޜk�O�2%_,jMx��Ă/�/�[5D�E��+�̖,~�X�q�	�s�zp�����j"�þ7Ԩo���r(�r�	<�4��x�XT���=��&��%1��Hp����1<)�t�}�E3����mr}~���?
C҈�g� H6gR?}Đ�D1j	5A�i�_(fDO?F�5�lw�2�^���}Y�W�^�po^w0N����}oi�3��YvT9\e�F�7@U��K9�DqM�IX3�4ᾮB��Hɼ�����\�c�_�<��Y�P_(		���{�Х��w��6�I�p��gK0��a�L���u��T-���4A`��aC��Y�o
LZ���CO;P�Y������=@��w��V��8�,�=X�!E�������N����U)[�ԭ��w����J*���ċ�&�����iGh���u|��ݒ�w0!/�A۽�sk��BKΩq�w��$2�Уh��+N�uG���/�FH�)�+H]=	EN�FAI��I�Rq�	v�����z�����0S��ޟ񨀫����X�=���A7��Q�˗�L�6@�Ad���m�O>%m�
�i>B���7�(���M�a<H��Ӣ��az�!��1��z%���
h"
�

�����l�h}@�2	j|�ް8p+j�b2�j��,RT��J�7��o���oq�R��e��ȬK�HI="�� 4iu������`$��.?�\+A~�d�I<G�!!��CP�*1٣y+�<����?�'�]oƓ �)�d�
c#�̞y��Kt��R��"+B�j���l0Ḻ�+r�;]�Lf�����m{*n�8$�)��I��8Q�}�Cn0�BdT�a}���8�e���*7&�c��l�3����t3 �����N�!V�!;d}pΆz��0�mm��Aw��b6��Y����!/ư&oq42�DM���:�s�����÷v2z9��	J����zD@�n�,��5�*~�V8gW��-2���l��6���5�a4,뇑 �-qV'�#_��(�+mR�O��pz@�<���u��A)	9��,LN��PtGd�VB�Ҵ[$I�%���	�4��e��fb\l8�gz0�*�!&uP»�f/��4��pL?�*j�B=y��C�z]�W��\&7�8����i{��1j���<�ĩ-+{9s����kp��.p��c��A���{����ˣR�cɟ�ML�P�e\Y�k�1za�����b_<�Qj=8A�!��_y�g� ��m���dTC]���l<r%�+����ZG쇁r0�u�:Lˤ���_M��bF�U��M�=�]��@�ѐ�AT��sF.�irP�5>�x��������
w���c�^w�`CT!.�+��T��OT%B��ʵ��?Z����I�y�f t��[�э:ס��G#`H+�b����:�i��f���{��?b�������tk5U��?�]�߿�cl!���˽�ֱ*��v�3��xD$\�l:Q���̍�K�6��+X������̙)
��E'M�1�xZ)��5���T��%e�Y	P
�`q��u�+:7�����]���EB}O��J.�E:�q�b�x+���H[����7��-+s=N�����,G���.����f,��2;�����#X��/?�')v�3Q�Wvy�Q
F�����j�!Eˮ�˯�<jP��~�"t����cKP/���%@����iMa��@F� ��^;�����b�Vl���3^�^tS��S��p^/��j`Ix^*1��_s�!V^�C��]��� ��(6"�P��^9��|����5c�^�uS�A3]){Z�QUG�u���&��o���<��� ��)V�~�!Ӄ$@0A�����ҙK�kS�-WH����֊�@A��u���3Y����d��]�>}��ncN�ф���k"w�
 	d`g_<^�_I3�j�#�.�3�=�e���$�(����a�o��6+Å���@�8,����;��ѐ��q]��}�HO�fAͅ�I���skϦ�9�A�<#h����GK���i����(��#�?8sH�^�ӭ�^^��.�ke�-���H�{�VQc~U��5�T��ؾ>�}�h�c��	@caM���c�X�z��'�K��|�b��"z�@�^&��(�;̏��R�~�{P%�Y���ӷ�XP���[˯yd��KgP�I���t����L�뵓��ߋ��ΕbB�2f��`��Ç�f��v��Bhx��[���Je3���(�����������ӂ&cJ�"ST��aP��V�5�3���'7����obI��2Z\�����^U��ro8:�kz&Բ�g�@GV��0��\=^7��TI�ƣM�b�ta���p�A��1_��&��2����ɸƬD��d�rL<-䦥6���ÎXW�l��p
�k�3h^����9�'�	Ƌ0��̰��
�n�{��N: }6��M���b����Ń�:d*aj�~{� �m϶S�+P|��ȸUm�=�����F���ߥ��i���B��?ֆY�����zl��UW6��V���H�*�G/1&|���Z���A��k=� �oNx��Yń
��%OX�Oh|���/W��-�P��Hݟr�=�"K����O��7������=HM��x�E M#�kG5M���)�/�,O�\�;�m_�����em,���^�X�lfp�����]�<߹Mfg�h�`6�_�5��9���������z%�HX�7`�d�5UNu��<$Z����ϔm�l(��Y��?\Q���Sj����*-`z<�(��K4Ҵ����RDM�Ny�c�y�T����
��9�=ȝ��(�rE7�"� f�t��Im%��<A��Ж��×&���;���`V�������X����y'�T���N�sa%��'oو������t�f�b��O��@�X�Z<S�?��}�����Y���UEE%�����j#�Oc�h�uhK�˜����-V��^��k,-�!�hс3-�]NՒg��]�?I�X�U`n��+�6}O3��Yz"�l��'����	�_˰�ٹX��JK���%�m��F+n����<��1��ܤ���j�9���A���OJS��bö��>�x�Wv���ׯ����_� ԋ��_�e����7�J��H'B���U��iE�n '��� ��B�/r���S'11[	"7j:�y�-.3loz�ڭ.�+9e����)�H~��]�k�"�m��7��$�(��Q:C9��!�� sn��R�آ�Wl(������������q.~�$Ne`"N&�J�%�uչ��f)N)�;r�aK얷?�e��S�loK���A��m�g|�U|�x[�#t����u�ؗ���Xu:���NC����#Fcc�V�[N��%�{�3G��>Y���)h����Β'M_\|M��i����	���U\T���u������W��L�8Պʭ�CR����\k��O���a.e��f�S��2k�;�|:
���Μ%@I��F�"���揑���]{TFІ>AE;�Ŷ�_E��k�/<.���N
nt�#�r�mW�RN-�-���aΕ=�ݯ�^���!T}����=T�un�	�:�kl9��4���Z�Ed��-W�S9���x�h&#8� �����+�|���n�ߟ��psܠ)Z� GĢA-WO{���j��eѕ7�Mcm&4#q2�[�m8�Owz�ǪQ�'-��s����69mV!I^�j������'�7�)g��U_q'V���{:�+,L�n�pk�,oU����F�`�$�M��5�5�f�_�닷�T����T�v�SG�N���N����j�<�B�Ǟ	�*�ˈXP�� �D���aQ�e$s�Z|��jbht%�0���Hn_��G��i��ϧ���G��vy[�X/��е��پ���(}\s�,_~��J=rZpR[��~5Ȧ�\�K�
�W@<��;�~�˞�/�����'F�:ܪ:qMq
�pQOa��̖�V����Z�:pz,õ��vT�b|�����Մ�qP�)W��I
��Y-�l8a��ʓL�ڲZ�6�s��]w5'����6���O��CpR:�>�ژJ=�Ҕ����Y�G�,&����48���p��Z���� ��j�븴^�?�����2;�8�H�L��O5" Md�%N\\h��,�l�A�8F�W՘t�=l9�׋Z��c|��phkk��ʍm/$8еҥ'����F6���:����'�e�)I��wn�<��%��d����Q���
�$_��z�[��:�|�i%\�4�U��=?J�L�	`*���>嶪�ɍ���Oqi�jjC�o����d��������OoE�EEe@`�����jzR��i�r�|�����m$=���j���I{�c�R�R1fY�����5G��ür]�����d�I65�z5~�8/�Pl��+�+���܎����Y���^HYh�B���r��Ք�池&=	�@3����~v�-
�zis���_6� �|���k8,��b� qd��mVKSiл[��{���������pUz'@4�֕�
"v[����C>���-Us逬|�l�\�;{�.�$��X'��`�9lQU]��{X�Vn����^���Sp�'���jA��B��֔�g+`
+�������c�R�?\8F_R>�����[}�HDݛ��Eb��������`��Dbc4rjF�5����@>�Ū��4�Q���D[4�!�%�_}��'���LH~��l�������&$��#�\��Zuix�v�!-6�<[j±O��h ���7�Ї���ߥ���a9+�('�.��̦
�3�:�uG���G��I�,���o�v_��~�G����Ku ��	2�)�pH�Z{�U<&����>bؓ����
cd6������0��7j��+cs��5�)b<ӈH��x?@ޤ*������p|I��t@�7A.���p�� �RI���lJM~M�D{]��Ov](��=��LR�$5�]9���@���p�dY�ى��X�9���
:m�;��������X���"�Ri݅�[��W��z�1![�0��YG<��f�ZnTc�4�]j��SFb9q�,���.�	|��Byz����`9U !P�-i�1��~?���j����d���.�Q4"IM�Q�jJ8NR>H$�)�@�gy�eĦ/���9F��!�!������6T͔#	U�N�LS�Q����ۖ�8��� �ܤ�9�r�a���_ܜ�����{0 n������G�i��(-d:r����?y'�%��h��ac��gCy��;�s`:8n1 �u�p@���',��ec�M��r�
��X.��q��"��0B���L,nk�H�>��OQ�T�b	�-��*)z|�P��u+�Ċe:��!/K0�Ɓ�ؼ� �N�tk��v�h��h��)�`�[���x�o�����9�4�d/XɮZ���$bXoV��� 97ȑ.�c��)��Od �[�r��Z'ߵ����gۉ�{B���~�D�쫶j���O�s����"�����G����T�,N%�T�SY��s�7�A��t�.��Ts�~��H����j������(���6SP�C��`KK�G����i`G9TZ�	ܯ%���܋��QJ/�ᇷ-��1. 8���A�,g����ծZnt����a`[�>}��"Y�����?�Qw칥��Y��k����zl�ya�m�t�@�ܲ����A�Ȏξ=��{΂�yEӠ�A��䰥��;z���7��yEn_����eI��t��c��]R;x֑�:�4k{��	�&dt��H4�-p���,KˍAF�M7B8U�J�޳74�I(�z�-cQ�����C�%��N���j�9�J�WZ_;�D�$ecK��?5�7�!~xqs.;�^�f��1IM%)8�mW��Ԛ�Xܩ�(Apf9Dem�}z:��ӳ|�K���X -Q�D`$N�X ������!^��dM��?t?KN7��݃?�iB5��X�0(nB:Y��K�d�`�{��3�R�GHQ����Wur@P�e�_�5$Z�@Ip�F�P�{���<ݜ����P�j��{)���a83z����I�B�����#��#�$}�)�q�2�=*��8v8�h^�biq��W�bis�R�BK�k.� ˼�-��sqD��C�"5�����Z�UP�S=��rs�T��$aNCet� ��g�fn�e�Ӝ�,@�v����z?��;O�7�@������h7��$h����+�n	W82�W���Ȳ��a<�<��d�N�t�ǯ�"M��a��~4|3$.8��(Q�k�W;��-����h@4�;Q`�ij�.����Fx��r>sgpp��? ж>@]<枩�P5��*µ�ȲnP�I�2nFH�{�[��:����|Ipg���T57`���F*H%"�<����.g�����PZ
�Ɓ�� ºČ*��b��W-v����+�am����}����"�c"��F����v��ۻ���]�����|����}[�؜���_�6��Cp�¬TǙ�0<�>�C�׶���ۊE!wNU���g4c���#��>
E�Q��ޔ��d���R�~W�����S��C�4�J-�j]�e'����*��+ᾟ������TM������}@9����ˎ�3b��� �I��5&�͡X�}cx����<'��/H���u��(&P��3�v�)�Ү�nd���U��猭i�M/��J�A�ֺ{�0E$�܌���8.��1ez��
� �d8?��\'��;�4L�N{Xp��o�f�ޑ=��ץ�	��j̧
���+���	���.�	0Տ��R�`\��W�^T�f�_� �b�!�w����*a���pYhM��A!�����pn��3�T7����2����	|P娂$�u�Is��V����]����Z&}�`^�7��m�o�O�8��k��tCcz�P-��=33�ܢ��ؕ��i���B��`�r������(���t�(̞R;�֕��bp:>0����>�+��$ƞ�G�H�#�5�i�r�����Q�#<;�.u��j"�
���	��fz���r>�`�Xg�XJ>��"�B�����A����(+~O"�
�Y"Q.�P��_����5��'Ā]�[�/�����[R/�E8��L�{�am8��e&E�ʔ9�7�?z?h�J����m�2�m^W>u\O_��g!��т��0�~XzA��Z��+��d)�}v�+����;�Yab"B��b��k���JL߱�d��U�qBUo*�Cg��!,@�[�q�����T� dōV�0��ʽ�>���X�!Z��m�Y��{��|���b��S�ʌ�)+��1ԕ�U_dw�n�{J�B5s%n��t�&���j4�ׅ`�@Ǻc}�9���WP��c��k��ֿY*���V�"��aT����,vk��~�Cg�k9f�w��)\vxT���:ӕ^�'�� ��}+��9X���Fm�O�ȴ��w��O)�>-A%��T���%�c��au�������X'�@c�+,�����Q�n�2�0	gdSb�vm7y�un�L�|ũ�f-��)���y/�hR]�&�9C��y/�O!D��4�w�>BS��x�żlx�݈���DB���	g�$_�g�g-TH��Bݠ�;�n�'��L�=����^���D�L�s�K���#���+�aՂ �3����&\��ʀf�'�k̆?���X���l�T����j�St�UD��P#f`;��cp�L-�g�������"Y`-��o�O����,�7�|�� �+PT"�:�m����0 ��:l"�0��k��s0>3e#k��T|��Wg�|}dO�����*��)�ɢ�L�Zک6[�b���xd����u������kdR�d^tV�F�O ��M����ϑ��tP-�f�B��u�A��'���٫�yh8���Ɇ���G@��^gJ���p�͓��c��(	i'[:B�x�p@���O}$s��ؑS0<��-[��$s���	h���P���b�P6� ]����}���>?������x5c�2�w��Tx�������p�-s�,E�����M�u�u4�E��ﾊ25�Q+Q�L�>��w�:X�E��i���*��qDA�����������A�N�}DSNBŀH������׈}���<�K�����Ϭp%�`ج���� �j��⭺���T�)���	=Z-�%�I{0V%�=��y�:u��\H�P���#�Mm�:e�����V�誠��E��"h��`V3��>{�E��_0v�*z�iZO� �������Ӽ����k���WH��D|
Y]�����a�+m�H�l|r��~dҤ�p]V:_D����Ab�ߐwR���(���kE
O8G�[��]���ׅ�Z�XES����X�<o�\�����(,Q��9�~W�Ŷf�>*�7�XuUW_��M�;�/�a��[J�� k5ۙ���M�52�lEV�*
��e����^,��ͨSQ����~z���<�"]�����~��n�����dJ�2���fF��<��w�QpHڣ(H77'�ݘ{��s�!�����%/�������d���O�V�5�沐�'R�&�s4��Ts�e طd$9
5V�Iod�{5����0�;�*��_��mE维��	$���H�}�p�4U)�#���QujH��|�$�=��i
���ރ7�X�g.Lx=Xz.@�.�#�3�|P�����10���|Y@�TcRn���ڎc�ML���_H�Yٺ��@jT������n_Ͷ�5�b�P�U�m�\`�~�M"�������c�j#'ü�}Α��hxlTމ���:H�O�m{(M`��R��mx(��tY�ͮ+�v�z4���f� Z��?�-
� �
L.j��s�����Pw���B���5�nB���DiǍsie��-j�������� �������[�F����TW+���?RIצAB`��b�ys�����,J����<OBŮ�|[>8��-�����Ot�u�Z��5c\˩y2	�=�^QP9Mı3Nܑ)̌�P�\2��ës|S�&��WJ���
�����0U���*�Z/���(X� �"m
���֛9GJ�գ`�)��g-���h	�ra3^�e��c)�Ϝ���]�;kMV���
���>~す�xW�65�eUB�[&RX���OW�I���]g�i�)�xȭ��vKr����& �9SY�տ׭_M�k��[�n��� �#�	��5�����$G7ȿd�:�x+�H}hS��o�BKK
��r{�J�1�>y����s��,���4���(u
�s"C�~��MH��Q��U��p�2���3UN�&�{�ݯ����ȷ�ʥ����=��K�� ~'�m���Q|����9�0�z�tG��]�j�l`�tT�a�`��)���^�o�\�*~��g0��֞@�~�3 5��U�����}�ǃ�K���n@^��2�Q�v.W��	P�JO�ENNP�Dx�8��=�	(�@���N���O�$y&9�Bi��Ӥ�v?�7X���ށt�-k��#"�n�d�j'h�XہFE��2��=�����s9U��FǯG�ՂU�X:�Ȩ@�f�_�T�j}�S�>�Z����4 �d�7���MOoc�ol'Y��1���<m?���D�JdoK&8�94�8%��)9��طn�3,M!~�-�S�Ā���mH�M��{RD� �`����<Yrl��@���c��it�U2 C��"���d؁(�|��}��;�.kSּ�LY�f-�oS��3f's���[��Y_ Vk#�Ia �N�^����H�'R]��򻀇ƂqO䖑��Ҁ���N��@�V����9)dPj�9��ˋ����6���z�_�X��>�w��W�����ERH-]{ty�kZc"#԰*�^b�q[apo(�9��kz������'�[Ä�����{q�h���nST����q��N.k����>qw>A��iol�vI���q�������;���ŉN��s���3�y���|�ՃB@�NY��볯AF��h5=*n0"�B������	�4�IV��s_�� �6KL��AI�y+[Ȟ즡�ch���ԣ֟�o�uW&ؙ�Z� u�Ѽ�G"8L$��Dg�]���뵮�:+՘O<Dz�,>@����XO��C��"$�)�V3��
5zx����d@��R��Vx�q�" �bw��xM �Wc�:��
 ��a�T��m��%M���7�) �����A$ ��bC�#	m����*�Y��3� �����w�}XL���T�w�6�	(�tr�dY�EWe#K�@Ln�$��zc��c&���vZ���˦۬�o�'K&��~�o3r��ر�r ?����.}8#�&�r�]��-� e�0�R�Q~��r�G������o#[��Dj�[l�����I�=�Α���~Y��"�ڱ�%"�Q�1��F��=�r/-L��-wi�Q�-5]w{��̩�i���R��
�I���(��!|��DW���\4fP�!|2d�'�&�����[�I���X���Ź�#�9�Vj��H�׶hN'֑�l�s�G�΅�,����09V�0��D�d	A,�
Ŀ���]݅^��F��_B�����M��TUln~*�bXϐ��ʎVzd 6�~����1��o��1���*�0�}�C��5�(���b�H7:h��4�i��J�R���m��`*�����4ĲS�5r�mL#G��N��p��񬼷�E�/G�&x�^������=yc0�3�=ґ���a2Dٚ��22�C ɫv��s�~����v�R��Sm��f�md������6����
w](K?\ƍ��8ǔ�&Lmp�}�%��w��Ǘ�M�B���»�0��^/�K�ly}`�W
u;����Ηv�����hM��t�n�:�����y�a�'`��!��h���?a9�B8���y�،D�ט��ϙrQ�;	�lкx���h�E�y���c���K.}�;������gX�<�z$�� a�<�������Y娜��d�c���µG�k��c`�N�@Tt]�^%IBd4�EC��y���j�r�׫m�+;]i�%�T���i�*���k���k��o�/3����;F�N�<�WW�������{o���)7TF�>���zs�T��K�N"�f���%u��N�]FR}2� ך��QU�^��}Q��񤴚`C��S��h���'%~�+dJ<D(�\���w�2�}`Jɴ��.��=���2r�QG��	���P�(0�RI���ƻ�hr0�!1(j0uG��T�Tj-�Z��OVxC�u�����.o.�z���u\��&�g[`:$_�J�i8�ӄ[�VJy�EE��p0�l�mB�� o�أ��8�7}���EE�dR`d�R�T�$ﯝkȾ�C�V��eD|�����﫹7F�Q��d�WB��^�4�,[�m2�öU��XkL=�G�/o�]6�s�A�v�������n�B��.���6�]
���������z�9b*��r^�g������o��X�㗹��"��J ����m��xn���뇴���y���˗��N5OH�t�j���x�Mf�|:�?�Ƹ���/:����ў?ؓ���E#��/57�7ɔ2!L��I�8m�U�O��8�Rs�6-|5;ϥjG5�1�o�W1K�a��f�������/Ly����ճ�W�B�T��V��.D��J���i
6-�hVL�'��O1��^�U؀���O	»̵#�~kyj"��?y�+
��Y�8�hdX%N��.mv��ZE��+��-��Y����'�Xg���qn�{L��n���8�m,��g�A������L�E��|n��Չ$����^(=�Rزf���}�\aވe�?�;ͥ=+�sn(-{i���\꟰���X.��@�~��oz=����v=���]M�N5����Ҳ��O�E��=d�`moq��r������G��[���)���j��z:'���vg6�;-�D��>��`~��%z|��o|	���a'S\���n�Ǽ
�,I`ɳQ2�_�Y�j;�v5R��V�_Q;�3���`�Q���R=�%7�OBh��%�Tj�ې&]�1=�1ʗa_�f�����hחd�3fIX3a
Q���FЃ���#lS�)`�8zU(}jEbT���L.�O=>�#��N���x�F��Ǳ���yW�$ Gl�S�p�7�&���\a�:����~ն}&&�W�"�M3�n,�$��X��\⓷bZT�~/?������E�/��f��5_��M��
�>K~0��o�DQ�k �˵�P,8�܃d����6Qr�~�m�`<z)��wq��6���V�Wk�����-]�eN�/�����hr�h��}Q}&fu:v�ނ��yޙ��`�}:�mA"5	W����iÎ�`'KaLn���Eh�B��@� �2���;��3u����<x��
a��)/i`�0ӿxϡ���_B�=���5�oB�����7��d�j��6_@5ѽ��H�}^f���L����֪zG�r��33�ήb7��Q���|�MD��	u1��X�ό֑���	K���b����"�^K���P��Mf=�:��D��cZ���-�� �N�ȃ�?��W>�'�Ndx8����{�ƹ�FZ��+疀�k�:?o�v�SW�i����L��.�.�RR�"Y��sN�R&:&��֗a�o��|,�*-�"��8Պ!�x��U�JM���cz�>�YYx�L�X)�cum@+Ʒ	�bk����fNd��"7׮r��|��A/F��U���P��S���6HZ���Gj��@	����?�P�"P7Yd֤�V���p9��j q��� �~}�Zŧ�����*��ҳ��yx ��u���MPx��a�3�{m�/c���a��I2�0�.]D3�ٿZ^w3Gʙ?���(5w�����^R���:��úP*��[	�zD=09�곽~�*9�7|�3�j���t;��lғ��_��N%�̞AJt&7�?��0�
{,����v�*�c��D[����VI��_Z3�Z��m?�(����;tqHm�\ɵ��w�<li�S�P����X*�"dz�|�(�u����e`n��{�&��\�C�L\�{�a+t8ͣt��)�~'mt�7+������!�+�,�(�kר�b�"�=�}�0F�!`wܵ��)\G.�����.���Z����c��EP

�<�EM�;H-p}�����C�rF�t�" �w|�#H��?"��Y��?���w��_[P%�OY��M�w��!�ʼ9�����4�)�.�E��<���l�iK�h�/+z����h��'1I�;�*∊j��휠:���1l��RnA?��n�����ñ�i ~'�L�=#O�t���P�)�4q F�������֮�j[�ʌ�1Y�%tY*�.����Aԙt+���j��d�F^�׆�c�j��G�����Jn�VT9u!8f��۽;��"�,�[�W3'�:/@�WHp@fn<� c�/[��c�ek�2w�s��Gi��F؟�@��s���t�&�s��+��s�/�W52wޤ8%'�xwsm!�a�I`��c@�OӅ+�B͔Y��4�9y5��!V�hק��0��Ga-X�N�@�߃s���"�?�@Q��e�I�A�8ЬL�|����i�l�#9� 葇}5%�m%G" V�{B��:$���Z��]��/�
����/J� �Y����c1:�|�� ������
����Zڳĕ笥h��MQ��\���"�����u��o�Ɂ���ӲYzEI�ݠU�8���]�d���J �nSV�9ֿ���n<�J����]�`��!qɑh�A!���r���	()S����{٢8Jr.D����@W���\�炷��՞^�L��h��)M�R���v�r���1�u��T�6��/3�h�5�����V�Ld��[M1`Z+	 z�=�bN�R��pv����Ұ�q�Po�b���[�a�0�a�<i{y����MF������ߩtv�����w��[����54~!<w����WSd�sn�y��}-T"BY�˔5	�f���b�e3hn'���~����ӆ�(�tp��%��L�
"�S=��jgF��0�3��Bq�G�
hONAܼ��Cô�K"ɠr�D��$�䋚kqȝ��+4���IdR�"��X$������j��݁ӤWb0�,0���!iT�]��	��@$;?'��q��u��m{q�	����B�f�\�TC>�?x�Y�x�
��-Em"���)I�;�(Z�㋕�ڄ�f�P�p� =-�wE�W��Xz=�:��P����i���YaS檧��w{:j�k�'p0}��A�4�jN�%}ܢ�%�qV�Qm24���}#U��hHc����|�;Ʌ��\"x��a�����9�W��$��*��D�CC��QH~
c1\�Bi�����-恗�k����,��k�tWs�4�n
�0
@��_g�.L.焚R�����SH���	�W̜����X��@	}�E4��5�B3�'�]�c5�p���A�Pڬ��N�%v�F��V���{����Sfj-΋���"s�@�Y��8� 