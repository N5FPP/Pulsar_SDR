��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv <��Ɣ�����hd��� *~b�<��G4�aY�M�z31�5s�Ԑ�s��
:���j���w�BĠ�9f�i��?!�B,�PAuO2ua�a�{��m	RK��̓��<��e?�2��ֺ��^��}J� 0-C�"��h%��p�V�}yKn�G2��}k�[ﾗ ~�]���53��QRs�Z�80�"a���~�%>J���v/D%�l2l�f��*8��^�Z�2yHd�Ɏ��/�Y\5��6!7�ؚ�w�T����l�CThw��mk�:�P<�u�,_��{�Jc�K(^w�����.d��b1?Բ?�p�i֙.&�]lҴθ��#a��Y��=�;ŗ!;T���)Q��֪�Bc:@�#���2��H�ͽi�'���"��N� sN��V��8Rx�g�y3v�K�������H���O�i@R�|Ygt��n�0�Da�	��@e?��v���_G�� �x�F�m�1 \a=�V���[��Qw!�)�ϟy�s���s�"%]ߜ�كq�M/?=hՆ�#����w��3�2MI�e��^�O��\����s��T�~ZpA���W���!����1�ʣ�N8G��>��y��Pz2���V'؍Ǻ��Tx���?B�=C��u��e>x��Dx��;ڏ����ϛ�c��1�}(SIG�߫��8���T��?E=v���'r�5�(��Hp���K]��h,�*w�A����X��%+Aj��nF	����19����+ˇ�,A.�d�
 �Vۤ� ��H��!�?�;lh���gcc��nk�#z���I5}���D>�D"��&}��c5�C�p�!���h��H`SR ����{�����d{���JcN����s��^��<x����3j;��T�T4J}��μ�<;�U5E��Z�btrRX��F,gB"�Q_B��1�V��л����q%�B��U�y�HHa�(���빪@m���a��� ��ƴ{0����6�-�2ԕh�����<���Pz�#��q�O9�Qn}l6ssY'P6=�Yݠ@����\}@���~a�B�yR��G+S��2��9�OBȣ��^S��H
�K�����MІ�|��RѿS��DJ���n>pիJ�k��O��:���Ӵ���t�w�0�+iz�=kS��X�:���f��hp��1W9�H��'�[1����9)�/8i�a��=���"���Ϲ~�
@��1o(��+b~�8�{��z����c������ێ�_��sؿj��^�ג�E�W7��]ʡEY&�����HE��V�`*������Ɋ����,<��g��k���>����"��%d�^�G��D������ǎf�i�� ��a���?̼���N[ߊ�5����¡q�3�GXIr�&l��aC�������(�%��QR���@c~+-k�\gJ��#���qF�c�[�_*��.�d��ɛ�o�?�e�8��x��0�-6"��dn��Z�gaR"����y�	�E94�����#���S7��EXʵ�%��.[3;�C \"�=i�1��I��'�|I.e�#2 c�E8>3��(T��F+��?����ר:���>6��M�s��/��l4_�����K�.nt�>UK����*D%.$��}���;���Ү4+�ПQ(���>�����a痭�6m�=R��4+̰]�G�M��#��$F������O��:�[������y_�:�X�|'���{��"im��{de�R���)nk�f9H
f��1Y4YI��1ʚ�f�T������:��lSd��~�,��S�=���)��6���?��2&j�/uh��[;0��@ʤ�qo��~b�@��N�a�*o�t7��
�0b _!�)��*6?n~�2꼢��Qn;�_��(��¾@�R(�w�^������$��i	�o���ɟ���P����yp��'�c�U�Fn�o��Je�=E��m���ȗm�;���(
!ꓩd�͛�8 ���;ro���٦oR�S�����w���`�<��A�5u�N�8PU�i�������><�~�a�'��d��#�8[w�pޠ؍D�a��*�B��_n�K�U�14�����|�����P���0�~s}�>d/8+���/7AE�MĻ�ҁ���2^�j��� >��+EԄ��Q�+�������n=�Y��,d5w�$����D�?�#�&�n�������T��3G��;�6].h� Z�?��x�HB����K\�@�uxbF��Q��8�Aш�r���uG�\E�#{�=���M��N���C��\(�����4t���9���!�k���C~>Ъ��pJ�9��IF__Pmi�i�&���P^��<t�h�c�q�,'����$��>4"@��čɕ����Kη�d�ӲU� �Q�5p[������
�A�d��w��p���T��p�&H�1m�|c���2m����o�d9�5j�jj3/������{�Y;��WS��'�Fǡ>�SC��b���~�NC�����&�5� ���쵈hD߂��e�̉|��`+�9]�����0Ct�8S DkbbU]��[�1f=Ȅy)fW���Ϗ��\�O^	Ҳ�m(ay~�ņ��w+@h5E�1��37u�V?���^����T��l�g�^��k!�m�Mc<��)z�<)���X\W�i�ߦ�|���S�B�<qx�_ߝ����>
>���l�fcL�ÉcOw���ǽ�<���mŊ�4XZ�`�*��yq��3#�n�����i������|o>�-���M�DT���fr�e�G ���ƠE�:ce�������P\a˶�D8�����Pp	{཯�D�u�M�xB*Rx4�O(�|>��~~[L��{6���X
$�U9�����߱}��]^���5���A����Gp
*�
�ϑ��z|2p��<�'���T�܊�x�7E��c���o��rO�[U������f�R��7yԹ���5!ULA�b=ʒ�=b��V�fR�39<Jwߋ�`���Z&�U{$�]6��A�̶��)< ��?:�S���C�]�,;7r��4��\H�3_#^̠�-�^ H�O_�a�k1���s;���/K�2�YIY�Å8+ci��N���N�u
�� �fT�jO��Ӳ��4g�sS�!(S��^��ڷ���p���t��5��g���8~�Hյ�{h^�i���8a��aI��\�b9�n#J�V��<��%�UP!����|�w�Є���v�7�k�,�q��$��y�/�:ks�-�.>;Q����?DHG	�1�x�Cv��ϔ�8�^��[���Yh>�A[� ���S/��0]ms԰|�S�|[�_:Q͉�̎����g�`i��uΩi�h�Fk|���7�ͰBB���a���,T�����"�%Pؽ(�uj��.�D�Nh��&�=�͈��Y�u�T$h�θ�wB:|Q5oH_}�M��br�䜲�U[CN'!����u���=�S[H��W�ѤV,L?1�b��Ș����?�{?���	!� +C�=�̊�o��N��Nc[dH��z�H� �y+��l���֘�E�F����`Q����Ǧ&_�RRQ����S`F:�D������9�}��X7�I�6��Iq����?gYtj�a���l`��G�*7}9���ST<��v�r���k;�Ռ`���|W�� %��B��T��s�&.���U'�����19�"o�'zUi;�77�̿����<�獛:^2�����L��M���[��g\)?L� �7��Gs�-h�A��(2�+��Y��Ћ,������9C	�?%��}���JY��-����+��O�B����N>t���4���'�ˑ,Sa,��@,��_u��˸�����&��m�8(�xM"�;��<?r��J�������N'P�qj����>3���{C>1V��1
�x���l*g���Sk&`��l�z�ʍ�#3_K���٥֭P�ҭly�&K~�iw�����n�M"�6����eF��2v${z��?��V��5^M$�n|Og�l��g26���|u�#��D��a�1���B������/:�k�(����H	`P���*�@�j���E�q%{��.ڲ>�"��M�4Ƃ�s�r'����unXh2?���u����+����=Mfs8�k���a�'����&(ex�F��Xk�N���E�.����9�1u!��ж�9N�u$n��*� 4��L�qN��+��9�O?�.0�+� /�&���n�E7>Q�v���	��~ ��j^��{��k2,t�Mj��yk��=�ʺ�r��P],0�� �=ǃ��lE�ԧNJ�쁔�"̯&I0?D|�2.��]ш�-�7F�'��3�o�Dn�c�Fv�Y�eP�~�_���("L���)�
M2�$I;�w#����%6�s} \�hJ�7�]<�}��sʓG�O�"���R���N����<��C�F��Y��c�+�6݆;UCɒCw��!�G�;0O��82
�e<h�8���9�����T�Ai�&���coW�e�r�M"t����T~�^cj Cg�J����Ðޡ�ȭ ���s��o����G��KK�M���WG�q㘜N=���Z��$��3^�M��]*5W�+�(3�g�Q��̿YA�����$CGP��r �m���J~�r�ƾ���ua�;	�%������s�3�c`��թ�Z����
��^�؉��l滴�zr���+7\�h�E8�%�
ZW ����N'�^2��3�'"M��eP���ZXm�U|��&1Ǆ��:���n%�E�@�
ΰ}(o/�"�!����Mv�9�3'#�1鵣"�v��� M�q�����=��B�W)O�4�n���~���t��7������}�/~*.�&ڌ�T�!��#jP��j���B��l�S��d��b��U�İ�~�\K�_o��~];���<n�Nm�e�%:p�3񽋉/p���P섺�v��*/�<���PD�-ձ�.㊨����_R7�I�e�%*y���$)��L՘��3	*&�߷���eL�<�F��#�����H��-�	���@�7�T��F�5�#CeC~�f=���Ct~/��ys�&��\U�Q�_F��},zu�vϗ�����E�X�8hm��?�����!�J�J�w �8�Bz��*��`���]IM���x�bu�G�I����Y�G�s�X���7�V�����bP���0�ص�?˕;�nV��.8���YM����iV�;�Z-�ET�X�:e(��Rv�,����l2��@z��G~�f`?]C��b��7��G]$o�N�Ryl��B���7pT�/B���;�n�]u3L+�����n*ؚ�T�㯢��A��ϣ[�8��&�� X
���X���+^�3nqk�C�9�qkбAL��L�L�Vf�d��"�����P^�����2��߯��Q��M��ؤU/%\Y=n(P	�����B��k�d(��VH2��:����c��#k*H����8�Dw)�H��l��\�~�N��zT��,�W�y^Ʊ���Z-k�b����X|����ˢ�)/q�:v�q߶ƞ��w5 ܻ4w3t�D�1���%:�|`��U��oٞ���;�T$��ueG���m�[�� Wo!���Ѭ��#wS�,�X�}?r��A��M̦%9����������b5�
�|Y�ݽ�k�&y�֊���,R�����Hj�J ��$�QíBogb�(d�e(΀/v��B����]G2�~��ȼ,왆W|y`Ϳ�g�$4*es��������v��)��0����%�<��ɿ~�_��?�cC-�C�uh�t�>�ÿ�� ϊ�JQ7���ڰ���'��c����A�Y�E@R�b��m��	oqҏ]"m��|��-�����j���!��K KRR�&J���Tțjh�=@:;�7��g ����b�3@;,a�S$l�j�mT�L��tjM�4�y�TF�rm��@��Z������ŧH2�[�o~[�`�l������?��[�զ�S�+�A>V��?��:,����ԩp�d��=eH�_�q�V3V��Q{�h7�\hL�"���L��m���v�V�u��I-z�R������)tV��@����6�Fy�SF��y�m�{@�������=�^�}z]��\��ܠ�l��c�D�1P�lb<kͻ��Y{q��ovlK�#�-�G�,�3Q�%F�i^I��s���Nԃ�Ind����؀ՔZ��L�?��f��e���1(<�\
!hl��X>F�+mD漝�wi�E%[�CjRS����	D]4v+O*0X��]n����Y�.��d\�4�#�Z�(��W�W�Z����g���� ��R{/�S�(�h���P�ďϱ���rk7��W�{��3\���(ŏ
���oJ:l�0����"�LR����{�jJ-(��3;B~�Q����"_���l�ǉ�\h�a�� �+�/j*U+\ U�Ž���q�pJ90Oِ�ͼ�*b�țY��:�p<���ދK=y��z����d���9�d�<���6F}/;�7�P"=>�}mA�>?�GlL�l�D����
�V��-L��Ө����8_�n��jg�� 6ϼ��D!�)!E6��'�5�U�M��D�c��-�
�'����cH��*��R�vhn	�;���
��ՁK���V�����q�ű3�֓8��g�~P~11у�����u<��Ŝ��%���v�����l�Y�5� �_�;����{��$ׂ�l ٌ/v���,����|�Pc$U�9���O�jm���� �ȹѰŇ�|(j��ޟ�c ���� �k P[ 4�z���Q�m#��� ��ýʔ����@oH�
՝��1v��DaB\8Z�1/v-�:N�\��Hpau���-�G����� [ ��P����a�3������^^�d�O�l�U�To�+pbH���D���"/Ȳr�!����!՚�����.t���'�)o�R�'7p|����(0ۭ�g����D�e�J8
���'�wX)l��	�	��Oyx,_�E6���d��q�'���?��r�/2F����s�T��=�N$Ey|oJP��A}<�4L;y�H��sF�+�J�;���y��y��>��0���A4��m�����fK�d�_
%ݷ���iE����=.);50��bJ1��#����&S�ZQb�zfֈ}�AZz}zJ~�8Qi�˾5�7�N �&�k̆apݠ���[��	�>ߙߥ?z���O���,���h�)�c �Y2\�dy�R����Y6�zyĻl��r�9�8.���d�������?���L�ED�u+�ݟS��Mׇ�4��g�/�km#�r#R���!��4�+����u�y��1R������)�h�|�c��R��2T�CY"������.�\��ɺb:��[�����q9y�V��*LR��C^���Ō^�jr<�}���|z�3��X��ؓZ[�ˀ0��0=�ׯN��y����3{p�D��d0z,��K�\|xd/�l+�0i��~V�~D�N�}�^�.�J�њO�:3��Q�ڡ��Ç=A埍id Iug�%�{(gϙ`����2�p��/���-l��r���j��y4`Ǧ��!H��Z�%!�5���a���,X� ,�(*\�*v׸�2�R�U��s�3o�D�w�����~[�
j@@���v��(k��w��k!���BT^Y��:5��#E�$�z��y<L�z��;A��"E��� �,۝�'W��.Z�&Ǹ?\�v�r���RL�jB�@��s��]��bh3��Vߛ�	43l~�5�9��mm���:U.p�rΘ����?J���A������>�"���&l$$Q���ϲ��~{|��֎�o��a����X5upFWx"�*��&�͉5:���Cvs #�Ķ���Ǖ��*�&��=y��ZyRXR;�N,|	�HY�*�*v��P2Q���}��V�� \G��E��ʚЌIfa��Z��5��@��R�o�q�҃!��r�@�vG��ؼ6��L}q�bf�;���䲅;y�M5�QF*]&�~+�r�?�
C��e��3���io�M��+��rVwC�aWX�s�朰��<=���j>n~�����c� Kכ���<]�2���mU\I�|� ����H��J6���+�O��J�� �>�
�%$�bG�}Pd�[D��π�˨b�4kv��:|��Eּ�f�5 {�<�V�i�HeI�(;iBmL��HA���O��(�i��O[���+����9�o�g�Tg��R��,3wu�8����^�2�#h_���p����ʖ"
�Q�5=Yo�����8űK�r �w#ƒ���#>��)I1N����9J"ĩ�«F���-d}خ��#����T;3<q�'E@{��X�C��4�rŎQFA�kX.��Jը�X���%�,����Jɖf��{��)lϮ��w���&�tP ���<��gG;�ǹ�m2�;�O���0��g��(,��U��.�w�pۡ�*�$����Fk�r���4�����:��Y�zҳRco�f9%XrhfB{[b��L\�# �}*y'܁�J�Jsj�n|�B��b�g�o��P��?��IN(�,�����<�X��ds���ފJ����k��b��8
���T��R�By�)�\a�BDQ}D�bA� ڰ0e�p(���$ ���F�{7����U��]�%0*Ѷ�j]�2�!Xv��8���������2���x�����USF"Ն��bZ�j˰��4�ů�h6��r���!��R��Б\����ԭ`�0���'�
�Ci��8�^&�k���s�����tN<{|��ɥ�+']�QN�]�d�C� ����Y�!� Q�a~<������2t��6flD9I'�˹�T9S�[�а��i}Y�U�L���^���v�x)^��\Tu�zq��f�����s$Ҵ�=ȶ����b� %��b�Α_HУ6N[�v7F�1���X��KޓAR>a�9��'��
m��C�)4sT�J�?=G�]�]��咻�1>Uy0ߺf1f����ƀ��%��6y�,�kk-3h��5)�͖��b����ё���
�V�+aO� �U y���^~��ҩ�>xa��.�EԼ��zmv~w��'��/�͞�5�_'(R20RHM�.h�3>'�p��'�\Op�%>����:%�V����b�rJt0zZi8�ٜ�%�o8.�rF����.�N���%e���o�-TaD�(�c_���BP��ͩ��L��_��>������&W"��%�:�GNd`q]j�"����B��\�¼����1�f�+�z�×/ᝌw3r�L����Y��`Z��&���eI���`Ť;�Xp5֖:�v�Xȟ�H��%�����q����0c&��������w�kC*��g.�P
���r����?8���8<�cи�_��)�a�%ډ���_3]>�9�8*w�m�sv�p֬�>��OOi���B"9��j�
��+}p���&��8�,k?S
k&ȹ���;X/㨘��v2G�E�^	��J�ϱp݂.}Ռ���\������W�>B4�PsE�-%�ڹ:�N-I$
T4i�ԁ�r}�0ڔ����!��R��;�R�
`8�g�I�=,��]�{=IT�x�Qf������%���S]Qʼo�B�9�U`��^�/�Q;1N^�&3�6f²f���%F�X/`^F;�O��GH�����XI��^�)���}�����U�țr���zB��#��I*Ϙ�P��m+&��Ǣ�J;��^�dx���B���G�FĩJGQ�<gp��eRq�����P���r��8G3�"�$F�K�ǆ�9?��y����q}>
��]��ؑv���\����T���8>F
��{n�X-j��D|��`�FI�*��dy�0�h�j�o4�MUC��{<�7��'嘚5i�ۂ'���J�Iu���Ty7P��8L����5B˔j��,����vĹ�>��<�C�ށ��G�J��0�r@�?q�o������VG��w���(���N�)�` �&iƫ@i~´����^��Ϣ%o~��V��t��f7yTHP~(e�9?s��#��~�������dF�ä�tV��E�\���SbDx�U{�ا���%�\�>�u�3蘎�`^36@N%U~qc��J/ά��V&���:%_�9s����vy��?/slg?n�>_�� c�t0��6�=�"��u�P�� ��+rH��_! .:��r������I�Ax��C�O��뵇>�}�<'7&v�O�j|d1��X�+�0��A��2���5�j]������fB*����;a��f9�؃�w��W�M���ï�K���DZ	�%�@͎`�־~�ݝ�N'���	��q+�E�PG�[�YvQdC���<�����|>��5��Ӂ�>� �����s9e�&���T�W�L\{��5�����\��o���.h^[cF93͒���"�.�mM�,;���i�8���
�#�B�h�֨��xO�B�`���m�,I]��WH�H�S�Y����;�}���ذ̿���;��Y����5	�^ɻ�����:�7.�"c�q�d�"�ﰟ��I|��V�!k ��w5`d�>�|G�BMq�!/�u�u�����JzK�4W�Aۺ�S����-�NļB� ���L�݂&���T�Հ�A�P���W���N���8B�B�m����j�p���M)	�$d�atS�BԮ;%�hHC
��Z�|��]��ך~�l+}�"�H�c6�#�DO���O	�����6�{qAr���t,�g��I����»�T��bnF��|k�[h蘿\��a�.%1:�q[��OE�C��ɿc�_�Ď�\���Q����GAR�B3���|���G��`%5� ܛ#�z��#	̚�<-9y_���W�|Xmd?IW���� }������?7.�	�6�
��H�ע$���J��Xf=ꇪ�mSt��o�����p�ݏvKE�@�}T��T ��{[�d�@�e������l_���U6fɆE�Q��U!�r,ǅ	��K#��#��4� �.QL�}@I�T�oj�]L�����;�H������y��'9A��ٲ����݇?�7������nV�k��:�k^�O� )5S�����[kAڶ���l-\��^���ք��Es-�4Z:���e�� $!:��)�~1�.k��>H�K$���
�dUWf�Ao.��������=��[��ݟ�o8���2($>h��ǉrq��7H��2�(���c�8�gf�쳛$^���i|�Ǹ����E�j+t$�=A�޽�:T�Y��TD��Knq�Ƿ�xӚ\S��X�?������l�D�^^����&�V���&d��杄@K�v� =���Q�Y ��n�[v��4��(�6�z����)��X:=�q��vs�I;:�H�u��V:���q�Nd뭈!#d�f�;2f���j�6Jj�&ـB�m�E��)�UP��Qp�'��}�J�� ���{�t~&3#�0�mxY�=��K�m0J����J<3�[�dk�k��&��f�Fd�Sda�l��4��D����
��*�g9��4`�9�-kS�2#�=�B �-
�%f��~Zeb���CD��j]�?�@�	]ˉҌQguf(nuJ� p�$��3QD
0	��4u�d/C�a����}Ĝ��	ٞ��ϰN�#>��Ę���a)�h�u]9R�N\��_�)I�%�0� �����Q7�$�,c���:�Ħ�q�f�OɆt=��2�k�>�3���&���2Wt��Tmݥ��e� �`L\7x�qD��a���6�	;�d�tiNF۫75�ws� `'����ՅK|jY�<�Ǡ�Kt�`�D�z(�ާ��[�Wq�����LlL�*���n�(�@��nT����	!�%��=	�'Sq��BI�\_�n��I���{�5bz��F���#蔤�{4�F��'�nM+�H�ѿWZ�P��c�!��{~9�@�t(�צ�lfMT��o���&���g\� �9m^RÃ�ǿ_��(9�L���h˽ON.M��	����Wa������RM���6��������c��7�=h\��6)���U@Z�R)�j����u,����̪/"V;��}:"��Xa˗��[�WC����"]�?&�O�[R�؄_����;��&�F:�&�rd��Ḧ́��5Z�]>��ȐS��*©�^�u��9D;Y<W�}4l��)�(��c�0�_�H��S�;�Fi���S�T_: h`�ryl�#�����L_����lW����E��pdA�PL����mc2f��Q���VI���� qO_C6�s[rM��
�LF5�:�<b�9�ɚ�!�1��5��+7�;�w��J0���������Yd#4��R����)|n��w��R6JOS㉰\�x��-p_�eS|a�n�����S�B`H&��f�a���XT�x}�5I��d���:��M3D��+3�P���,��U���TFox�3*K�O!h�Az�*�x3�2T��_���<�t]�@�����4>�}�륒�GB_�C}G`�N�Sو��B�)t"���l�%��c�)�	��Չ(�>���X�_��<���K��b�=�l)zx��b�>��̬���YJ����l��sY�����ž�l�������˹��}
��&��<�����<��\�Lj)���et&�\���We%�$�1��/��H�(�w���ׁ*q�����'Ǩ�f�kmET	�/
V�}'��j[�k�4}��'_��"N8չ��`���U"��������w�\C����n���{� י�4p�(��]�r��ݤ5��%�9ag"lC�y�8]��������Oe\�IV3�W�YH�6�s%�0�?0��Iˌ�	��$F�;i�,���è�|�E$Y�팉J0d�O*p�D���mW�z��k��t!�3�o�><2���9#��-c�]��t����ܔ!�7���ߟwO���#\p���j�dX"�%��CM�#_c>�;R� w�K��Az���:�ӎ�}nYJH��Px�e���1�����W�q��z�#�;�+搲U��N܉"JR������.v�0+Ĵ�+� �#��0~Q�<��+>���t����Uך`��ɢr/�N�'*x�w�eۓC�qr	
ID�)%�"�S�)�gլ"I��]�f�Yy�!�\���A"Su�#"��7�T�g7�`�_���XV=,��?XMN!s��&��HA�U���p�+	!�ǟu��7�%ȭ��C��{��(��e�p�����Q�[�0c����j`�uF���!�Ŵ��z��fd�9��d�b�Kn�N�$4�ۛ�e����VY�M�yg'��q�,�m�\���FV����+��*�X�ρ�a���"j�,�6�F��Ib}3j���P<�3�e�nlX�,��=�� ���μ+T}e�ӡ�,���q��ы6�I�*� v��܍�#��qpNx��H��o�4�3�o*���{@��_ct�Y&V��g6�d�t�L���L��t5�v�zN�#SL/�����g
}�'l�,s��(������^<Zm�vp	fs'��b����3�ů��gǞϢ��Fآh{����yW�5'��g\4h����b�4�Wr���<�_w'���ylM�7�<����r���\է�(M���A.��n
�7=��y���2�0 ��$�X���(,��ͅ�k%��)�D��y��-;}\���ל���f���>x�,C>C"2�״A���i��e�i*�	h6Zj��?T���So�.4�,����$��귐J�"��H����Z�Z��_%�Z��$6��nHW䗆[�uU�:���o>�jeXa�9J����s ���0ت���/�y[�m��|�e0�V���3�J�m>	��$x�7엏�l�����D_r�NH�MQ�l0�r��5a����<��j�XBc,����ӊ�+ev�z,�86�"g�k*h~c�����q����E=����{��O�&��IE�]�D|Q�$�/�p�X��̛0h}�F/a���&�w.y3���07��v��ts�L�ؚ"E{�������o`�T.�����̪3�
�J\5!��%@z,��W�ExJM���x{���)���p�'|��C�n��!b���=���|eUw{v�2��{����8ǧojIBT�WBr
��Q4���c�xC>���1P�b��y��N����'�c����7�DVeSj�	0��??e<iOP���r��%�������n�24��d9r-{B"Z\�5����\q�Z����i.�5F��ȵ��o�, ��?��#���Z������~�:]�2ө��|��+3%a_��w����!���*W��������`�O�S�7��Y��u1��o5l��uyR�n
�c���"`��K-LA	|V�ʥ��:%�$��9��|"��>��t�jK2�W �[gz���$F�˄q=�>�j�8�f�?=7�� ���F���%ϸH�nt4��;bS�P~�.���xx����_�S���EA�[�&/���6���=��hl�۱��O�41��D�8ܩZ�<�
܉"[6J��-0r�@^��`y�D7�:_x��@ai��-�Q���B$RJu�[�z�	$
���Ƒp�D3�b���ws���%Xn&��g��u�M߷�N_~9�.e���g�����B{4�K�c���'K$��"��+�j�Txk
�ܢ��&�Ok/<��}y�fHcٖ:n7�>�Ӕ8J;�/*��P�,?�g-Wy����^��<��5*	����Mp���EZ_~ 3�s�Z�y�xp���^dI�T�F�;O?z6��R2^��8�?@�mhg��S
Y=RA�xILPf�q��YK�{����p{(B��zr�� �k�J� ,�Q���Wt��s�
'�\��4%cƠ�km�H�]w�- ��/�r>��q�� �"*YS��a��""0��d��+(�1��Rֿ�,��UQ낝���O,�ѩ��T-'ed����e���#x.)�8�ݗ���}���|y�T���	I\���=&ӹѫ�!�;�˱�$����	Ȝ��-�W�ך��b}��{`�rҞ�f�[�Ћi�0�Na	�7H��t���ߛ{�_I����
�-��$y��+�eb��x��,��PNu���^���0��{�gmA{'���'�?_$�������)t՛���%� ��+��
ˎ:[�hp��I�)�k�`�р������J�U+W l������R�j6����,p�����o�&�U���)T �ەT��kw�D?"��(��<�R��Dq?�}���P��S��CU=�@ȕ�A$;2�8��^��ǌ��]�+���s4�?r'1L�{I���q+k,G�>Z�����{Vt�1�Ɏ��K���Z��zе��(}��t�:�v�]��g��y|�{Q��i�~�{ke+j|z�2R��q�D�~n|��!�Ǵ�2�q�Z;\dp�֋��#��i�
#���0��CEY��#[�ތ��#;�N�w.���.����=�$�K�C�l+�6^�$f�]��=^#Ng(��0���������7$����n[ҡM���'p��;�R�\�.(�O�Y���P(�.=�dk�|eZըT��8w	�j�C�׺%E��E5��5�M7��7����X��H�-�5�	L�����_w�',h�;!D�`��G ���uc���S?���姑�Ӈ��"Dܯ���(�KH�1{�Ջw�K�.B;`N��Q䙛��ʽ�U��(��mY�V��C!Ա��"g=T`���2��4A�� k-����R,�����"���xBw��z�6g	�HWK��[�vְ�;�f�_�%��7�ʏ�0��SW��Z�\UQ�ȭ+h��Q�IL����.�|5���*y�3T�r[Ṕ1(Ρ�8�g�]�G��v��llq�.裶.�Y���	��~_p��R_�p�4@�TJT\Z_�O�a�4�8��7G	Zܓ��g������09B(-6����TiI�C�j>*��*�!3�'�������7�clu��H{d<#w �r���-%��)�wl<� �d��E:�n���7����̬hM\*��n�$\w(�����#0�a)�5u��<>EX��t�*b�&�&�6�Ol;�HJ;�xς8PLj�{�n�?O埂��ɛ6��}=�m�9p@�R_j���>2����KDs�m����y.A�a��g_�]���f���4�>}�~j��ԗ���i���&�{���x}����ս,�6B�����f�\��6E긬=`AT�.?�-�f�wl�g�|U��N.��:N��"@�$\vk�z�?:�R�洚>�[;��lh��Yj�W�a9�?����)�4CY�9�t_��u5�L{"��6�H;����PO��~bH�	_(q�_D\h!��&��NJ�8���G�ֱY���d�T~u�ޒiG�T(�ܚ��|}@l32ۨ��s+t?��w|�9�O��؏HϡaOZu�^��Xa��jV?�_���X���l<(�wͪ�I���}�W�[�'!�p��..Sf�l�@@�r�|@��:Y����wQF���d¥�x���TO��R�F)�b�VH��no��ˌ�""YF;	��d��x�j� �0SeF^	0㝌�ttR��h��9�܈Y�:��F,���3�,�Hi�/)���
4Ҳ)���4��r�GlĊ�jqc�xU�u�}/�D�z��A�F*��$[��n�~Ǎ���ը��$߯>.B���]V|쎀"��������6���.��{3�p�:#�v�*�.%2�c�-l�g$y>j�l{HC�[��؊�+���P��|}��41lc��vC6S�pPG�^���>x4e�(r��p�.�8\�W��#�DMuI}H����a�{ܻ��"go�m��ӭ}���,4��@����~��j�w)�<��A���������i��6!�Pa\��s�>3�;,���@�tY2�������q�	�!@��Vx���A�LWҁ1{�J|i�䂓U�('qџ��o\C��bL�c�3�PUr뾆;��[��*��N�!hx��IW���:�����2W��F�+���/�Y�$l����ȟֲ���'��6�C&br|��M�f�a��`��d���~h?�8��!�Cʩ�\��0�T�f����ݲ����]����L��A��cA/�����t�8D� ��SE���~�+=��m^>��.���;�}��M��LR��j0�;�6`uoha��IY3͑�L:j�3�
Z�	�"	-�������AնAk��C�;!�m����RO�$ni(�����&������K{ZCf}�@��� .n�>˹�_�9@�m��RT�W*�`���~���1��s���E���/$�
���!���%�Z�AZx�:��H��Z�	˱����}�
�m�g�1��eP�r�(�������E�������38��'���`D��M�sF��ӄcf�/������>����E1-@݋�s^Q.�H�2��NA�=3ʐ�[��c���yNqk�k��0n���(m��m�������9˫��R���mRj9�����/6�2�^�K��o�p�:`��<�7�x�w*�G޸��?K	R�nK��(x��Q��l7N�����Y���ԏT��Ɛ�����B���b�AC�;�o�o�;��.�I���q%dOh����H�+�G���v���U�-�tF��՘m7�C��Z:N��Y�ž ����yg�ǥ�ώ�֤#��sq�֘Wa倽�+=6�^m�8h�<�Y�l�xjatf[� \XB��5�{�(��_d]��S����
j�5xd.戰O�Sz8	,�����^<~�n!������q�lD��*���g�D����~d!�/��f�I@a62��LRR1#]�V\[�{��g���EW]��v�ӫ���k��[!pf�
J:v�(�h�^���ևƽ<�g=ۛ���B�`�9?M�g�s�:3?�M���J�x�U�j��㲑�O��ќ��� ��6 ��\0L��K������(1����xH5+C����v�oN9\dVCF��K܃]	�W������\�_� �lo{_��ۮ��'�,�˰&�W��GK̃u�)R��\�k����2fsqH��I	�p���_��̱EQx\�U���]PA�SWe����'XS˂d3+Z5��,$��$D(˵�������>���j��s�]+>��0Z?7Y�
�f[Mx�z�n<�ʷ�	B�2ު,��A�2g!E�������W0rB��Fw��TE���?��@��� r.'�o����_��7�3�U��x��k���6�i�3��C؁�vŠ��"�Z,";S�� F�/�-4;��� ш��@�{���'��RA�[��t�z~��-�g������u'���H�#: �V�����z��)�h���6�W+6�;�e�K����,��(x�1�����۲�2���V�))����R���x_�VT�(i�Fl!K��j����*s��<��T�5BM#L��2>�o5��'��ڔ����{;MW�̪6I��{R��H�F�C2nc�*�+��g0��њ��9zo`�	~T5E�D���Ɍ"ҳ�"7�ެë���6��7��˖�z�)W�]I��?�F?���g�%g̀�Ž}���)º��7>ƨ�,�)y7�90\s* ��2ӇUK�;�^p �l��o�@{��bӼg������I��ۨn�����< ��@���]�w�//������A�r�bt���"��G/
��;-�#֩6d�I��\��YŬ8�'��u/���^���Y}�lҗ��PW7�����O��g��ʨR�Sz��+��(�驣]5k��t�O�o��N������;� ,�全�O�VD);�d��i�ȑΊ�2�Q����l��� Z�9
α�g!�"����������ػ2�|Om��<8�FSN`,&!���?n�:D.��_�#�~��BV�2n��:[��;�)������Y��j�Y	�-<��1�o8����X����`7���H$g����>�Kqq�Jt�al��]^�Ċ���:@���8ȶ\��s!��!dĐ�o�)a��#�c]�bnȍn�_���d�/+wS��]������h�\�G�~{�a��{�Pokx������˫�}]`w]��f#֧B���l,Į������lيH��s���2$VWd�q�oy����'��R��Lv�Æ���O؀*}�C�`�K�*[�&�Q4�=ԟ+�`�u倩oKgF43��sU�K��s4WG���J%i<���	�y�#춮��iR�;�ݣ�	�e	A�}��B��/�/�d�H�#�o�s}D�S��%����k�ӿ������b�,dR=�+W��s[�gY-���i���K����p]�s���M�����
%�WB�5��<����� P�� ��8�?��
?/��r�ɒ�]�'��I� �6� ���	t�8��8��>HdC�ܣf���()qzh�ι�Ǯ�(Q��T:���Ɵ�D{�Q���0u��~�������ϫjw��o��1�6xW'���ww�|���+sʍӺ��[������N�S,�'q2Z�����X���'���l7p8�0�������O�����������l&\/��a�����	[�O�xD].�X[ ��.xQ@��lc�����!����8��Y�a��H��Ӳ]��,�I
6O��7�Җ�S��O�{r����D8δ�(h���5���#�6�K-L�je:R)ii,[��M�X�1X4��`v�n;�3d&���vP3'1�$�~I^����Ԟ-(�@Wkk.�T�`L��T��v+��ؾ���^Ɠ�NczG=N���M|���[be��	E�w~�/�`�]x�x��|�����M1/vޜ����#ߤJd�Xͳ��j�X#Ǵ��_�iw�8wc\���Dw�屲��'n����fb)�P�;���B�Z����y������M)�+�{ѷ���XQB��q	�:�Q�[ݜ��,���;���$�@�\Ъr�*�`��m̩�#6�d�1ڭA�����[3��;d`f�$"�����n��$+�f`������\�����-ٱ> n~(�͑���z�5����NR|�S���I�8�>?ϑ9n�γ���e�Ӌ��Flm�\t���w�pSۗ�m��B����т�M��M��ًn����9��d�#����כ:=Ctz���0཰oakе'Ԭ�y�����-![3��d"Y|�?��ny�p��*$�?��i��~|�c�y`B:�^��^ç�0�$�i�O�����PN�@M�T�)]�{.:Z_�+���^Xp�k�PO��m<P7��Z���U���>RiSk��qsff9��в=1�r0�]`����߯X��R�1�t���A�ܑ:9f�3W�nA�å�����>Q���D����e�9�:#�@���C��at(.�Pm���%P�#�x-�M+�>��7?I!�0�SbC���,�Z�px���č��i�s�Y�0�nv�xB���5�����t��ӫ}ڟ^+��̟��7 ����H߄@-���uå��
��4�$���I��T�����ûЏ	�����#q7�Z�,���$x0t5�����`���z�l0r�ڍ����E�������TQ�T�/Z7�Ҍ�)���*���b�_WFr��.�i�C���r� �eﮗ�Vp��7Ȧ�����P����Z�6V�,/���L�|� �h�1� ��9�s��c�c��^�i���D-{0���E��g#E	����N�޻96	Ƭ e�t���1�==�=M����? �ߚ��7-��r��429ޱ���̯�!�F(rt���UK)u+Q� yR�k��U��5+����Q�N��c���Kؗy�D-<�ݓ��.1���:�p�-�\d�D�L�]E|��B���ށihdk�f-�<��Y7c��h�`Au��'w4����H��W.�	O�&��P_lX�i��F�OY�9�y]�Ҿ$�-A��c�=aZ���	�i���h��l?��'�[�@M"�{)�ө���ؑM�+B�N3���Sx�UG`��F8��u�|Xj0���o�.ځ���Xaԉ�(g3n�d�LJ״/C����4#���ê	5�Ѳ�����k�|�vE ��}	 p8b>٭�}�Q�y�ԫ＄�Տ�N�Qk��p �������Or| u�A�H����e[`r�����k8�}����k[EJ���`f��L�z,_^�J�B��IW%N]��HQ(R�yW��-���e�*�HN �T�v4�z��a��s(�',���!�$�Lgci���8x��wy. �Z��]+:4�<��=7�	�	�=lG��Z������x��� ����0P>瑀O4~�Z�C���N�g= �,�D`�8��wB�;�E)G�By@���m;^��Ґ걨��7�,��~l�֭)�1�x�"��C?ϲM�M/L�^�bU*�ovp�&z\9ܡV�&Ы��{/��=j���;�У�fr��J�o	M���6��R���R2Z8��^��Iȋn�So(Nz$��I0aY���L�e=�����:��i��WNg�ָ��|�^s��yJ/WgR��W@"�h���k>��)l��U5����亟㒲�/F �@�E��L�.vl�J��4؍Aa�ۛ[�����yH!W�Н�`�T��z�]r��a�D�(?�q����Z��?
L}C��F�	ay���;S�n��1��4l��ߚ�À9Y�<�Z+�s�/�5�<0�Q�Kť	6�W����[=�����3u��@/
�JF����e��w��Խw��r��I�am�Ť���9�_�w�N,����U��=��r#_�<����U�����g���t���,��cͽTd�Tc(%qX�?��f!1vꌊM�$����6b�6���o�@��ѶX�I�Y�[�����g'-)'�����O��+貖���n�P�<.�����L��]{�eF|��A0��4�����=�ȵ�hz"��`���G쉵�E��ʀ
S)q&t��˕��Ɏ�֞~��X���c���i�u��^��;~X�t�F�]	�-����t?�8[�8��@���/0��Ԟ�o�5 ��c)�&W�i��