��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VYq����x�0Yi-�#/7��*!;��;y���b�kk]�ȋ�0��4,^�y�;(�|H�K�NZΫ	ՍY���g�:�Mٞ���J��0��ĭ}�2�bFD��ָ�C��1�1�-T�5��X�E�EM�3���͛���d�1��;)�K&�!x���0}Qw�G�l�
��\������u�u��m �pdC�E�z���l]��|j19{�%&w�FB/f���׷X��Y�
����^i��/�	7G�V������I[-�[���K���P:w��Fz�w���X��y�D���p��.x9ņ �<fć,2�;c&�h��Mi8ޢUx
��Mby5���oKz/��Jk��ǪrSOT%)嶐u�C�"��F�z�Z#����w4�(�(Bu%�L�
��������9���/Өc���q��6��u��U��{�3ת�d\3�nh��\�U�χ]"bM��W����`�c�[�t�����G��ͫ�{�.�c������<��>T�$��O��f�����݇�9��y�fD,�p��U�F�#̑�sQ�ru�1�Hf��������N�8�@�9B^9�������)��Spk�I��<�4��=*3^r�􇁳vn����(
��e|�I�h*a2�yԻ�B~syw~;�+��%mƴ6���Pjn��(I��tW��ۧ��^���dLƲZT �B��#	-lx�J�����9$����J�9�J�]��� ��|�*w�ω�0�p��3H����n���3ȭ�׈Q�PVu���L8�}ԧ~�T*���;A��M��(M{X�{@/�j�\g�˭t��>������bY�"m�� �v>���lFz�
�c6��a&r��á�G|5����A����[ܾ�wΘ-|0���ʓtw�Xtc"j ���0bQ�L�����L��r��nRsj`͖�g����>@s��ЃQmwc)����u�Q���FLIE�WX�؊�m
}!PCX�M��YOa~��F�/�	L]E�#���sjR\j�it2t��
��,��֧�d���/��7�3�Ȯ�ɇ�gf��ݻ�%�~I瓁���>�?$�rA�7��}��a�c��}�M�a�K�Xnq݇��U"�Ap#"@E]6+j�j����˺s��0����|m��x#4�E�ˉ5�i�b#��.|����)�Pр�p<s��H%4^��a���S�a��'���@n���y���r�Yz�WV����-<kau5�� �?�6���C_`�n�D�V���44�{w2��\	�⍣Q �@m�8�W�/;YA�AV�whP���pNS��Y�t���+�K��x��Y�[g�4�)f[��]�i���3�j@* �~.$v�	��lWN]�>�n���#�4h8�h_՘��1nl�C�����A�����y��*N:��Np�:iA���A`�_�`4��^��τ7��S�1p'y�!gS��t����p�D��ͳ��?~!�o`�\x��U�WwIp�jB�v�{�3Xʌ8!�4:Hި����`�z��8&ĒZ �`U!l%A.TqY؀��������;�R� �1��C�D��A��-�]�l�H��D/tW�JIE#s�i?��x��'7~���:�M�r���dڀ�,l�3��fɅ�Ҝ��%��[�V���JY7��q8���Ct��)�.���|0?�� ��)���F�u��&d"?i�?>�����|�Y�N1c��2��`ݧt�i1&E��������
�d�O�%�o�"��4���(���~m�72%�*
,F�������]�\ng&]�P��^�k��඀��7{w�Q����]QWq?Z] ���ѷ�Z��op��'�ٙ�Z���I�n'U{t���՜��v�}�B]�a��/���1^��bn5Чi��F�
��tf��&ѯ�fT���*� Km]v���a�������ț
��H����ּ��	�$��C�t�����<�*������"o����G8B�}ǽfZ��b���I&�+����� ��a�ڏ��ϸ-����,�˿I�@��j@����Y!7��w�t��5OLl�%tXێ��z�T�?��x�LE��?��`x���G�Z����xO��۫8���:���|�Gep���I�C/���ڹr Z:���P�N�E!�D�⥅�ܛgX+U"Y={F�|�5f�/T�ĵI2��+v]-|ח���͏�&�G	S�S��D�$�T|\g���M�}�����b��엢��q\���]���12i"�k�}"��*rB� ���d�!�!����2�~8�Dd�YF~Kb�j��I��]Q�t���"���6��W�ra����pe�P�*yH\ro�K���f6 A��oP�uȔ����i[���]���b9(�a�z�
L�3�ܛ4��H=��A�g�k׹��2玺�����r��k8O��d
|z~�қ'7�n�   �J'��$�����M4����#Nha�[�߫�^���4y�e���X;4�p_HA]nw�2:�ˍ��$�1���%a�&AS6qz��D=�5-!C>�e��WZ���������g����
�u�؝�c�/:�u�9�WYxC�?9m�d�A	#�&��2ه�#Q��u3=�����
�bA%�G�h/��	2�u���g�t��+��n����b}fO�řt����o���s�)��-Y�>~�|u
���GٵE�^���iL�#�/�/Lm������x�-�s�AN/z�w!G[�^���Z��QN�߱�D匋hM����pOaNU�b^�)�ֶ�d+��T��	��!_ˑ�{�޴�|��f��[������J�sq�^���Ӝ�Fp�T���8Y:�E����͛â>��O]�H`!�*�/C���z�R�k��������X'O\��ݗ��^]	h�����9�T���GSZu�^LZ^^������zB�M��#8ꭠ1��P9U)��4�9:h��KX*n[��{�1�̍��ɏ�h}%��f�)���d
��
�vٛfM�;'(p���Wφ�Uy>�S�d��������/�Qw�"���2�&r.b��r�w$�h�S͛L�k������DB��k����b���k¯h���n*6�'=دW�4aA����v�l���D!�a����7������I��n���v����$6f�g������"��')M�\��{��+ъ���J�?ʽ	ٸ�,jm��-ю�s����m�:�»Dy�gu	/@�$Q�)ˁ�ۙ|��J]�L�!�h��2�I���L�p;����]:���{��!Y����J$�;4C�߃����u�]Y\�Z�s��n�>_Bb.���=E�䭶�� i��3�����R�0�WJ�A}�}��Q۳6k��"j�Ax�@GG�@^tb'ݼ�����,�{�eg�Y�Q]#u�0~}bNo��5yn��>�+}��Ѭ.w�ܚv@cba�ɪ�=��L�B��_~��C�4�p�&�d�+Z-�w��\�^�t,H?�#��'�q�9���<�������=32���	��5[�<X��N�&}/��(��s�-&B�TɊ\�h���6�%��$�8D2�+
��.�24Qӿ�n��%�d��YBY��\��l��QQ�TN�bj�O�� a��ҳ]z!�MHJěy~P�j���m<�_�{�G'�%�n"������=n^Z���E�ݻ$uJL��N3�.��/����\�*P�I7�RC��I�Lj��6��_� u8�����%�ȝ�J�0���<{��/-��U���:RF��r��Q�O.:A�LA�J�4�8`#�?�i'����4�}z.��S���
��]����B���	8�H3G����)�y's�lT�'�М�]���ϼ��ͥ$�|��$��d��$;B�ټf^�m��M��M�jr y��\��IAOu���9?v�dˋ�V�iD�:d�"�74/0��+4���7����)���t�v�E}A!DX �y��X�0e�1MB^�:�wN�+5���u,��n�s�^,q��t�C�����Ȝ�ʿ~�9��,��B-"H��ֿL�0����f����{,��:ѥ��Q�.>oP��p�T*�RX o���zc��@=rb�����R��G4�𙵔�wc1W��oy`�4�Жئ]&>�F���M����S�F�{
�����