��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4d��oc���_LG����*k����۾�T>x�/>:��e�=�C5!)f���86�$����ԤE���oZ�&�x���� ]1����V'���Hci������I���-�;����{�g+z������b-�ݦ�e�Ow$�i�y�{/ʳ�q�c������޼������iqV�8���~�u#Q�3��hKu�Q�>���)����	B|=U�K +�������0�$3,��;g��o`�!�eb�3��Td���n��J1�:���W�0We�c��M�Ե����{ԐQ�JHR����@�����t�h?��|���� ��rEd�t�(�b�^�ވVh�tWq��y�ca���[��^�Al�t���k�qq�ةí'��Z=�;�$�Ly��r��هe��4�t�b�*Qҧ w��@�@��$��^;Գ�j6�Z����������8�7��b�lEr)K�qiD��{�ZԩC��I�0��O�[��z���e��fڏ�y&��y �����Xj�g������j�0L<pf�Q�"OB�kL�� WgA����\}�V���<,D�~',Nm�)���"!bK;��M:�"q옳;,�G[}��8W�F����FM�a�/����h*H�k��Qqpޢs2����� :5j���'qrC`���'��?��P���K�C&��n��Ϻ7ش�������RŪ�1��@:�B�Y:�Ə��8-���iu�ݝ
��S���?TE��.��Av�J2,n�fQ<��P*"S��r��K��O��_�Z� U���ԡ�^Y^�7��EyWG��պ��a �%g���5~���ʜ������1Bώ�Dx��~�P�؝����N�[%LF�w���W5�y(ѽB��ƺ�?Y�J��9�J��-�N$��Sr�\����8�r��6Ŝ��dz��ъa�s� �4^]A��~���{;�F�{r'�I[�Z��,���6RU .�iˬO'eB�QC�$�_�v�c��Z�Ƣ�?�O2�9.�@�["��U&74�B|�Zo@v�N_�\���S���$m���%i�=�F�[-.g�æ7O�P���T���&p7d������@��A#�/V��b�E�l���д�ԛ"�hoZ_��Ւ�Y��퉗 qLnu�y����?�G��w�C[\�.X)����}s��,�i�¼��dZI��3QR9��VTF�v�#syA���=g)�8d4a��5)I���F1�v���|S� � �&L�b��v����� �f��>^�X%�K���!��x�:�"��� �㩻e�f$Hd��*�A���7z�}1�^�������a �u��(|�kQ�=+���O
H��8�r��� �-��ߍ�M��62��%E�7�uL �q9���t&�r?�6�(�Zdڧ<�9���jХ��7���p��_g�Q�h$$����d�D�����Z���m�ӬA�S�I�/!��6���=s����X�j������gJ}�
|�u^�K!��y�R4�<�U�r��#�)�,�j�B��	8�G����޽{��C�96/e�v��
��ɞ��92�t�g�{Z�K�� �i�,1:����2��j�[��ieP"B����5Nq!�M���-�P��S��8h��_��$�/?:^ywhK���)��N:�
i�������
N�dП�{33��*�H1��l�H��O�L6WE�k=���}ש�e;�IHi���<�c,����f0L��u% i�`��Fݢ���ޓG�l����R_�K[��s{�t 9kT��Bn��g�JGb�HYs��ߟ�N�w��Wh!+2V��N/�?�j~���}�t��u�п�?P}�eΩ��_R�i�#���RR�j�O�b@���p�y^�qZ:'��A�(��|��rQӏ���>�%��4I�}�Q�ye�]uݓ{�S��H,k�������ge�,��V��RC�DC�����f�8S�l��y���ux��{J	�r�|}�D��s�����~��q����۔1mRȨ�Mx@���9����	���wY��	煃HY��Ͷ���(SI��*�����/��+-.t�F��� ��%��^'����6�ȈѶk.��qD��Ix����YK��������|)��LZ<�� j�M��.1�%�kf�[2�iC� {m���0p��VG���H<��>||� }Ɗ���zCa���.�B`Wg�
8v7�~>Q�\C�E��
����"k�w�������O��i���!�W��O�׌���؝߰��_0�h5'�*~�2�2r�����l�QF��S�Jtl*��;����n�K�׮�'O��(Z�l7<����r;�_k ��9�'+
AUE���^yB��Ñ8����$�r�Q&{��o��at>*:Z������3���g���K
Pz;Q�,���Y�y�k�����ʣ|�"-t�:
�[�)�DㄴX#(�P������MZo�N#���!b:���)�>C�E�<HJ'|\�ID�k�0�ڬ~�2�Y���_�޳�o7����rd�P�3DKo?z0:�E8��;�n��{=aޫұ�#��jS�����y��L�h��5�)���Wf,M\�W.��E�x$0� �%D��y�������L�(9�R�T@ 7�E�Y)�,���	��E#�B-���s�x�p����D�K�&�oi��0��[�%���+� ��"�E9=\���'����n�_��w�/��+���0@9���_��#�Mh�l�us�1�7�Q��tu��b 8�Ȳ3��]�����(���^��)I;����UbW�yi��
�}����S��=��*+� ����:�X�T��&�~̉�@Z�D��\89e�VgOT�FUH�t�������<\1f���}ߤ�!���%דIp�I�R3����0���[v怇DR�{F��'�L��G��V#��h�E�ɢ���������@�e�6w<�Eil~G9��Uy��%��50R�C�\����$C�G��%�
��QϬܯ�8TP��eT�'P �40�)�J�`�&j�haޱ��m岉֡˳H����Q�Rd$i�"�:�.�X
B"%�03�|%Q[N�P���4�n
̆�ľ*�eFq�#h-�۟�8��rl�U(R^�~s�Ҏ�Ti~�&�D(���'�=w t�� �'��I�n]ꅨ<7S��A]f]}U��<W�ˠj��B�ذ����L-$���'�~���\ʚ!��~��Ϫ[0 �Q�dvK���'���䢹3��Ր�CFy�J�.��Gr���\ lU����W�G\~m���HM�/��V/5�P���D�|� ex��A��"�Ji⴬��Yx�aQW�M�Fu��qe���:i�Y��{�V����_���&���83�X���+���Y��#������ܭ���´�\bf��7�YY�>��X����:�'W:�oXCL�9�:��Z�u˃��Dw�h�e�EA\�ba���g�Tp=w��%��w\ c��$��9�hϣ���\�Fls���<�Ka�O]lx������U��7�J�W�����G��rq����z1�P�7��m������e��l|1$>sO�~ĊI�P�������6�@�A�´��������FAb�,�[��O�4�S����62�XUfZ�(��^��.O�nv|�kNt�h+���jKBeg[���D��
���Ѕ��_�NJH	�f٩=`Ψ8*�Y��.��>��%R���B�=���l�ur2�8)f-��G��d=��w�ǳ+�W�����.�r�#/���.�@��G���rV��Vݶ��N2P��-$H�U���f���EAb멪l7v@�?D��������4���W�l�Md��H��@X��"@;�T��<��%�Q��8(�ԥͧ,�l�Y�6j�f+1��H݆�fa�V7#cw�>�(uQ�ņ�@{'%+�ݫ�@�߁�/Υ�G���̎��]��w<�'W�
Ê��L*4���%C�K=�h��J���=�/�r��ۨ��/�I�mnS���cP�+�Via.�;��Ƥ�ՙ����G��T�])2��Ց���|�?*,��V�`�|����S�Bc׋��1`b��&���P*�G�by����A�\�b����O�e]��Ey�fm.Lx��)���W����P`[�Â�Y�yf�w��J���P�S�C�Ϫ�T�C�|x��΢��M
��@���T[h�BH��P,�'��u/�ڥ�PL;�ҧä�Ț��k�;u�����ո��Tm�E}i�z뀼l����3"|9�N/� �FC��vh�N�Ƣ��ˍN�m������b�5e&�m{���'$5�� ����2\i2�B%w��3'� �#�Es<�yPZ�kW�s�oA�@D������a)u� _�7���i��i�"l���������*jΆdԔ��)�R�h�@%7GDP
3���$Ƿ}���Z�UX���>�R��a&A3�����Bݟ*�ԖM��;��%u��Zl�����G�(�d�U��Y쥳�~��3��r��-�l��f�j�pAA*� A��1j��6���Q����.G���:e�;h��x3bV����M� �`#�<gٌ�6Ĉ���:Q<E۷b�Ehip���;�*&N�M��A4�u��%r
]vIC~����(�uE�±����[��^g~��$:�%`jf>V |�kbIz��c�\zݍ�p�j]�w��>	B���[1���}F��MbM��Sbd�~�
p�9%M�k��)��x8�rA��6�$7���L�Ȟٷe�}>J�#�+�٥�|�I�mZS!��ׄX�R���Z#�[�m�'�.������lr�Z�-&=!���9��q�v0 �i����c�OZ�»G�6�P}|���1b�K�ZGu�K@h�x~�Bf�/[tܝF	�8��>���˂�(��j�4�@ ��E��F���3k��]'̣�AF�p���-ueo5n�������G��6� �k���t�(�y,7YN�a��֜���?���׈�2�7)-��?����w|�3�<����j\*���9P�<e��	�2��ڂ���X���,�� �J�x���ye�`���������G|<naH�lO����� O�j���ۭ 
��[����R螠�zL���`X2�z[N[<�������̌A�����*mS�/l�Uƚ�b<���s��j��2t��Y-���7�< n�̜e�%v P��D��<��R�����ڇ�g��?�>�-1�!��M ��8��%3QP����M�������2���+�r��i"B䂲�Ӫ�k���;���e>���2�s�=�_����KA�}tZ�(��c�1o�c+[�gg��^�[=����E���hn6�5˾u�4E����uߘ��6��>�9[�	�O���Q��z8�0H�h�B����7�"An!��[����'m��D�'��U*��N~��U�iE �1���?��HX�$mn��y��!�c��݋ :�/���'i[���S3���.�2�(����
����.�kz��d0�y�[����2;��~�F;��́��hKg*��)a�0���K_Ǵ�7�j9����hϡF��߰ν��@[�S� �iU����Iuf5n���uSʕ̙L��c�c�F6 �VR���1-�uB�D|Y��������
�f#�u{�����B9W���~�Y���1*�/2�
h0��&����AѼ��b���Sj��o�{҃�d`��1�YY�/����<}���\Y�Z�/�n��U�j_ũ�V)��%�)�9�N,5�ϟ�`?�8˳��7�ca��D�:��+�� ��E��0D���Q�[ ����Jpӏ���X��l\�i S>{B(:K�[��^����QK��ע���ܺp��C��ڗ�0��@�~���ʴS�Д�ٖ}���Pj�'��F!B!צ�M{=�2ى��S�yߠ)oY�e����]���q�f.7Ϡ��l*�:�8�(�u3���Ru���01E�|��	��UAz	Dʾ��.�I���%*�zy�������6�T�h�W�O{�e�uv!H�'IH��������h����GŶt4}ʁ�9�~���s�x�7A݃+(�_�F�csb��1T�!���DjA���1�}&�]�wؗ"�:[B1üW�fufz�X��&�,�O��Eaܔ��Ƀ,�2|]��_\a�4}�wV�>�����$>��gr�n���(y�AY���JDg#���OR���{�YZ�yw�p7UA��#i9�	7PņOh�!:��� f�`��Cv�@�6��L�c��Tp1߫�6�Ӂ�����Gƈ���U�F�LD�D���]�}�]A���Qҋi@v{��K�Ȱ�?4�ޏz�[�V&﷣���K���X�����g��	���$��]��Y*0)ذ���
�Xq^�������FXԘ��P0���>�W0c#���*�j�ƪ��^7O�x�
E\�➱�g�$�R�u�`K����\5�����G�Kqw�"�� �܄N��%�P�X�D�z �ﾥ�*m�B;���xhq�r���-J� ���i�&n�2�c�\zk@\����{*T�SL��_�K�W��b:e�:�y^�T5�)S5�a����Ъ�� 7	�(���0>����j����Ҫ>~-��D��t��y�S�gk�G�Z����;f����`�)�/n�f2�?�s�3Y�;ns$����vqC��NZ��Al�\6'�]���\D��4��d����� ��J��4ڃ�d��0x���C�$k�����n77�Mё������vPQP*�� Wc=�@H3T�/W�!-��:O�8�-�>I�@bpaza)H���ChH��݇ۊ���y��i�j���Jo�W�?'��\�VM����� `h&9W��4o��M�(sI��is��2'���c#�3f���t!���ԅ�.�_��ѽl+��'۔���3Q�@D����j詁���-3B��z6).��}{��M���%��O������c�)�����}˕�_��9y��/Ʀrq��"���q���6�O�.�Ȧf�^�׳��0gEw<Lf��Mf����[O��Ơ/7�lŠi���MR�B���f��j)�d�7���9�����Jыw���1�Z8�OQ.#p�����݆h5������w� l������?I����&�����jah�^f�[U{z�H�>�:$(�1ɣs���A^�p�!��[��h���bΚ5�C�����g��;sJ��̆�ӱ���%��u�6������(ձ0{��)U�+�)���p����<:@~�z�{e-ӅU��>�l$�ƺ�6�Ew�,3��U��SJix8��\�A��@�.����W#
I��s1�ˑ���quMY�ǥ>�j�)���Ζ� ��{)wC���%�i���6��DDZ���dLzr���庺����H����#U|y�;�1��w?�ߤ�4}K�e��p:ܙw6�HE�]'�X��g��!�C�,�T�s�R��\b��5�pO#I ,˧,�g��*�KJ����s]v�,���T��&h��~��~�s�{�fc��<��j2#��_%�_��CU��V0�Ow3\�Q�&˱�{-m�urVk���a�/��X��\�v/X��Y;�N�����	��
e� ;��[5�"�;H0-��~��5��]�H�Y�"� �x&�|���]���	���,��`?��q1�]�ş�O%H�o�[�,�����5'��eI�%ɓINk��f��4��,l��qWK��R��>9�	£��!d�W&�N��,���򯽜S�I��ns��nܓE��n��|^5}0p��v������~�D�vz�o���:��n���Ef�Y���+�͹ݮ��蚡fW$U� @���٫�D;]PO}D��#Rx2¯���x�K�.%pޞ�{�h#aT9pr$��E��-����pEM����0)[n��u����`��κ%cI�Z��0#;9�_ Wc%+�Йܠġ+�:ؔXv�q�ޡ8�nifz�����B�9��$�ٺp$�o��l�o��& WzW�&M��u����}��_�p���Ւ��)\���#���0��q�����(�^�Oa�wV��� �F�ϼs��MC�Ec�m@�����K�h߫O�E�Un{n��b�MN�
I�u=耧��C;��x��Gn��'�\�%O�5���