��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|8���e5�I��d8<��1h��}���:z��n�Z@�8B�:+%��Hx<2r�����OuT�m{�I@Yr��RB���*(�!����:|�wB(�{>�3h��nR�܍.�V���_1
iP(?(&êI���y/+S�u�b}���?W����X�\�d66d�xE��V�1�4��������q�X�}K`��х'�p��D,m' I'�F��Ҍu�[�9��ￛ>��h��n
W��5t�6	׾��pI�(�g�O�-���Uq@O�-��Z��)�~��>d���e��".f��b�Nm'
�	.f�%����4�17��"��;�Q�t
��Pyp(���~�$^�m��&��Q���3mW|�w����s/+\��湳�WH&P���+p�?����p5][gd����u�f$�:�K�R���������ښ�2�4M� h��B�I5���|��D�!�����3�zq�G;,j~��\Х���5��R��>v� �d>�/��l�Z
-�s> k #^��A�J�<�//a�+a�Sk��D���6g��,f��ט�(C7��ۮ�k�PU���Ԭ6J 8(*n���pė'���8Y�;VF��e��^�GR��W�مo	w����7V����%��8 \NO���LqVR�_A�Q��w ��M�<be뮞l:[WS�|��_d�Յ�o��?z��B�鱫G�\�u�ޛ���m�����"�I2�@��H�]�� �~�����	�(�e{�?VOb9�~+�.����t�W�u���8n1tBs�G�t�#�e�j��
	�Wn��!��FL�8����	�t��׻�*�i9��F,@�ֺ����u� ỵA(e���Հ�#���S�~xٓ��u#U�ЍIl�¡@H+.ss���*��^z�a4;C�x�24��H��JlE�u�۫ˬ����)�̗�֭��7����ׯAJx�"��6����t����r�c<���E��{��M`tra;�1�|л�F];����5U<��ڨ��p�'wv�d��)�*��`%�W��\2�hG��F��\��%�vk���T6/�Z��T��ȋ�Hov]_��&�.z�.]ݔ�jLO����A�3��q4�jw8�eƨ�ir��۰�{�~Dǻ��ٔ��D��Oyl� �H�LZ(J!Z���v��'��w��;�nZ�Y��K.�ìm(}�����ï�����"	|H%�T�-;��f�W�	=��䀳���2�:�L�8����u��MDP2��?�.���1�>���� ���EJ��g:�?��1B7U��U4��XϓI#�r/�6~OSp�S��$v��$TR0�ax���iV��GB��X+wаBi��$�L��m��]3��6(�M}�:�����Le�[l��mLs��zL��@�]�� ��|xݞL��g]�SO,{��S�}����j7S���ep^	U���p�y�I`�5����ۊ�nи�����v���a]P�v�]ɓ)�|!V�j�y�s�n�^6H���V˻
���Q�sXc�|�ι��Se�;6���q�������b3���vF�L��vX򽏵����?����f�h��X��e�fr`�����.\ґ���&���|٤.J!�����G�\vx����_��.�h�2I��&
�Q�����d��w�o�}#<��uЖ�_�f5��m�b9��0��n���E��(��J���g�=JrpɜVΑW�\�=='��6�5�$����>6mju��[+L���D{E�t�J��W�22��!~'����JȽ�ql�����3�x����{�ޙeI��w�^��`������ ���!�4�;�}}���kj<Sg��G]�UPu�#�����F,
}K �c���Ib��M��l�f֮��Q��n����>X4r6���SI�ր\�Di�BF2*�qir �W��R�������.�l`_]2ԛ�n�[+���6
F����B�ߑƙ�[.�%_Δ��\������q�>���A������'bL<�A�T�g���w���a#m�8Өu�v�;�����;�?,G��:������Ґu���J�o�R	��}����ϐ��o��n�S�:��@�Ϫ��c�#c��^��+�?g�?��Tew��'T�����j�!erٖ��ƜUZ~�<$�]�j?��'�ʷ�|]ZƜ���o�a�d�yp&�z=8�F�Cuk� �վ��5DQa���*9- ��9��z=7���G�an���(Y+��Ef]��ȫv�ק�M1����S�}�z;N��:��s��U�l�`jD�t�o��Ug��E�;�C̵*�_��4ѧ�p~A���8)L�!Zi����J#�-�QQ�y�v��8���v�L�0d慙%&Ay�;M�"��"pQ��-�L<n��2�]������_�?t�)a�b�;�A��6B+������8g^qjP����38�>*�_�����&[X\l���&�C�����¿^*�z�3*3����\�Fb�ʍ�z���g�4�(ԋ���<L�-N�R?��m1m�O��eĀV����h���%m��S���G�2��k�}��/x��7�%&�������8c� {�Ԅ2������Q�Vӷ��q��3��q�}��� ��A��m�n�P����`�M���^88��[ xl�؝�.ĩ��/�����&��"�=�<�Z��҈����d�l�7�y�9��[������+�X�Z:�(�De?��/TE�����*Iv������i�c��E4kz��fS�n���l�|^��`���l~��C�#�@�n�]�;K�� Rvz:Eu��b^�%nx�XP�i%%�f������wKi�Zli&rLb����}f��2����m�T�e���ջ����Я����ִh��%�3"m�j�k�	��^��?=�m~�,�5��M��Tl�a��� ���-����AT�Iͯ�c8~qp&m�}��ؿ0/���̢}�$G�w���amQ=�R%��^����,�������y���9���)K������n��>$'�k��PqC����tN9���̶a#��T-��ӝR�uf��*�8n%b�	�	�▶%�&p�����~�O��!�X����U�WQO�J;��'8�
�e-H��YF��r���*�`�D��븫0+���Q�tP]k�����7(�M�Іi�
Z�jBa�kC`p܅!����WĔ������`��6�:r�rz%�	�*LG��\�����c�	_��M��Ⱦ�g��V����C �e5t��-y0W�y|�Gtq�<�M\���p�
��FI��X�ؙL/��,�(?��+3�������2T~
ڡ ~R�6�?c��?��J������5�����&�mu�qen�Rg(���Squ�Y�<�����'�q��Y���nΌ���ܸ��d���E�Ұ���!-c�"�IM���ު��+%y��)C7k�4�|�z��xN����]I���V�� 0ư�ZY��O�G>��`��l<��{�\��E{1����@���7�FKx�@��_\,ƀ7�V�P�^EXT{�x��x)-�א,~�+B��k���F־�d������#���sE׳ �G�}��JKb�L�)z��W381�bם�r�P�VT�2-�t�l
v����Ψ���dY��f��+��7�`,�2�p=,:#\2����Ϊ����R�xI�R�*�T��̳�����UŤ�~wD�|Ӥj�i!c�ߚ�έuʞ9�Щl=h��i1N�-�X��3c6	�s�HX���l����t�N�z�a�&�5
��$�xB�6���+!�0�|��U.[�S����y�p}��T���{bRi<MU�(JU�e��EЪZQZr�,��
>�.97��6qb��5G.��q%p���v,TZSf��"�P+�E!��ɎD���ج�k�[;}��C-�W0�=[&�Rh�+��4������Dݯ	�/,�B-�D�,�i̘ly8�@�An!8k�N�m�ϒ�a>*��<i���'HX<��Ty�L��wȥltu�f�S�h��6D$�Up��VrVb8���ơ�)�?q���p�+<�����>+��-�p������⅟��^~w|����D#\���lms�9�����V�~Q,�(B�����!�Ŋ���ˊ��r���b�M�J�h����̀~�� H���y3�`��&�+.;�4m���ٻ%l^y ��0LH�Yq���j�+��*�F��|� ��Ci09X͆��{9�d�	�M	nwɡ(�x@�
)`�<͗�%�r�Z-!�AKԋ:�BgEw�$<Xq2�������[�i�:���9*��K�$H-ք���<���5�4`�H�%Fp�6�[�my�R�Hf��{�a�1Uٯ��0��J�U�O٦a=���>�2Q�r��� ,�N���mra4��D�c��`��V�n����v�e���W6��\k���ҷ�����ӽ������|�0�b5��ݟT��ExN��0������y��=->�F(#��>�kl,MK˙Z�A�����=�T̤�0ۋ���������l�g(0o�͐�v/�l����꠾�zr�$�z���R;��.q�zŽC���Ȓ6j�����"OF�9Ѕ���7���o�$��,L�o���/N�J�$n��E�U2Bɦ�I�Z�ޔ�=*� ��]bqը&ogݙEg��]���6���<�%����0|~���۪�����������U�d��� ��儼�Dą���.+��{�.��
�G����
�u_sӗ՞��y`�$�����rj���ž�̻�`�� �C֥ T�7����.t|X���A�&C��s�� <���7ђ�1Br�T����٤�e.,���G���5�R�^���>|����-�l@U>�Ih��xU�a��K��*�m��qR/���%�%dXu{�	M���}�K� ՗��B�=[�y���k7�L���E���$���Y8�G��ٽ���E�!d�Ͷ�,�Ta凤V��1���o�=���]#�T��q�3�?�Y�:���D&X��'z��q`t���mt�)�**lռ񰾀�G9u��eO�Tn��D�2�����&�LHi�ژ���*�M���D�i�6j���S�c��p���{-SoE���A��a	1��Z(�R=n��0dH��l����T�SFNc�EMץ@��n����[%���x��7��
l}̍���O�D+̾�\�6��9i��%���$YօN"u�k�1/$���E��!d"�n����(3�H��~)Td��}�_�ge� �4S��J`��B��^�(�㔌�+ܕ.������/��\��.�I��ػ����r�*Co����FR!ך�D�Fϑ({`�R�<��<�i�-���J�F���yU��i*#
=>�u�1�͗u ��T���K�.&m*#K�ٳ%��q��j�pi�R�7(�p$C4��Y��	.V����/@t��#�Y(��Q��B�b����g�>ŷ��������vlY>����٢�",��>�[��0@�@6ʤ�3�[ɑ-{���b���9����ۍz`��<y�F1
����#��kh$8���+��=Q�������]g0@\s4U�}�/	盿6.:�	���B�Ք;����d�S��kem��&1�J���N�۝9�.}��Ҽ.��2(yȃ��V�/���M����Ź|J��օ�׸i��룭Dp�Bq�\Q�Q@�6#�1�'H�~a?ލ�����M��A�,�p�j��I?������l�&eO`�Bu��~�m�����r���~����N�!Qd�惇���u��r:��%]���S�:j�'�)�sB9�p��}��GDf��y�nLm�$&��r�ce�X=b�_'�0�J���c|9U�ڏE��'u������Ps(F?���3�⟶A > σ�G�</����<͒7'E�o	a_9�O{ފ���GH_	k�
��r�����/�/��⡱� 8�i�g����S��%^E��J)�*�O|S瞙�3ɺ�=�1q�8�@NcxJ��F1�Mh���,<�Q��we�
�b>g��v�?�:���e�\[�(��JM��. �K���}K{�Z��O[�tߒ�lI����������OQ͊��Y��,�R�nÅ���F;�#�p�7�ւ�:�4T�r�}M����+
�Mo�  ꂄv�n��0�d�ˣ&6L-gt�gU�3��0�]n�<���bi�l_��pZ�4lb�Oh6hMc�^h�{��}�Z�$K!i�t��|;���6���Y���"��;[��GO#}O��Z.���`<r�z�J��|���G�Rp��-�R�Tk�5��v*~�[+�<�d�;�Ω�4��	��Z怬�\�-����� O,�W,x�q�٦�:^Nr?=�?7�o����y7mA��Y�ox��h�E�����PX��p����5!-�V��V��D&�g��am�ܥ���z({��e�&�N49ǃ��E��~�8�d�[|ʋJ�9L�f��[S�)Yk`v��,�{8ׁ�xM���g�-���g��z�d���Q���L��%�����Ý�'�����"��y����<,��Y�
ֈl�_6;c�5C�L�i���-O�1)[~[��6W�Z�����4�tS�k`U�g��1����qs�P �U������z��k��CT��e���X�����fՄѼ��dWzX���%���;�����0���vlDP1�nw��Yp ���\���@$^�3�YS�]��kk�V'�~��RC0_{�bg�BН��"�r��Zl���% ����_� @\<_,��1*o�&��Ua�W�����gA�\O���oJ��#bA!cn1�Tu��,��N�Zs�<풟��k�d'���Ӽ~$i&U��'|l�n����@�-�0�:R���A	rk��]�y
�`i;�dF��cv����:_]R�z�
.&��	V��8w�N[S'����I #O(+8��`�'�@��F���+����~�0�t�ϘG4I�i8W�N�ޘ��d>�ӊ]9a�^�M��M��):��,���-ydpb�6ƨ�~�>�$̹���K�%�R��,I�hJ|����������N`����M�����M2���zs%��	���&����>�����[��gT3<j��X�9H�V�.�P�2zlхi�L�i������i{�0p"[ZrP����΁/�/��e�0���s��ǐE������?�yq�a�\cb~�5R�q�G��+�����CT~��t�=���4O�N(�f��s�d�� �%��͓0&֬�>	|�xz�(�&@=�.�$7�\��u��5c8k�O�o;i�-1��d��[g���z�Υ���_cu���T���yf�5�J��S�m�9B:��D4k �L�q���k�Oj�S>J�}3m;����~��ZI��e<�C�Et&�="�¢X���c�K���L��lHҾ���P�!9׉{��ac�Uq5���,��Ǫ���"��jn�I�ppv.�!yΆG��[���"���o�g/�hck7.adU?_p=Dൃ�����T����R���/�yƑd�b�cIұ��'Ԟ,d����$;p2Z�NP�����~�Lu2�~�t�x2��ތ/P'��)�ࢌ{��M���&pD��0�`��!~,q<Fn��|��ٿ�1cW�0�Ż�k5!�C]Evn�t�q�#!6EbX��,�r��t��Q8���YǗVH��8}	��XbK3�
�,�K����̸
��֙�M�����_}�K`����̓	%�n>�6G'OE3ځ��Z�nn��mY����*ޠ��������r{����):_���y̔k2Jt�����5���muE�1�!m����gӌ����I=�)��Ѐ�oW��nn���h�</?�~�I��PR�/V"v3to��Q.n2%#"����ax0O ��*��Բ%�>=�'���R��vuɅO�NƛK��!Ӵ�&�#��9�����9�4'e�e�iu�DH0�������
t]�z��a�d��A���$�5(��l� ݐm�@v-;�]��X����'g��]���Av���Bhb�N.@�l����B����r��ak.h�$1;X�K���N	�垲-ja/����{Z�긕�AB�
}ߒ��2ĝ�Uz!{�<&.��O��d��P� +3�f�t�xjiP\���VW���4�{Ŏ������0�g�8���bbb6�v�$AÝ�zgJ��Ý���z #��C܉)F�ٙ�w�)E߄%�Ѫ� $_"ft��_7�Q���d9��H����]�.�kW@����a8��+U�X?&�������p#���^$�w���C��M�zE��m�Fz\�Ӆy#���z�$�n&c�F���VϨabҳ�
DG�T~\�M�XN'M#|����(���혫��N�\`���>kއ�AE�D� �-R�lټ�t��Ԓ;J���sl�rP?h�I�j!~��v�-R��`������fRl�*��q-Ҍ)�����]���g�������e�+Wl�/eb�B/����1b����,{/�S�=͞:���C���\�	�s��c�!<I��Lf@gQ����[�F9#�XWT�^zM��v��ߘ����O6|���K�]Rf�t,B��?�gx4u�.4��ߢ5���M��&��p��0�C���������<����7?;�!���)A�����=R��Wi���ǩ�;.��^�`�-���	����LPW��=�)n��L�ͅBC�$��9�'=je"q`3n��x�#��=�@��p W_N��SGh�"�|?enE����ڀ�:�i=��s(��>!�O��i��Z-��U?�ԯ��A����ߎ�cc�aTNE ����{����o��_�O�B{s��.��_���L�~z3�[*�c���kʔ�����^�oм��~,9h~]���t��	�_��2�I�aB������_I�cUx�C������r��3,�k��h�A֤L�"�*�7D��f�+�(��Ӟ׹JMްP�t�@*�kX�,��ǹ��NNMR{��<���/ل��"Z�u�u[#�;����9����r�QY�W�3 ���%�ܥ��XA�~!�W5dA��|���qݱ�HS-��o��B���$���_��zW��ܱDO s{��Q1[��%B@7��Ga�v�����<����n�s�uCz����n)�]�rm�c�����r��/7B?�6{�$
�D��qe@A�����<+>�G��~SOH��m�D~,����%D��Z�Μw��6�-=�h�F~�l�E@�HX��$+p�AZ�#��Ms�m/��**n�ͬm)SãD	�mp�G�Z�!��Q��@P���;���4�6�bI�2��a�*��C� �G�p昧��Խ�q1OWȴ6۰�����Ԕ[I
�i�u\��p+�vW��^���B�\ޚ�e|��L"iO y��9��&��"�����"u_fl�=4R�V�|*�;�����7�y�Xp��^�-q~H�m�*f.��sGsP��t����t�Z�D�m�r�]��~N��6��_�s���w2f��%f���s`��_���D�$e�$μ��7M� A+�(uNj�`���ȫB^�.�B�;e6�\-���#05�X��!m�c����u!�������٠n��7{��\�ϑ�Q��$��1-�!c����m��9�6�',h���[�Iw�D����r��䚗(V4���!5J`�wH���#���/�P\���P�
�Q?:�Qei$
��	��&����r�i�����T��~�	u�x+��%9����<ċ<���ĕ*���m�#�ÈW_yr->��;4ff��k�iE4�A�jn_kv>�~�x���m�,K5b+�A&��0���	���	\�����6}� +<W��-�K�M	�P!G%�W���<)^��ib�j��ğ8[���Wƕ�V��-/٧U�_�1���>:s��f�=�{b���ED6��7��g�z��v`,�!&�,ֶ%��2[���Ÿ}_|l����OɈ�vQ^�>45�XB�����:��b}�k�`N�0Vk!��-�I������OԚ�	�{�Q�ޘWn>^�̎�����~��ʬ�.�/��}|��D�J�d6�(�g&n�뭨Mxr�&�R�����ekQSn�?�E�O�_
T[$��W�����\@m���R7w^R+pn7���%�2�t�`��B���w3�N�ҮZ�-���)�l��n�"�N�Qp�]'�A�Y-����9����o��6dX�X�
�޹&�[YH2��Q̟,��GM�y$3�a�Ԩ[)\j�!>��>�h�PS����nbb\��(�5�J�İG�%�Y��������A����)(>%G����%�M�}9� ?�ɯb����l�T��e�eJr�|B�O1o�b�����j�?{��9Ks�mzM������=��Y�(@[��Ŵ���g����.k;�+(���j\Qe��*�Y�X����Dl��Ý�w����&�eӲc+p/;X4aݓ��Ȅ����Js�OMtajF���2v��|v����O�-j�K��ꕶ��7ϘЮE�&��9ϡ�S�<=�󎋍bm���b̅��c3�<�f����=��C�c$g:�@�Q=0�Z�}��RR�mK��.k�tZj+�x)ރRM#�Z�QȪ�3x)�����t�1�g���jx��"15 _$����Cz�����m�T�� �� �9ޢ�X!����r���ZX�ކ����9ł�z��"UDK�m�3���-���Xм��{s/��;Do\>T\iM��i���w�<�<(�����T���@���f�����4rz w�`$e�1=���P4t��f�0�'�:�ntcS��Z���rՋ�u=S�@rΎ����^ާ��3��A�7�*�Y]2ku1T /�ҝ&!���~" %FZ��k�����v�l��&`��S���C��ص�]��3$KX��hƟ(g6y6K��N��.?QS�4[ǽ0��7�>g9W]�\�ج�E�Z|�k���h��]��y("�gH(ɓz�a�
8aς��X6u(�_$�ò���8E���+^̤������<���LE�Nx;;"�^_�jP�T��ٯɬ�-E'5��I��C��/h��jI��3�o�ms���I
�C� ����Wuk8h��9�)>�E��������g�~	 ��S�븝�uo3��I���^�87wLݧ�ݝl�'�	�g���C~+�#Z��P�ɧ{��qp#��?<��_Ox��jF�Z��Ex#����WZ�Y��7��Ɨ�'�2^A�{.E�C���xXW��LJst���&Iz|������Q!�.z��5��Z7�l�j�|���Ʃ]�.��2���*�ٲ�Η/s�L=s��Ԃ��*�w0�^�L���<Ho��'��Ni����s������"܋�_v�"^�)����4CJ"TĚrU�&.�j�'�}5*�X�:<i�Q����݈.1�$v)�4�|T�3z��S>��O�����,dK>k�H�g����9ǰH���;����\�d˫�L��:�_�-���Nmm��������G���A�vȨ�s�����ԥ���n���ia���7�5`;��� �{�f�OiS�}��^N�����W~#�(�b�ۭU���gߏ%�lO5�&�A���}���L�
S��)�隆�^��ό�k"|IM�H�fT㧌�i�p�kײܮ����Zq�\t �0�<�j~���daRT*:��Xc�Ȅ NFWYuKmȁ�#u��l�f�,�K��D$w��JFb��I��w���؋T���6,�� ~]��b����7�8(��>קL�j��p��xa��낯w��U����gkTF61,�&�(H��mΤ@	�t$����X�ǃ#a����'+L9�Έ��p)���VFE:�A"�b[DAԅ�@`e��4��wUH��y���'j�P�M�OƗx�`Y�Ӏ�V��Ƶ�����ډ�J�vU����Ϋ��Q���F�Rn
"�6N��L�:�>dQ�ɹo��������	#�����˾��[en�d�,�����ށh�k��$�8�����ncDʼwj���Ңߤ��G��@.��7��5ɝ���S>^LV���&����;H�SEԃtƐ���)^4�܊Ӟ^,�9�I�VΤF�HZ��s7Ja��M�;'�(*��q�ӹÃI�j�n�'�$hRG��[���SxVEkx���H���HV�U��PJ�HU�k���~�7q{���5N!^Zz;�B'�I���uH�Vb�/=%t�S��VC-n�Q�[���� �3���`�j&pO�G�[&F�kf8�y�X�ol��.���rEVX�y7���[''�f�D��ˏ�,�Д��7`M�����:\VF����6����%̷n����/*L�]�p`�.�� ���@����O@"�����P�%��c�QE)6�-�����ƶ�=�)��9�~X��V����{�:����ȓQ�d��H҄���G��I0�w��ț��>� H'�ji!�3��O�����N��~�)v����5�<�IW�?�7�I�N�`�~��X��e'��vLsn�Ӳ���!�ǻl7y��p��lE�]q)C��~�O��>N��`<�ʀ]��{x��,}>!E�����d�a��&��P�߿�sBS��ؒf�-��@��e��|K����/�`)!]�g�&,�u��A=Nf ���y� -��q�2�Uq�eU@��2Ȟk+���dc��_5���@0M���\����]18�K B庨Q�t3��=.`f��)v3�hMCS�Vؔ���2����"��Պ:�ٝ�yK?�V�qtOUea����b��]�<��6�R����s�bF���s]��~��5p:�`5+�ǰ6�����Pt#@��t��+��*�'�@�ѥ4�U���	�.'�?��t�u�g�K��x�#���,Od|�&��>����k~��"C�A�_(qNZ����=�y��o��>#��-ouԌ����/�$�q��^{$�3�3��o�A^�EZ�����գ��A]d�P& ��Q�t��:�
C3�c{C��܍qltNN��0����,�!˂��-;O'�#~żdd�/e����p�htE�jA
PZܓX��Į��hVY��rK4�k��
��ڜ�*��p8�'��`x;��.����2�p�'
�'�x�+,ˇX(��L))���������Xߍ.U�*����'*����a��F?D�tһ�!Vw��A��{E~*Ly��!bQ�O�0��NL8�����?ռX��y��t��j��$�M��7E�S�6Qr�|�?L�N�_P=ET�$d�ڐ�py�*3Â���e��b�>/��*zɨM�z�'�Q$��_�`X��ǈ����2�W��Y��Gɢ8��T弚�����L�,$Ս��
���y�̌�L���3{�]�n�tQ�ޒ_̷	��9�z��%�a O��ۗ/T<�h� ���.�Zv���6g��t�������F��J�-��KXx5��j���� �M�o$��fW}8�A_zkr���c) �CVy	�'��d$7!�{`zLV�U� b�^*��J��b%ޚM�m��Һ�J�G�BU��̷����ӱH�4�� �`��!���d�&�>����������F���h���VԊ�-��;��>_V�K��&GE ������l	S�øLǳ`�u�O��%C�]�k��y=|?N;��������x��|�+�mx��"�5S
�����a]�E�PK�e��J�觵�8e�(w�D���	Yo�78�t{c��x/�ؠNr+�l�&���=!���b��!�7�?rBvu=Z��pX���ͥ�ޯ�U��Z/j�eg� (u^o��1����� �Z�y��L�nC�w�1\ H��MH��
��l�f���2��1����̒�=�[L��g�H�Sp�j���sg�E��3j��r�p�fWE�o��!���	GKQ,�Q��_+�0a&���&�`���ر���L\N�`@�u����h#�w�>o���j�B�ׅ��0�8Lq���(<��'(��˫H�0�|+���j:��Lz��,ݻ!ষ���������V�9N�`dE��(�3~�\ۜ쐈����i����j�߸��F��F���<mc�`Cg�_э�3����`�t/M�tƛA�N�S�3;��ȕC�5�]�c��6# �t"�dC����H�]&�����w�FF\���5,y#"�.�l�h������c܇�L�]U�K����ԡ,ى����7������Qq�w��ܲy���s�(���Jv���^*��`le�M3�,�����/!�!Cfs��#�ǥn%��6E�׈��<��WC�K�Й ��Q^�a���	Tbki��G���� ��`7���z����O���.(�pg�B}<3�t�r��@�a���<~g2�U,1+���,��i�@� ���M���lz\^66( �`qM�V�X���b@%)du��K�y�c���6��KF^/ւ6��u��C�MC3��uf�[�F1h�䧮�^��+)�6$�:]O�.r��`�	�D��=�ʰ˺�p�%��&Jr�/��yS*6�j��L���[����ܕ��-�|͓Ȃ��l��dd7��a�Y�����K|>w�{���ט� Wưs8��s���!�!<U%R�8�H(�W{l���qie`���pW�W�O:C�����~�(̈́d�����P!+d,U�����Pv����b�4Kv8W�W��Kh�����w�m� ��,0�jD�X�>������j8�Q�<+�g��3�f�zEY8�E�}ߋ٪u��%o�>���qX�F��Ǽ��=�f�i	��&����H�RH��	�ѯ��hS!��[��X%\�ֆ��쳛�����/�UB.����XVAdS�a��	�� �Vgg�+����7 �A�!=%{�
2Lr�n�T�O�c��⪣��Z�x�#��
�jE(~�Ɛٚi�E_b%�`�&r٫���x�1|i@a\��	����-�E�r��a�@����� �N`y~��ǲ�mK& �B�w��nxq������(ķ��
Qm�e����t؋k���_�O�,G4e��yKԉo�;G\�<�̏Z(�4��L׌����*��Ĺ��Ht���\�Z�F@��\�^}�-w�2Hv��&��O~�/�x�s0c��s�K>�?J�����g�K��4�X��3���+�V�Y|~V��F�
�Ĳcr�	ؓѪ�C�|����KKu1 r��|�K�g k�ώ���0�+�(������ibL�&ڜF��0F(~��K�v@�J^��k��'�V+U��:��IMIW�ٵ|'uA�:id��俈�a��ŋ�|�D��ކa��v~(�č��uC<e7\���F�X�D�A�E��c;�?Ȝ�u���Q5������wV�I͛s�Ej"S}D��j-�7������J��B�9ˮ�5R����g�s�]@"������l��B��O:Uk2Nn^\*��\�ӂG�p��EN ���̿�?�O��C��MdP�W*} }M��9���*��	��0�t�α5�YԈj�º�k͝v[�;�bqL���LJ�#����`�8$�%�S�G��4,ϋ>�dK���1d��^���{�vqݳϣ�/4�-����i���(IQ�g���c_B�?J��>Ky�V*����<K��La�v��{<j(U���d���RGf���P4{W���Z�������}]�29�)xc�:�,�z���n���DA�Z(�L[p�"0�ܒ؎\��ujǇ����Y��ܠ���;h8V�}m0 ��&�4������ͤn�b*G��H��j��pf��ҦӶъ$�Аi�]�Ж{�����'؅�]�je�9�og:~��z���'9�	�c��Ȯ�݈8���L�Z�e��#��ųPa�r�t�.A|łk�؝�*B��F)v]�5�Ґ,�������Zr�X���Ч9O�l#��ʊ�zL	Ƥr�n#��H�����򊘮�1��3eT�SÆ���T�_�9N���2�@�2 coHhܤQ�JI�hG��K_o�c8��s8�?�5r��878!��z	�;�ؖYA��X[���$k��������-�Pw?�lK
v�E���J Pv=��i~ķ}c����+��	�^�Oċ��۔�~�V�O  ���$ob6�Kx��'���;j�~��I�U�ޔ1@��\a��Ɣ]��O�<�kuhU�&���Nu�b%=�	�UC����M��f����ϲ�e����٭:��k|[!_Ⱥ�XR9w/�;�h+�Ҍ���M`���{Q8e�Vu	+���"Ϳw�Ɇ�AQ;-�ќb������p�z��}�lW��'=u���Gfo�m(%Q.Ü9w��W��!����Q޾��ܧ�R�����?��G0���HOg1�Ӻ�;�m��
O��1㦰%۾,(���!0�OCR{(#x0�("����MRE�&��V�гw�@Sdq>���O��n�����8��(@���V�fGK�H�����]�CR�~�: b�>���^�$��8�T�O#C�V�$�h҉u����̹�pn�}�IҤ"઄ٻ�ZC��k�2���Α�]���;�v�n�u��@!��?Й�q�����A;��r
���i�Gx)J��vK-(����R l��5�C�ե���m��qBS��[GD�4[��7ʩ�`�:�9]�${͘��-y x�Hc�����7�pX���	VZ���6@qw�B�!��f�`Q���a�v�d�	����E����J�t>����aropD�#�/�,{���0�5*0�c={�,����rz�@�y8R�v���^.״��b�����J�D�o�k:'�l���JF�S��S�+�����<t<\�=�
����T��%�iD-;�h�e�{��	I� U����Ak,YyUؠM�K���դ��)F."D\F���]�,od}	��s������X���ݍc�^[��^9xd�
��GU�v�C��-#:�V�����p3�c|~�<BE���Z�[f����:���q��*�w��m�`��L��L@�>G��:B��~(%�Z����d�w�e��R(S��������Xv����Hn��s90j���r�>A��f��q+�'���&����[�
��(�X2��	(%��A2T��^�}��ؾI�6-	��q/�1G>i����p����oNq6���L�i��]M-����������_a]n�|$��RX|�'�A�4'��8�4�#���q��&��و%S�,�B(7,:��&W�OY��3+��ZH�&��9��/����t�R�T�v�|�#1r����C�(���^��IE#�^���p�!
�Û��n{\��LD�U�6�������׆��I��X2��J��1H���{�,�?��|h�X���F�S��T�>1�����������H�`�~Ŷ��O��/���=1��`�Q#�L�?�>	p�PUqR�6�m�3ذL���p�|�K��TfRz�*Q����1}b�_�6�-���\8���ZLk(|I��
�$��󱒔��9)hh�BK��e2;i-+C+����G��;{�*iXJ����Y��
���k�J��������qGTAc+]()���0���h��{��b�@���'H)�1}����2?�0�f��1J�|�t:ȿ~i�8�]I��="����G#�ǹ�焚T��B�hL�6[����аU;q̻��������2e3|}U��l�Ke�(`�
��d'���I��b��ļ�,4��b�(#�M��(0c��+'7�gEA����jҐ����^�,݇�f�B���u�O�i�	 so�[��U޸�/�L�H2(��Wܨ��Sw[���^�|a�7����k�Ɖ�`�l��z!�K&)J���/H�ʳ��v7��{~/8ȭ�F�i�6h@�c�$S�*�E[x��w�uBV{��C��pNZ�t.e0�P��r=��SFi���]p��Z���a�A�fu�Gq�)	�cy\����>A�N�a�t�(�+��{��3^M�����93@��{)P%1M�B5�L2�9|�MI
�jW^z��������K�3��&Ƶ���ش���r�r�8��M����n�J��Z�#}�2�Q��D�����S�N����>�4İ��J��Ѷ��_T�i��#|=i �;���4���sR�*S�6�fV9�E�$Iy�9�D�A`)��� |9^�\䅭 o������K�ݣ��W�Vq�B��&%e��߰�5�&��K��n(_cl��� @���z�_7��� �͋ �#H�3HA)!���hB���;�|�Dyr�<�����ʑi42l�j�8���n�u�'�++�y)g2}d��zi��0�.޿���	�ʙ����"�j�P;�Ë�tX"�8`�z�g*��zY���3 0R���D�o��̪��M�,�	v����!���Z�8Q�p���r��+A)�������ϋ���13��p�|�� Ln�{D���D���1��V�4�1��V��4z�g� _7X����G46OO"��D��M�*���/��&�?���;|)��S����sW��~�`~sAQ'�; ���L4^:R�HX��*��H�>�}��)��������.�9��vߓ���wY?C�w�5.�먻�ɀ�|�j�M�,~|,�Һ���7VaC݅;����m�*$P�s�(��Q"xMѰ��i	����=��~����'~����ZYP�ϿwO��(�O&	A��|��n(/��oRS�XK�^u6o����[���Ïv3}5	$Y���xy���F�� Wbܔ89����ݚॕ�t:Xwp�6n.��`H���&�\� ���]��b��(�!l���[�S�rݛrr!w�M��9�}Y@�{S�Mp�����]�P��`{k�p�v_%�+���3}�="X�
�Q��&���B��/��2�!���Z���?G�(+J\	�b�����a��[�jW�ֶCJ!�$�{@D��2!�&�x+`��E��`M�s����|Q�q?lھx �B�0-^�ŷ#l���53�Ĭ�C�|8��6Y��Xo|�p6Ks���_������n�TJ�ڞ�>@���ˇiV,��@P�n�0�R�m���W�M���[$n(�-�0��t��4�[T���J�ړ8 .�h8:Ps��T:W* ���L����`����f�1"Hr������q���Qb�p� �t�����m�� y�T��K抟�C�)������E�Pzt�P@8e��Ī�tㄊ ���bA�+�CX�)��Q��\�G�'2�p�^Xh�=η�Y��_(��T����6���ٛ��2��~J��lబn����Lڑ ���5ǧs����0�8��.�,2�ZU��C�O����P�g T}^�e���K��3����1��{C.h��T
��?��0ғVJࢂ�%""�v9�S����G*�$X���j!{���Tv"9RC��]����7*�I"
t��I��4.V-I���A_�Ҋ'�m�TK���'ξ�8�$4�й��^�sD�z֯K�N �x���V4�<��şO��XJe���.1��Ku��@��(�C
H13ǠD���K����a@j�߼�]�5�4�yq��M��(�[�))�.|j�m��B� �:-���yk����z��Eyv�l��m�;CĎ��w��*��=���3 >p�K6���X��t�55���W�^�b�e�(x=�,�9'�5�L�Jחp�`;2?=Ϊ������3��(�e��H�V�fO�+�ڔUl��-w�b4S#졂� =;_���Ld��?�_&�;(�4�T�_�Ӑ�Q|�q+�}�退4L#���?��$'׍@3��hO�b�F�Q�L�%��v�o��2��8��2�k�\�>(����#V�̒�Hꏡ������c۷�3p8�Z��#�q�y����G�7t�x�A���k���D Ie�c�GŰ����X�O,T6N�E��j�(�E5�y��=���fF��Ӧ��
 E͚��3mpZ� E�X��f0n_���O���3GH�E�a��cQy/�!pu��ؗ��x:Wʑg�=�@��d�l��5㦅lW�z8r�y�1�p�{�z~C@�$����⨚��x�����>���iE8�ė$��e��n@��&��=@�%�)����z�T㝣�-:����:����σ_|��6�M�������9��*ջfZ߾3]���F6��\�; �Ւ=����gj�c} ���6h� �p)���¿K��qw�ʕ�.�u*�"|�~�����đ~#P�۱yp�"� �c���Z�4��z �<�#u\�]NY�PBP������ac僈��bM�A��j��ZF�a�v=<E|��ܘg4�Xhn�X�d�S��$��/�H��Ɛ�4�%��)Sl�roQ��6�K�+�x��+��zaH�6,K0l��j�����_����-�dp:xؾS�Ð��-���{����a1��RGw~�֍�3"�p -�o��>���!mҲ���u1g{EP�c��fK���\DM\� ��ܧ M�}?Ը�U����>~>A@&������Np����m�[�^6(E/`)LL���w�M�q=�l�%'R����~�U	�4!��:Uṕ����5سޣ���S����Y?۽l&�ki:�ύ�g^�Tk)�a�����ja�(��Òp�c���� ��������p��ֽQ9�ά	O?��XS�(7Dp�3k����"%S4ƧW ��E*pc��k��?����]�?����e�\�V ��ͤ;�����*�d� �ٿo?e�1\�h�����~�TAH�%��<����u�i#�"����~��0�8Vސ��T7�_�2ڞv3L�T�	xE��$ؕ��	i��mˀ~;��J��9�S��K�#._grI���m�Zm��R� Ϝ*7i<��zt�䢿��Q��+e^���Ưܹ��`�X�pu'Sd��asTDN�+#���f��f	��mzMfa���C��0.�{κ�%�g�ܐ���v{p��eE6EV#u_1��V�*@�������Y￣�>	��^7[�:&P�y�$s���A���8A��3�0���M8�Q��Z��%]F&�<E�ɓ��]�*@;��)���[ג�ұnث�G��6$rb�뺙���+����'�SՔ��;T+�=�|���y?�#$Y���e٬u��zI���s�����!���S&�q	�/�������6��U&���-�}L����
��u5n�7íˮ���f��Vt�0�{��[XO�;0�,�sVi��w��(>�)v���*�2�����mݮ�Cx�|"��A~z�ad�Eњ�]�v�eH�`h�M�y=��{%A��y��)P8��w�{[�M%�U�-D�v�w �е���f?���L1�P����l�:_G��ki|!���k?Ɖ+�Li��9s�b�R��j\�%L>(�c6���̖R�ʫ�� [q"�5�8#�b����=dev]�2�܏`�3�W=��d���(��6>"����"ҒLiGE ��/;�g��l�U�?K�=R�ʦ2����hq�=�������w����s`H܎�L���U�-�`�� M��۱t��뷄M�_�6=�m@hՎ	Ĕ��N� �E�M8¶�?`F~�dY� 4=!gė@��Y���-��C�\�+��Z��*}ŀd�x����n��2�VW�
�� �h+2�u3`vD�B;��Q��E�*�v����a���,��l���]� �D������y�.��H0�0������4��0���mG&#�h� G��M��xR-Q�&�fy�B�����ƥ�Ź��*)*��1�1.���*ƶ�vx)�����JV�����x�� ��J8q/��H��|9���(��T�%w��2���AW�Vҝ��v����&����P �+�"U���In[�Z"qn2�e�7���|꺃 XD�(��!�Hs���&¥��#�@�1��C��)�%�̀Ʀ��y�Cꏫ�����g�����yIL�g��/���i�ڼo����+�5�@��G�2��GX���=RW��0P碲�S�iF�A�&qS=��Շ4��u"�~�{'�ɾϿ=�4e�ؑ��4�P�D�]p2/0�4o�y�g�����uG5	59��Q���=,�b,T�.Ց�i'�^��q��	FC��f�5)�.�����;)�\����&!v�|��=�'7���wߟ[�y����Q̠ �k�h�<�ss�V�ڭ���'˭�Ç`DYp�l{xT���M ;��]�I�����rKͽ�0�����Tk�≃��*ΐ.J��("�1I0=���(�cI3�~�v�7�F[z̜{lG�y`�(���9F��t~����\N;�J�ꥎ�]r����v����)��$H�2�;|f\���Hg_����a��y�������fM<�w��C���Ǧ��dc�j'dV���C6�����[��'*oE�U���4f$aa�;|SW��H���w�I�[B>&��TD� |�	�?8�"PzN�ýo��j�2�z�s�cpRV�^ͦ�7�	�D���t��Ȕs�HSLG�����伓Fy���s��Jnp���c��A��؀/׳�,N��[p,t�R�v!hK�*����p�l�����������a���K�a~�#��u��)P(�Z�**Ҡb�n$@w9j	�����{�Ҷ�:���~f�O�-�8��G��p-V�I�w?�uaqNxF�WbE)��d�N����nl=���j�D:�5,�wϧy�`Z~�_��
ܫ�V'q�Q�I�07�%,�U.�Z��]�D�Zo4p%݃G?�,���E���x����o�*P����1u�w�Ѡ�oޠ����#�$��4�HvG��cs���|gϠΚn�gs��,�.g��؀4���9��S��ʵCg���R�:ϭ�.�UŘ�������dqb�z|��uBP-b�z��7A��h1S�m�ٺ�i�;vK(�jq ��;�a��ə�Z%����H�/��)�R���o�u�Μhf.��=��x��u�L��rV$��� �Ю��5vX������]ϫ�]vV�U\�-�I)��!��x�pp�W��<7���
A8朞,��̊
D�_:��\z&�|�6��!�Y�(c�.�~�C��� �JO���COGS�~I�߽�PAT2�J�����?�'6�����S�U��J�-Fc��,�����<����5\��x$l)�0р�}Q_C��O��SI_�n��o�9�wg�zV���y6m޴P-�&k�����ذ�|��8�w���,]���YKu>[����[x��*�l6mc�l1��6��hA�:ϒ����ܞs̜m���I����y���D!�����=��	0zO���@7� "%a�ƶ�|��8���$h���[��32b�!�9��oR"���jV(�6��d��܅�Sb9��DH�P�߿U��|��B���\����?#�媍���{��D��K��_�ijQK�k��"�OЉt1��O�q l%b���X�ih�|�T1����p��x�����ŕJ���Cn�Rt��
I���9�M%�~��Z�'�?簧��%vpn�^�I6�+�:וi?��%�{�Q��
��z(�r<;��O�CO>�w��\j3#'6-��y*V�(Ӧ�sX}n�<k�1�N�����ex�qxJ��!aڜ�Gz�g��)�6��
r&������m�s7�ˁ���F	F�m��KsV诒Wu��R���2�J��)����q���K�VX-�6�⎕ �lh������ڲ�����ZG��m'�8ƺ��e�o�u�U��WE熢o���6euT�/7��|�8��C����ӖȜq��$%�C����V?�)���X��QNG�
 �=��Y����c�'Ӱ�ԍ���Lx7jT�,���-vL�
��T}0v�ҽ�|ak>���A'�83�D�f�H��ҝц@�p��(��RuۦJ���pNPPv�ʒ�m�q��0b]=��~_�*�"᧎�Tf���P���S7�+�ɏ��rN"+��43h��x�D�>Yʁ���'�B���:\����p���5�Rz�I�[q8*��$�X��=<,�N%D��iy��������E������7O�T�m�N��+���|ɨt����,u�mt��5�XiS�7�~���C��8�/4վ���R5'y���"ir�@��`�C���a�=��*��:,�������&�0UQ�џ����N��\�"y�奛g�?1�J��t#�9*J[SJ�1��F��ף����[+�[���e&���@�q=�UYJd�
r���.����I���A
r~�����ki�}=�
%O�z�o!�8k�x�צ1�d3?QJ%��*`ݙ�xrX7��z��Ab�Ʋ���v�:)�m$	�7�ɗ	W�LG��"�O��x0a�g�<8J�_�\/JU1F9 -R�����m_��$��9R�'2m5��IZ�'���M�h�*���ɉ)��o�O�{R�($$����F�t�F$�p���P�}����,j�_	���m<za	�t����= �#9��GN��k�ю�?��q��ˏG��|?���z
j9F�EY��FN�\J�BwȿR1���"�{�ca�g�ٿ��7T|8�z�D*��Ɖ7;{T���\�e���b!f(�S��h�Mv	�:$��j���?`-c�0 �� I���.$O��/L(ѻ�M����/9�U������
B���p(Y ¢D�/�AZ�PWx��XJDK���?"5�9DS�Uq���$��v0��SQ�jЁ%@��h��gM	�T?���Ɯ5��uY�X�T�uk�iY����\_���#��.|:�����N{F�3�iY�1�N�p�ą�ꪨ���Ի���hL��3ԣ��{ʕ
����&$�b��kQ��OoO��YV�M*���-�C z�[\��������@���?!o����'X�ۋjq͋f(��>e����	�������E�C�d6z�M6ȃ������1|Q���2��~I�̾�G���w�lq |�[R
;�]_g����Ty^�;�j5���J��i�A׼M~���/�kAvlFA���19�"᜗*u7w��gF늣�ښçb��,��\*���%��O������jYٌ,�ӊ�z�|�����@����c	�I�N��F�KA(,*��`�5���w�1n������'���@�wJ�թ�'KC>�Hg4�����Qw��U�pL~b{"K��_o�9D���D�q�w�"n��7�
I�����6�Pe
SJ7K?��=��zȧM�ZvC/I�JPГSbv�N��Yx>�Ŏ��C�a�蔯����o��+4�K�X���!w?��u�.�ȁ�� .>���?�3*�o&�� M�����`P�}<�TX�c���ᩙt�{��E���2��6�V�)�;�"/Е�5��NK&�7�<Wv�mO����d�=wqo��:��i�-���H�'!tM�&�6��v1�d��l�Y��er*�����B�v�3��v��h��t���&MU����'�S��/�j���]+C%\���>�d��x+�$8��Ht-�;��ǋN����,�Kߦ"��f��:� �v��
[�+l5c���Q8�E_V���9��+�;@Hx_�ԇ[7(�[ e��R&,]����B�Q7�i�B2��(`�����a9��/(�צ���G��K��`�w>�흿?�k
vE��?��7]�����͘�_5)��J�$ʝ~��9N�SnU�ܥ���@�`#e�̚���u���@ԁ��e��G�t--�ll�u�&~�Q�G���ڵ)�~t_�/V�W5�;�#3��Xa6C\�r'vaЭG���/Ա�Ә��X�E9l}pWLߗ�����rY3��Ϊ�
G�PCq�C����Ī�\�A�ן.i���߾G����s,u��|�ʸ���vؐp]"Ak\� ?L�����o�{�T�������il��Zk|8ϖ`�����⥎ ��O�ڔJ���J�|&�-����i���*U�C����J�7���	������:��1�t Yp1|�R}��O�a4	`�"����2Q��cǦ���մ����7�����^4������n����?}�<��pR�,�9{��z����1R��e��,�yN-F^^���(�d�g���:��^]�U�vB����8#�M7���L&F�) ;�x���vc��k��W7�	��D����|:�->���*��hrd����I&a�%xs]#��j=���]K�r��������Y$�m]����i!