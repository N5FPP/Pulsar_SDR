��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��e�ik3�������w$����g|��J^]،�[Hވp�`g��=o����}v�t�ב�$�Zy
"�WZ�At<&Ie��?��Ǚx u����Ú>�n���h����y��k^~��Χ���8��@�r�^��U)1�&x*�N��<��0fD�-��c3t�5C����`䃄�M8�R9r5v���D�H	$yS9��C{��dxG�SX�6x'�9RA�:!&�o�L���� 8�Y儼�����h�{��Q�����J�kD��6��U���� ����Z��us��!��:ѭ`%��u�ah�PfE(oе����;ѥ�=<�p��>HK|��5�����-Pm|�s�)Et��b�p-�
 ^v։���_(���i���O�����Uv%^�ln��i�{�Ƶf�!�d�E�}`c�:�� ��z�K\��x!���x�N�@&�ѩ��0�Mk�k��Ŝ��˩��k���0.��Dl�"�R>�{�Ӷ�"� Ҹ�¸c��׈ނxC�j�IE�u���S҉���i`B5�l�z�c߃�������r���x����em/�����kb�T�v�t����q�Y�i��_��x�J�������͹Z�]>�1�Q��0)�c�	�7Q�Ym�<�hX�ĺ�You�V�ΫQݧ=b	�y��e1b�߽}�����Sڜ�x���ZSi=]3���L�\�z97a?�`S}䧑 e�;����U~cK�`�+v����I9�ݥ��i��{�vS��$識H�����Su�#­�jf]������;��!5� bo����}�MV��f��/O�5eU��眀���kCz�j)[���;b��5����k�P��o����V�9���"��75Ci��"&#3��G��bd��r��}�'��*���P�U\��HF�Y�$X�"9�_�(r���%�m;ҘH���&2�9k�J���b.�a�2�����#&OrGú�V2ɝV?/b�8�:�x�\8E�_�y3��:�A�θ�M͈rz$�dK��q�`�nM<�kqSؾ?t��$qh^��5�q\�a�p���j��9>�u�oz�̖��f��?�u6��򨙙m��f�G_�
,����Y�/�j�Rƪ�}�?W{�	�ш�v�z����R���غ�e��O�v��I�"���Ŷ���e����ݶ�L�{��O�YV���,6��?gۤMD]�ݦs��2�4�ʝn����0Ӵ�N��ҥ�k&%.j4f^e�} ��:'c���$w����su;�4c�7.Ā�_�%)�!X��͉���K�%�$�JN
�N(�{�kF�ǚ{|��$y%ȕ�5��I �lQA���M���"S��
����Z����$"�h���_�6˸[Q��W<v~T�޻u~IOC�����w���G�Д&z<�s�����M����&+�����4�ZE����$M��k�g��6�<� ��S �g*���~�X�Bh|_�:*4�5�ƸۯN�J�\��X�����t��2z������.�gu�n�h?�Z"�j�ϟ�ڳq%�	o8h��L%__4� ����=�<��� 91i;Zt��1i�Ih��)@3w*�:�R�p� �IPq���nV���S��� F5�Ҝ���L�?��B�{���(+����f��������P���HK���[@;H���(�K؍�8t���:4�^�E�v(�U�®쑪���}�T7Z�dD��ϼ��m�Z��@̪�ud%�.pa]��*V��S��b1�Yj�DZ�� ��!#V���Φ�ސq��yNs����E�z�f?Ñd@���`�q�����S�忎���Y��
A .��fld?ٞ5;GAr�a�q�ep.cU��~j/ʪ&��f�k���u�:u�f2�ӭV��ݴ(.\0���eY���x��:���LvM�,���	��`��A%�����t��[Η�8�j�I�e�
��. �I�E��4�؊e72{�u;���Q߲n���h�J�V��IKF�+�}5�ENW\���ufm��~;2��L��-R�{o���"�����lD,����O0mo �ܤm���$9fp�wA�P6Bc�?o`�����ѝ��2&NN&Sj;���3�@�́���*l��[۾rϥE�`�噆�c�{4�+�5����A��;n�к'���VҐ>P����Ld�8^3�:�v*��>���XCX�:�#�IRhBg��~��<n��V�l'��UR-r�����8��������f<���3i�!�J�r�� ���K�}�9.�ڀ�c���`�] -�R� w�����zf��r~o��+�(���:�v��	Cp���6�h_����#�=�g������6�g��<�����W ��:��G���Ҋ0�N]�Ї�u�$ә�d����ݑ�~/���|'�-�P�1餭M-�H;�x>�����`�W�4=V��X��ҌMįl%h�R o^�d�@��-I`��;g�H���%=�#;����#m���C�JA����(	F#�قf|��Fꛝ���$?�P|%���fzʥ��1vP]����I,���}�,g_���=>Ym�.��+�G�zM#�f��S�[��p����[��I�|=ɊO��}�&��o�ˀa�z𴸳��Q���{����6[��\�z� �$u}^��%�X�bZ��Cz�U��c����� �'@+���U:�T�n."R�f����D�J���g��`5ͧު�gU�d�Vi尐�T�����L�&m��p2��M��mM_}*���Z�7+b�P�������秂�V�߇�0�`@����
! 	=Q^�DpV �2����!�vR��wIkZ�ڹ���� ŀ^�Y�o�d1oY�a��mL�m2����G��R�g)�M��-�?��a�:b��gx�s�r�\:�1c���<<��ĝ���zo�T��.� �Zȣ����,�b=���9��a�wqd{u.A��N��+�j������ Z�'�Ǘ����zݙM�2�#��|9�I�]|�U0�����D.H'p�i���k��6p���T}�ҍ�K���g#crO��X޾8����Ⱦ?��.=�# "^)F��|�����N�P��l���6������^��z�YD&H9+���H(��T�Y7�h�/%�C��CE���8�c=�S�?��r��qq��H:(ڗ�O&/��$�p|g�nBiF�>�g�!
%��Y֨/�N�4z�v��UD�QYp�9g��ٿ����f�y-a�|��I��7��ㄺvvݐY���	Z��,�p�������c��ni؍m.%^A�a#%@����^�4Q�����7��z���w��@~��0�i�l�e ��-���T҂������+��3XW�c��,�'�_��Kp.�}��rGĊmxi��d!� q���c�V`1�Ac�w���l�*��F�7��`ep*E��1#fc̉0�+�f8�����;�Y���@�'e�P�925T�b��D(�#'2B-��ZT��
$nG���'U :P:��<�%�I��g��6{5B8�W�=K�d��f"��K��(�q
2�|a�ܓa^���e^�@�%@��D	��1g�^����6 Vl*�p�>�)?�^ �{�Z����<t:[�*��(!�Ϛ��1�z��#b��h�-�MABu5u���>vf�H���]?8�Ko�Sq�+�!ee� ����C��``���u<����`2�	`h�����6l��I!'����^8�f�K�ͦi(>��$�TFh�j${��t��B�jH�v,��"�O	��d	p`��Ll �(�I�]��;^j7:�${�� DeK0~���H}I�k�T��qq��[��SD)駛���b�=����婹��ɋ�d�ܶ�`��ZR���(YH����eA�R�xx���ʽ�h���l� _�^"��Jˋ�`<�ZF��o+]-<(ݘ#U��BOl,<4y�~VL[�IA
i� %�� �X�씈�Ò��$�lA-
 �bwtc�W8��'�Z�qۛ�o������ѵ�Aǡ� ��݄�G1	����o�H��A�ne�1
/]�Za�/��g�s����(�0#�ꓑ-�iW�&�@e��#QO�H���gwMn�%�:^�_b������cQd����� �ސ�*�l�ԶC-�F��	����~Կ���w��/QAF$5�UyKZfw��V�_�-����KDb��PƾCO�[��G{t��z}�V@�mu��"�mIq� ���`��s[�#C�骇�M���Cޔ$R�|�j�}��3a���d�4^{FA2�1�>��?��Gh�c��T���}�of$bEx"�,O��C�BK�ыc��*~3d�Ld�^��$��A>�l�Y����e����e�z�s�U�?�kF�ˢ�VJZ����U�Med^���i'��� �J�at�
�����j{T�J�rb$5I|�zu�͠�s�uE�)�Bǀ!��\��2{f!:趌2*P=ƅ��OR��|/��`C���L�CpP�wA�!?ϊ��kT��t�o�w��d��r"�i�bP>��y'�GW�B�ۛI/9�Ɛ6=�ʑFڒ.��(@��wH�<-9RN� q�c���`������z`T�>�����ݲ�!(S�"���Bg�pÌ�βC�x�va2ڒa�:¯����x>��v����(h�M2ޱbKQ�h�](2>���ؔ��Ã�sK�S��O��7��y~�t�6X���'d� ���rơX���;��B3ۗ�F��3F>ޥ��=M!�e�X�><.�T��ӟ��H�6T�-p�d��$��)T'�%�3��ZL) o��:�N��M��o�?"�f{�!�k0��2J�\���e70�[*�tt@�֡Orfx/����\~v5���A1�ȨǁڬAK�*��fݠ�B��ȭ2;��N���d��dY�n>�E�{��2�t�q�pm��l�1�[G���@��͈�i������Xh���Ju{6
���Cn�GM(�6��Ǵ��-�hx�*W �F�wp#V3�I���7� I�0N(ި��V5�ϐ$WSF��8���v��_����΄ ���~ɰLE�}+�<,kt����~��R+�
T���zԔ����.��� ���ί�^�|��2�t�"�̯��eDҔ �޹[�fX�X�^���s@>�����U��#�,��l�Z�>�C���6�G����w�e�*+<|S~�&�!��9)؅�T47q���9M�vd��l@*ˡ�v��#|pR&˻G+��P'c�ՠ���H$*��A�
�RF5��_|A��ۢzS?�z��k˧�T^5� <l��E-�	-�r�D��}�|�y����Y�����( �tg�c�0��/�3�A��i��[����r�QU�ݯӗ����o�ʲ�_v����e������}Ư�dh��U�_k���{���{���?��,�3�HoK���o�u8g�4�	dT�Pi�~,C���� N��	�"���&\�[�2GAާ�g��!�g+<�z��b�:\�e����wx�e�H��G���T�=�T�����Q{:�Z5���k>�	��uK=l��V冪F�a��F�NX�h�5�A�J��X+V-����lsE˅>����5�_�[�!-�&I\%<�yPv���KN�B=A�����q��ņ���mG��\2E�b���;�9+�	%��I��Sbe�gt�0�|�\����J֖6����0��^|f��m�Uo܆χ�ɬK]T'�M1u��9c�,���Å(_Es�i�H��x�|��W"�k��v6aK~'�/#9���E�]�q(�]2n��d��u$o�3�>8�Rz�EIF6��XLJzvc��>�GP;�K����~\�Ǟ;qE���.9F��2�l���D���Q�蘰�!�c��sy�?�ja��f!��0�aU�ŝ!����lP�6tW��6�,�!I(v��ݓ� ,��z_����(aDR]���8vd���ׇ�����R���)��B����(F�/��7&31���=��Lz,�)�,�G�m�z�5�o�L�b��'�N_��@�F�<�[)p�)���I7p��z���)Y�
4�xS�
�T��G��^�	�?Ύe,~��5�P#த�b���΋�u��(�X>⫐�����4�t��(��0P�(���o�^,Z�`��*OV2�Y��O�N��������C5�$� ��m��?3�3�T�t�����.V���C�$r��ʃ�r��Fr��7��X�a=
��<6�y;(eO_�b�z<Ve29]B: �`�	��J��(q/�J��~��]��C�ut,�9�?�Z n����9$t���pq%��RX���]z�8�n�u�<Q����C#��UL�q�$�z\\~�U�-Rz�����,��ظAϊB��6�|�
�h��hU�{�ƨ:A�2$���2��t�xGN��q\Q���A#`��f���K���}ï�J��J~P^�ޯ0�0�̯��E�~�i�� sn�4Ac�v�(����Ԥ��X�/ �?��^>pvx)뻗���;}L���ᾞ�ஜ����o!N�-��ۏ��#���?xkH���Hk(�Dϳ�ȯ��:��EͨrY&�Q�g��0��"�`�����+��\Bx��h��_e]����[�80�#�__�pQ��^7��	�Ӛ���P�
ˤ��/Kw���Ri�Ԣ��1��u٥��TQ�_�O��UǢ�h~~�)P���	�=IV�͒c�k�} h��3�]23���3&V�ӏ�S��p;��
hL�4�VVQ�}����E9��K�85JC�I|7��ܴP�nX(I/ҥr\���˛=��b~�$�9����}Ò_ܷ�{�$Ձ�wA)�e'f0������8�@+�q�hF���F0]��V��Z{�6d���>@�)3��G��++�ƸzxkH�Y؜Udy�`�lp��o���m6��%�f)��,P�A��<�É!nN<%{8���5� ɕP��h��<�e������Ri+w�N���֏�d[��ڒ�~���`��u�I9 �~$�Q�0��}�|���䣲'�ETV&�����P_sU��#rjek��X7Y6�s��Y�m����;5/��X��"a,�q0��``�9��[���@��)��~�2��1ۤAr|%F�m+�3=T�u���!�rG���C�r�ް[u�R\�H0����"���7�L z�z,�N�����nך��ǫ��z������WOV)dM�G�2�~����á1զ
uDQ:��"O�hk1��ڞ��Fx�z8o�M �GH��	E����Z�U�ڬ"p��N� ��~8��c"�ۏ\�c�^n�P?,"��p@e����6��˨�@)�d�>3~r!7�X�_��r��\KW�.dd���4:A� }���r���I7�=!��t_}�:�?����'�êjx<bS�΋P�רoXp����h���P)MW��(���y��,����iJ:�&;
��n�\�"K��͞/�a^���;�&��@�7"s�$��ؾE\-��⢼��p��P�m�-cԽ3 t�҇��q�F�=Ŕ�=�, 䗡O5CS���YltW$-]�9�(�m�J�!b�d��$�:����p_VXf�|wSD�`�c���]�mP3���Ա�r���q�[v|ư�1�����fh�Ĵ^߁ݾ߀߄�K�<؈ޤ�S��<zu�Bwx)*;�x<�KR5��,��&~�L�=���8��9�$�?�d=�)?�NK3~����/��}av��I`7�S�|ee`faY����Ǒ^׺������]7��JR~���=����h���3��J��^�O��#��0���;i@��L�R�:���[�|V����K���:��v����/�cp�!�Z�:�|���S"�ǣ���<�]��T��W|�wՠJ����̺^[���r`Æ�zr:��$H��J�\V�m>6�ΌLr�.��µɃ���s���ү�x�y|n�)	� NޑlY�o�7����cu����D��AKƍ+�mR�a�.�j�E��4�?�0�{�S�}r	}~|ȹ~E)���xJ����=�J�&����7y3	݉Y��y\W���o5�%m��N�J$��;�aez@P�¡Z9�!�
"~2^S>�B�Ϗ��e�U#��ho>�K�X���"H��}���æ���63�T_��bA���>A�22���%Thd�ʴ���F�^R�We�b]���df0��ʹ@�4c9����^9�	���ۘmZ�^�v,Vw5�~�^�џ�a2�e!��O�6Q��ۄ�t{���A��?��]�6)����Sx��^πskd&N ����_!7	F@�i��or��Ac~�@�O{zD��f�r�6�
;��7?:Z�Qa�zS�x�6�y�a9%���l�j�R���:��7��U~U�E�ZR��Tk̾�#_	O"�'�v��+'��K�Q
��=m܋��zu�������
��7~��'`|�(�Y�4��J� �F�����>k����q���8�#�P2{E�z��_$�ЀMZ��/�W��V���5�0>���������r<T�C&���
{}G�d�ܠ���T��C��ޝ��`9�#��u (����w�����yu�����h���M�zG�9��gM6:����\���djfT�=M�*y)4�Rs��`K�tؗS��6ץ�6t�4��/�ō�w��3��Ż zP� ������T�EJ�A��sU-� W�t�n�����1<�� |���e�\Ŝ�	ť�:^��4��"X17�T^_�pٌ-�=�Q�KI�P���t2.�`�3��w��ꤥ�c�^��ҥ_?d��~�g.zm��/�:r�IM�p�џ��Y�@=U��0�-�d
2+K�3:3\֗��cr�Ҫ�D_��� ��P�9����]>���~��ygE�*y�X[�ԌެL�F��tdzhf�b3xya&��{��Uj��cȑ)ܬ������'�h���Tz-W�y��d�� ћ�������?4���'����h��M�u� n"��
c7}7����b�ӢX?2�XB=HI#tɶ�%�����$��[������l�	;�3��5ßZ��5�\�����<Yԏ�X�:��������x�i��j��Ba&�ʇԐ�6��>��M��+��Q�@|i|������0��}�ן}��o;y��M��q��.�F����B��~w^r�@ߞ꬟�}�cM8E.�Pq��XJ�$�Wk[�q���#���"0l�ƻ����)ܒ�z��z�2UH�:�Nʜ��Rd`��I������$�;�N�-���&��N���%PHumLtTi��KG�1����'�qH��5����v/��� �|=4�(ȃ�li�Ǡ�!Q�"�4�f����/E�J��.�эA���ޔu��?_��ʺU��S�}h��(V���v�/P��T�n�nJe�_�f���;��YA�J,�$m?Pi9�Ж��E�v�x��T�,�<l	3{fۤ���#����b��s����zw��N�Ck� ���7�2�zi+�^S�S�_���e����a�mE>�G#8'5�r)��l���~����@��'��V����aI}�8,/�Z�x�0j��?u���	z.9����'RT���>�~Vk�29��L��{H����������������<������������~&��R����Ey��u� &��@��U:��sln�� [�hs.N�#P̷"�|�_r�e1C�������̘�mPD]�>g���*�X�d�����V�䬽?����"���$9�L��$=��V�����.W�PUն�D�U�-|Zb��?�4$7��o����7y��l0��__]BЛg�v�2���*+/��R�%<���<˅XV��ΞC���@�r��Z4�<u��n�.{�5TX[m�pkxۯd���f4�U��1�V/�Z}��I{M� ��?�9Y��e1ry$&�`^����q�=2;�3��NY��)�22n�i�"}�3+�=[�@n�]!��hԟ$�uX��kg66��_�ׇbΗ�Rk9���R%��X�5��Y��L�ءTj�Q/O�R\⃍b���w�N�"5w[��d��&�1T��co�P�bL`�A��sq�#S���F�N�_a�g�3H&s��&��[u8���Jg��G�F_�.:M���6?;�&�Y�������)𞵞�<'��ᅳ�o����W�*d����«�1�� �7|N|�0��NE�<�#���V\�v�ڨƅ+�HY�����ʖf5N<P�Z�NC�A*6���y�����|oh�A�,�zf��P�n�?k䡶7{�9�
�����D�� sh��!:�<A��}� >[D�����2�؜�Ӝg	n�c>h-9��<{q0�L]��.6�}Eݰ�#[��xZH��ڡ5O�Q�].�X���ʹr�]%��s�˛L�g�H�$0���'.�Α.��_F��_��kl�h�o��u�0����7�����U,V$Կ�<�e������p��6(�lc �h&!y��4�4j6$�ȐkD�n��z�U�j� ]�<����*�|�F�F0��5�;�ԣ�
H���No��JL
o�!�*��I�;6�D���b����CM�0�6xI@�e��k���μ��
K�~�݁�$Uf��龜���:wQû]w)�zv�2!�.���=9���.��{T 豝޵�Z�^�̉�C_��&/7W1�P[� sb��i������ӎ�0�(�m���b�F1�Uy��0W�ޏ�\cM
�Rb�?H����Q�1e��&��jZ�����`__�/�W �a-�wt����~SM�9�r���1��
��z�uY������O<5K�@�n���?f`|�
rB���ӛ)��Aǟ��:e���鲏���i��5���r&��u��p�E��Z+P]!O����x=O��hH�^~�úK"{���������u#b�{���ڼi�üO��o4;�m����~7�h����N�`��Ib�&������/�ϯ(H�( �^ג:�PsJ��5�*nr�Nm
�ݫ�wȯ��������m�m�/N6U�%1����ݲ���>��˱�L�+|g�&NVz�jS���|��L_��v�C�4�������XIN,����bf�ݷ\v# ���y��}����¹ۼ�E3e�?����p�A��q���U��:�����7��T1�nD�9Z/I���+�|.�L�Wo3]�C��Ϡ��(��h�#N����-��M���%}�ւsM�=���o�x�d'�1�-ʢ��2?�D���m��:Mm/C9�{B��taԔF��"w����yo�l������r�^xO�OT���9@4Ig�0 ��v����3��D3n�C�Ͽ�z�:Ά�F���B"��u*��������K�$I��g������-VHo���W4;Ǿ�}FZ ��$������^��u~�i][/T4���C���|�E���/�.ȳ�k,����#��SF%Ǎs`Q�[�
o��3���
؀E�� Z,�Y;�a�H/nM���%a.�g�y,�}ރJo$�@~"�&{п�[S���Q��ݴ����0e��9�O
�L���o�}���5��ݏf�E���&Y��|[Pl�V�Jd�o�^Jv:&�i�sC���Rn����V�����`A�� �ZK%����99HV�5.٧�}
�:
��
gr%ݴ����	��#7(a���k�����e殞�F����l%�D��������_�^�+G}�)��D|��)��("[W�`k��b)W�y}v����z�lſ�hآ2ۮ�7�a6��Rt+�*�0h����f�a�%�����?��k���&�o.?�?��$��:�@�U	W��SK.vHL�Nyq�&�`�7o��Mg��4��A����������g�Ή�����,c?��ylBx�ߤ;�*6 �Z�b�8��v�1Ddc�sMU��|d�qA,���f��>y>V�x.(�1�]���vᢌ�k�?�J08me�������4�eziqS�w�w9�m3w�}k�,0�m\7�.@��)������}L�S��Jbq�u�����ΨT	���J
=��a�4s
mWHф��C���m��P5a`>�e3<��R�6��v�^N0uH�Z��*<t�~$�p��͖�����l�F`_�w'�uڌR��ؒ�CA�3���K���,����}K�u���?���	0C����{?BQ�^�t.�kG��;���� �����̶�<��뛅ܱڃ����Q·V����O��B��~�H㽽��ߩ8����:YإS��: �3���˪//
 �,�H��yt�Q�Y�ˍ�� [�i����؊�����.�EaB"��f�9x%/#w�x��/JA�����9�Z{kW���Cfr�/AS��x<�����n���R���H�`K��jh�]u��Z.�2��N��3�O�p+��h2����T�O)'1����
ZЛpny�]����.��S5/��:�,e���b�
��`zPQ1U�cAg�Ta3z0|D���fM��"i�]r�������b���0��� �{h��髳xN4���i��ӝ���+�_���ޘ�$���Nz㞑�D�B.j� �ȴ7��֫۸w�@�~:��������c� 20�v�r�j@Cj%�
�r��G��z�	ZI}M\|�.�L�k��3+��3҇��
��#��yV)�{[����)�S�����+�XC��lUW�*7�����׽�mG��jM��A{����A>�g,5�MHM��A�����s��&�iE=i rX�����=~��Y�zݧ�F��&�T֤tb#o0��!�P��!X)hu�o���7�Vyq���] �<R�ZX]��?r��ˈ���&nSx�a��T��\DE�1�柔a�D)z���ٞ�QA7�����9�ojyl��p�oݭ��C�`��K�W�ѝ�z�\+i�-?�|t�ͰYE�
�l����Q�[;�?�H,�50	5�s'�;N�))芬XuF�j�2C��E��Y2�HwW��exe�I�b ��b����;a����Bs=&[Υ���¼�aҡ-&Nnb:�I>iZ��Cc_�ʞ��Kl�,��[�xeY�|��ڟ������%$����Z��kg�G��l��y�y*z��7��l��2���U���@��~pi��H.!�=?4������g��"��ߩ<j�F~"_��P��~ŨK J"f��n[
�a�Θ-�9�4��r9_��	ڈn&I�s�r�e�'P���Hnz��`V�/��cg�����7�>���i0��_��:�B�7�ܾV�T��]�"��Ʃe$��Usv�<ڂ�zT�"��@=��?'{8`T�Ho)j�@�z�vJ.�ڨ2`�K���.u������3���X�v�g���G�'����M����}n,;�zl�uш�*~t^<�*v�k�zIr#����\�I�d�n�����ɻ��X"8e�Q�Ӧ���lF#�ax1Rt���@�4q���z#�&�p��B�#̿0�Ԣt%Zhj[����7��	�k ��35}_	�Wv{���KO�C
��� �V�3��[�Ct��u^�Z���ƚJ�D�|��R׏.�K'+p�Q4���ܬ��c�o�l8!r���Yt�¼ k-o��=��+O�l�q@<�>���ĳO�6�,Wtc���qr[' G"rs¢���N�PFH�O3��Ab�B��ɮ:5��MB4i���%������n�@_��3��sp��5�����p�ޕ�\��$�+`�xN��U	���$WA���+{�;����o[�/D��Kw��Z��\��e��Nw"�����?yA�k�\5D,���(1�`��|-�/!Ha�rb�X�G�'g�ï��Y�v���u�@rZ۾�3?D���ߎ��2�qSm�iӁ���T�5�aP}����M�9΄�A�^p���s����>��(���*S5��{��R%À�}��9���|�"&%7-O�ُ�G����8��+YbAmL�N"�^�s(�f�Y CT�^��Tt ���ϮP/*����*��	5�J�Xx{���(�HQy�w�R㌭I\t�}2R.�E� �>�$�*�[��̥�L��[o,[ܐ!�c�����R#�S+f���?`�h�j�ţ�GQSM��i��Oo�/#SS�sme� F(��i��J��)�~�Ź7uU��y#�H���X���w���I��-��o�{
Ax����j�9��ɾ9PJ�1�\3aa��}���-�U�cɥzr��0ס\_.~�t�\S\5�����zK&bz>�j��n��K���~p�0{�}��Rm� R3~�G`�g|Cer�9m�R�3�C�\������B�\\RK��S+�n�����]�C4�U e~ش�vi���v�t�����G��ݨ�Az��Y��}Pž�E�kk�\��H����'���'޼�>|�����/lo���v.9�X�e���Es��*t�L�5�:$�\�6�w.���Tm�_�bx}��f���=�|Y�����^�a��z��v���6�w���+��c�e�bI�c�9d+#k����ױ� �����!�k� �@^.�J�����������]`�`:�����>�a�*^o��{�ϖ}�i�<��POJ�j{}�0|@�!V�6�+�G���Y���m�SR ��Ʀ"�NMcF�����lg:�l  �D=������7$�O��9��u�,;�7|e]�	j����2}�ٺ���P�f��w��P�;��Q���CK�叄zy���d����(�x\ H�Y��8�����,��f:�6��qa��Za5� R�Sjͫ��G��T`����eZ2ꬳ�Bp�sO	�0�+�t�)�CnR�ޒ�aDwLU������)H�;,�5hЧ��`��aSR�g�f#�{�b]���*��$�e㗤���n��)_,)����jwP���I�dvQ_iҵ2�g���V�!_��L�_y׶����F��$E�O�	��rX����!�fg �=J�����K����Aă�b���L�����i�T~��#:�}�QK��)vkх�yo�w��#N���+�Zy����m��/'��\/=~��r&����P�Z��\t����%����E-4�\b���<�Q��t���S�_.`7�[�G��%�C��a�96�#�u��W��L��P�gE�9�L�
1��R��l�|6�io�m C�����YB���2Q�,h^1t��_E��@`r���dUG1�m�	45Q�����C�{�9������j��ا��R����p7ю��\�sŃ��LM/��N�s�j�|֍����XR��B�`��!�^�ڂ�q(���ԩ(g3��u�G��-�1x;ڡ5˩�y�i����.�����s9�̒�F�U"M�������u�����#)���F:���	�jlʓ���뽘�o��Y���s<��Z�֦hJr7Q'�gA2���������Ih!�,:�\q�"=��1
ͼ7�v��tf�f�P�IA>�\�W��Z�G ��.?�]�z@���N/*�$0?."ZF������g'7�,�im�^�>����Hu��F����q8��	Fa����_G��V��B�P��\啃�#Ʉ (O��z@i���
G���Ү���:�q�3M/�
Ab���&�U�KfU���̾Bų�:ER���
m����"��������3��⨉n;�3Ze�@*�]�M1M��%jT-��~�0T�]2�#�ُ��zh��V9<S�a�����VM绳����8q��/{�s&(aEiR�҄Cdi1���ܨO�.5z�ic��(��B���R0����FǱ^��C8�'��8-i�;�K��9��]����t���?����dFYn�6�F2|o�]9���C���fw�2�]�'s��_z�3]ڧ�%��f*��$���4�]���g/�������<qb��xy����Z
�qL�dUշ�ު�ٻ�ȯ����"O��%Ӡ�}ѓ6_(z|@��Q>t�=�FF҆���p-)P�>��Q��V>E�s�#zb̛��0
�W�W�<�L�k9,��j�za�2h��"o�ȬL�H�0�Ӡ�)1@��f���zG���>%�����٭�	�S�v@B=i;Z���zb���qb��[K+�qtS�)��~�GXwlH�L�i�v!0���I�Ǘ�0W����[=���;龧w����ܭ�z/�/���Z����5j�qYP<�5䃁����&�R{0�1�&�+�D�������M޼n��T�#��ӡ��z��u�Pa`����+�Ji��G��He��t��yR�4�?2��Gf()̗4�^쥥BwL��>�J��|z���p�oPD�K�\yk���}q�P�� �Ai/Н���U�����Z�+�&KN��;�g�wMM;ԝz�JKD�DZtߟ��g�����@jQ4�L5���c)��E|��D������w	�`���i�c�^�o�S�/�>8�0X@|��%�D�Ѥ��	��!N��k>��e��L�����P�`���I�7�KK�(����كkc��)�d�6(���`y-�<��^x��zT+�-'n�ǹ(Y\��0����'�ɦs#�; �2�]�fL�f#�k"7��Pj���+��̦�c�[mILx��~N3���Q�YK�s�\�����?s/������Ż^e�'�pG�1��1�gZX�ȏ��
���le�&DN�C��M�/+G�|Ƭ \)��� m�i��Z6^&����7>~�)ʐ�"@��sؙ���#Q�a�#w��V�sb|�a4���$c������K%�h)����T�:"�xE#��Z��ƕ�a �{���-E�v�:��I$���ݟ�HZP��qQE4y<Y�c%a5���,l��WYj���2�{4�$�����z+%���L��@�^G�!�%g����?�60�h�AH��9�ĳ��T쐞+O޵2�RV�ߐ"֓���3��&a���ת@ꠦ��54��/�$��2��Q�BZce����	F�@�8K��wG��+�d���egu3~�[C�ȩu�;i���뿓���5�װ��G�yJ?����K�ߔq���͈/}&8��3���h��_'��?���JLZ�}��4� j���;���O)���i������>|@�������Sy��K������ʈԌ��tS�ekj�L������D	ʄ��S�\#) GnS��Ĥ� o�f2a1�`��q�4�rO���q!^�\Ķ�IA�똍$��}.����Dd��&�cZ
<�ئ��T�7;'�1`m!GJ픾�� �aˏ�};��~���L�[�sZ�;�(D@ҥP}�fݱs�	r�y�HGB��q5���0����	��Ů{�4z��[%�S9�dJ�{a/g�4RF��q��훠$'8��.�^΂�n�t�R�ۏB�C��x�c�h��2V�]\���!H- P_�7�XP��d�7�+O�Bi5Z���=��՜Xgp���ZRB��q h��&	��l�e<�x��U�u��V�<���qT����㕂7krc����*���8��^�ze5b
ڻO\����R����6685�1��
h����M!gHk�VJqY���8�Aݐ)��87��%�w�]�5NFCS�L����ڣ�R��j�<0Ԫ��^5�C�Q*�L2&gaɋGn)l�v�"08Z������O�}�-�I6���92�v&��n}�yF���K��u�Q3���>	7��т��p9�c7/ڏ���w_�Q*��Hv6~���ӏ����G�K8��C<�Ms`���_��\�6������X�%��)���J�� p/�X�W�$Zd:'G,�7�t��{���V'6-V/���8`���nZ t��Γk_x�������נ�d�/�"���U��#�X��L��6x\bB����^"X�K�����d�|Dz� W�v����An��;\�~%`q��,^����<�� o��5��1u��g�/%đ*��@�}��K��|�ԍf]�PX+��A%7PG��v<<��9����{�ȋ@��^�.oЇQ��lsSb54�*��M00��T1�=�$�~�/��~������p[�λ�x�3�)K�,�E]s� Y��fː>���� e>��4��(r���T���p ��-��Fh�<8�_���󰷷[�T�&���1=�˩Y~���J�&�)
�9�"0�N����*�?�	�b�v%f�c��x�KA���jt����VhH�6��3�3�~��[ ��sl�� ��3�C��6SW���	�;g���XI������L_�M0snjL��37,	�mi�8���3�/ɛ�hH��}[
�,�c����<}`Ķ��_�RX�T�������s�Uw�?��ԇ*����w���m� �G=�v��te-�3H>JF9#r��EM#&�$*�6_�m,8�&���C#݋�j�S=j�,��#U�r�+�����0���=�G���r��E_q�T�eAK�U�,���)���a�