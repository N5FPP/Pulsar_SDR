��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY9?�C�><�Ǌ9�O�
3��9������3KA�rԨd�/.-�|�3�ߐ���NE*���]Al�y����i���K����}�$�v�l��X�D3nh2n/Z��xvnKZ�No]���n6��d>�2(b#`Sɠ�9}�I=��;L�AA�g��$��z���\%�p.���J+yy[��7A�M�`�`��|z�r?�q�Mc�#v�$�e���=��$#5+�}��P�������J�;�C� ��ؖ�|%�)0t�Y#�#w=4��"a`9�X���k*zYOU�u�8�������9
Cd@8ޜή�#�u���B�cu	�:6�q�H!�W��D�������{lĻVrC�r��ךc���}�'�㠗���=p��n��C�iͺ虣۩%����>"��-NT��0rI�g�(#�LK�+������Hh��<5�j�Hh$ ���F4H�d����$�d��|0�sy�^r��$��؊�Q������q�`�$7�@U��v�|���Sҽ��~�U�s|rN�xоUn v�=ƶ`�"H��W
Qr#�l_�;��y��c}n�a���}7͗��3E|���������/H�C�#]���L+T1H������m����h�C�L��"���b�
Cɠ��@���j��;{�_�S}E���t����	;�y�m�0�	�׉51*�쯵Lݹ�����ŒV�R�|3��F��Z�Jՙ�|�&��,w��8ogZ{�3�u��	��z"��Rl%�WΕv^��;�����Z�N���cq��{�����0�
�(d}F�S�,!W��T�|�����
C��t4���)Gy�8b8�U����{M�x]��Y�=�o�9�A[GIs�ߣג��v�~� ��w�h��E�4gj1˰)c��3*�ZV�VA,,$��S�M�F���� �؅���y2㵏��F�Ȫ���4����5\�>o�i�na#�]��
sK��T���4�7@)��W����� [ K�[�k��%6���1=;����ެU(r����d)u�z���Ό��:%F�'��_�� ������6m���>�\��y��R4�Z۩�]#�Q��0l�ސ���΍�G��Y�wht:.�`�AǨݶ�590F��4���
��?�S�MjFr*]�{�n,ݱ���F� ڷ� &�)A����������ܧW��NX�(�֎����s�����|*�		�F9�˻m����/��A��Z�W�A^�L��@* �n]�H�m}}�r�:c�����E��i�Q�;�	�ZY�B9��U�6�_7�Waτ�9S��Nm'G� ���q/ն�.!�Z��SUxv�5�t�O:�z�ɷ�v<7>�	=s�b�g�>����/X7���� �M���-;�`�o�9^�_�		��	���f��@Z��Op��_D\u�=�yU���22˺, K�`�_��N�C��e0����lO6zs�AƗSE1̅]�#d��gA��|�R��"7�'oZ?��]��뜲�