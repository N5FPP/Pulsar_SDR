module altpll
#(	parameter	bandwidth = 0,
	parameter	bandwidth_type = "AUTO",
	parameter	c0_high = 0,
	parameter	c0_initial = 0,
	parameter	c0_low = 0,
	parameter	c0_mode = "BYPASS",
	parameter	c0_ph = 0,
	parameter	c0_test_source = 5,
	parameter	c1_high = 0,
	parameter	c1_initial = 0,
	parameter	c1_low = 0,
	parameter	c1_mode = "BYPASS",
	parameter	c1_ph = 0,
	parameter	c1_test_source = 5,
	parameter	c1_use_casc_in = "OFF",
	parameter	c2_high = 0,
	parameter	c2_initial = 0,
	parameter	c2_low = 0,
	parameter	c2_mode = "BYPASS",
	parameter	c2_ph = 0,
	parameter	c2_test_source = 5,
	parameter	c2_use_casc_in = "OFF",
	parameter	c3_high = 0,
	parameter	c3_initial = 0,
	parameter	c3_low = 0,
	parameter	c3_mode = "BYPASS",
	parameter	c3_ph = 0,
	parameter	c3_test_source = 5,
	parameter	c3_use_casc_in = "OFF",
	parameter	c4_high = 0,
	parameter	c4_initial = 0,
	parameter	c4_low = 0,
	parameter	c4_mode = "BYPASS",
	parameter	c4_ph = 0,
	parameter	c4_test_source = 5,
	parameter	c4_use_casc_in = "OFF",
	parameter	c5_high = 0,
	parameter	c5_initial = 0,
	parameter	c5_low = 0,
	parameter	c5_mode = "BYPASS",
	parameter	c5_ph = 0,
	parameter	c5_test_source = 5,
	parameter	c5_use_casc_in = "OFF",
	parameter	c6_high = 0,
	parameter	c6_initial = 0,
	parameter	c6_low = 0,
	parameter	c6_mode = "BYPASS",
	parameter	c6_ph = 0,
	parameter	c6_test_source = 5,
	parameter	c6_use_casc_in = "OFF",
	parameter	c7_high = 0,
	parameter	c7_initial = 0,
	parameter	c7_low = 0,
	parameter	c7_mode = "BYPASS",
	parameter	c7_ph = 0,
	parameter	c7_test_source = 5,
	parameter	c7_use_casc_in = "OFF",
	parameter	c8_high = 0,
	parameter	c8_initial = 0,
	parameter	c8_low = 0,
	parameter	c8_mode = "BYPASS",
	parameter	c8_ph = 0,
	parameter	c8_test_source = 5,
	parameter	c8_use_casc_in = "OFF",
	parameter	c9_high = 0,
	parameter	c9_initial = 0,
	parameter	c9_low = 0,
	parameter	c9_mode = "BYPASS",
	parameter	c9_ph = 0,
	parameter	c9_test_source = 5,
	parameter	c9_use_casc_in = "OFF",
	parameter	charge_pump_current = 2,
	parameter	charge_pump_current_bits = 9999,
	parameter	clk0_counter = "G0",
	parameter	clk0_divide_by = 1,
	parameter	clk0_duty_cycle = 50,
	parameter	clk0_multiply_by = 1,
	parameter	clk0_output_frequency = 0,
	parameter	clk0_phase_shift = "0",
	parameter	clk0_time_delay = "0",
	parameter	clk0_use_even_counter_mode = "OFF",
	parameter	clk0_use_even_counter_value = "OFF",
	parameter	clk1_counter = "G0",
	parameter	clk1_divide_by = 1,
	parameter	clk1_duty_cycle = 50,
	parameter	clk1_multiply_by = 1,
	parameter	clk1_output_frequency = 0,
	parameter	clk1_phase_shift = "0",
	parameter	clk1_time_delay = "0",
	parameter	clk1_use_even_counter_mode = "OFF",
	parameter	clk1_use_even_counter_value = "OFF",
	parameter	clk2_counter = "G0",
	parameter	clk2_divide_by = 1,
	parameter	clk2_duty_cycle = 50,
	parameter	clk2_multiply_by = 1,
	parameter	clk2_output_frequency = 0,
	parameter	clk2_phase_shift = "0",
	parameter	clk2_time_delay = "0",
	parameter	clk2_use_even_counter_mode = "OFF",
	parameter	clk2_use_even_counter_value = "OFF",
	parameter	clk3_counter = "G0",
	parameter	clk3_divide_by = 1,
	parameter	clk3_duty_cycle = 50,
	parameter	clk3_multiply_by = 1,
	parameter	clk3_phase_shift = "0",
	parameter	clk3_time_delay = "0",
	parameter	clk3_use_even_counter_mode = "OFF",
	parameter	clk3_use_even_counter_value = "OFF",
	parameter	clk4_counter = "G0",
	parameter	clk4_divide_by = 1,
	parameter	clk4_duty_cycle = 50,
	parameter	clk4_multiply_by = 1,
	parameter	clk4_phase_shift = "0",
	parameter	clk4_time_delay = "0",
	parameter	clk4_use_even_counter_mode = "OFF",
	parameter	clk4_use_even_counter_value = "OFF",
	parameter	clk5_counter = "G0",
	parameter	clk5_divide_by = 1,
	parameter	clk5_duty_cycle = 50,
	parameter	clk5_multiply_by = 1,
	parameter	clk5_phase_shift = "0",
	parameter	clk5_time_delay = "0",
	parameter	clk5_use_even_counter_mode = "OFF",
	parameter	clk5_use_even_counter_value = "OFF",
	parameter	clk6_counter = "E0",
	parameter	clk6_divide_by = 0,
	parameter	clk6_duty_cycle = 50,
	parameter	clk6_multiply_by = 0,
	parameter	clk6_phase_shift = "0",
	parameter	clk6_use_even_counter_mode = "OFF",
	parameter	clk6_use_even_counter_value = "OFF",
	parameter	clk7_counter = "E1",
	parameter	clk7_divide_by = 0,
	parameter	clk7_duty_cycle = 50,
	parameter	clk7_multiply_by = 0,
	parameter	clk7_phase_shift = "0",
	parameter	clk7_use_even_counter_mode = "OFF",
	parameter	clk7_use_even_counter_value = "OFF",
	parameter	clk8_counter = "E2",
	parameter	clk8_divide_by = 0,
	parameter	clk8_duty_cycle = 50,
	parameter	clk8_multiply_by = 0,
	parameter	clk8_phase_shift = "0",
	parameter	clk8_use_even_counter_mode = "OFF",
	parameter	clk8_use_even_counter_value = "OFF",
	parameter	clk9_counter = "E3",
	parameter	clk9_divide_by = 0,
	parameter	clk9_duty_cycle = 50,
	parameter	clk9_multiply_by = 0,
	parameter	clk9_phase_shift = "0",
	parameter	clk9_use_even_counter_mode = "OFF",
	parameter	clk9_use_even_counter_value = "OFF",
	parameter	compensate_clock = "CLK0",
	parameter	down_spread = "0",
	parameter	dpa_divide_by = 1,
	parameter	dpa_divider = 0,
	parameter	dpa_multiply_by = 0,
	parameter	e0_high = 1,
	parameter	e0_initial = 1,
	parameter	e0_low = 1,
	parameter	e0_mode = "BYPASS",
	parameter	e0_ph = 0,
	parameter	e0_time_delay = 0,
	parameter	e1_high = 1,
	parameter	e1_initial = 1,
	parameter	e1_low = 1,
	parameter	e1_mode = "BYPASS",
	parameter	e1_ph = 0,
	parameter	e1_time_delay = 0,
	parameter	e2_high = 1,
	parameter	e2_initial = 1,
	parameter	e2_low = 1,
	parameter	e2_mode = "BYPASS",
	parameter	e2_ph = 0,
	parameter	e2_time_delay = 0,
	parameter	e3_high = 1,
	parameter	e3_initial = 1,
	parameter	e3_low = 1,
	parameter	e3_mode = "BYPASS",
	parameter	e3_ph = 0,
	parameter	e3_time_delay = 0,
	parameter	enable0_counter = "L0",
	parameter	enable1_counter = "L0",
	parameter	enable_switch_over_counter = "OFF",
	parameter	extclk0_counter = "E0",
	parameter	extclk0_divide_by = 1,
	parameter	extclk0_duty_cycle = 50,
	parameter	extclk0_multiply_by = 1,
	parameter	extclk0_phase_shift = "0",
	parameter	extclk0_time_delay = "0",
	parameter	extclk1_counter = "E1",
	parameter	extclk1_divide_by = 1,
	parameter	extclk1_duty_cycle = 50,
	parameter	extclk1_multiply_by = 1,
	parameter	extclk1_phase_shift = "0",
	parameter	extclk1_time_delay = "0",
	parameter	extclk2_counter = "E2",
	parameter	extclk2_divide_by = 1,
	parameter	extclk2_duty_cycle = 50,
	parameter	extclk2_multiply_by = 1,
	parameter	extclk2_phase_shift = "0",
	parameter	extclk2_time_delay = "0",
	parameter	extclk3_counter = "E3",
	parameter	extclk3_divide_by = 1,
	parameter	extclk3_duty_cycle = 50,
	parameter	extclk3_multiply_by = 1,
	parameter	extclk3_phase_shift = "0",
	parameter	extclk3_time_delay = "0",
	parameter	feedback_source = "EXTCLK0",
	parameter	g0_high = 1,
	parameter	g0_initial = 1,
	parameter	g0_low = 1,
	parameter	g0_mode = "BYPASS",
	parameter	g0_ph = 0,
	parameter	g0_time_delay = 0,
	parameter	g1_high = 1,
	parameter	g1_initial = 1,
	parameter	g1_low = 1,
	parameter	g1_mode = "BYPASS",
	parameter	g1_ph = 0,
	parameter	g1_time_delay = 0,
	parameter	g2_high = 1,
	parameter	g2_initial = 1,
	parameter	g2_low = 1,
	parameter	g2_mode = "BYPASS",
	parameter	g2_ph = 0,
	parameter	g2_time_delay = 0,
	parameter	g3_high = 1,
	parameter	g3_initial = 1,
	parameter	g3_low = 1,
	parameter	g3_mode = "BYPASS",
	parameter	g3_ph = 0,
	parameter	g3_time_delay = 0,
	parameter	gate_lock_counter = 0,
	parameter	gate_lock_signal = "NO",
	parameter	inclk0_input_frequency = 1,
	parameter	inclk1_input_frequency = 0,
	parameter	intended_device_family = "NONE",
	parameter	invalid_lock_multiplier = 5,
	parameter	l0_high = 1,
	parameter	l0_initial = 1,
	parameter	l0_low = 1,
	parameter	l0_mode = "BYPASS",
	parameter	l0_ph = 0,
	parameter	l0_time_delay = 0,
	parameter	l1_high = 1,
	parameter	l1_initial = 1,
	parameter	l1_low = 1,
	parameter	l1_mode = "BYPASS",
	parameter	l1_ph = 0,
	parameter	l1_time_delay = 0,
	parameter	lock_high = 1,
	parameter	lock_low = 1,
	parameter	lock_window_ui = " 0.05",
	parameter	lock_window_ui_bits = "UNUSED",
	parameter	loop_filter_c = 5,
	parameter	loop_filter_c_bits = 9999,
	parameter	loop_filter_r = " 1.000000",
	parameter	loop_filter_r_bits = 9999,
	parameter	lpm_hint = "UNUSED",
	parameter	lpm_type = "altpll",
	parameter	m = 0,
	parameter	m2 = 1,
	parameter	m_initial = 0,
	parameter	m_ph = 0,
	parameter	m_test_source = 5,
	parameter	m_time_delay = 0,
	parameter	n = 1,
	parameter	n2 = 1,
	parameter	n_time_delay = 0,
	parameter	operation_mode = "unused",
	parameter	pfd_max = 0,
	parameter	pfd_min = 0,
	parameter	pll_type = "AUTO",
	parameter	port_activeclock = "PORT_CONNECTIVITY",
	parameter	port_areset = "PORT_CONNECTIVITY",
	parameter	port_clk0 = "PORT_CONNECTIVITY",
	parameter	port_clk1 = "PORT_CONNECTIVITY",
	parameter	port_clk2 = "PORT_CONNECTIVITY",
	parameter	port_clk3 = "PORT_CONNECTIVITY",
	parameter	port_clk4 = "PORT_CONNECTIVITY",
	parameter	port_clk5 = "PORT_CONNECTIVITY",
	parameter	port_clk6 = "PORT_UNUSED",
	parameter	port_clk7 = "PORT_UNUSED",
	parameter	port_clk8 = "PORT_UNUSED",
	parameter	port_clk9 = "PORT_UNUSED",
	parameter	port_clkbad0 = "PORT_CONNECTIVITY",
	parameter	port_clkbad1 = "PORT_CONNECTIVITY",
	parameter	port_clkena0 = "PORT_CONNECTIVITY",
	parameter	port_clkena1 = "PORT_CONNECTIVITY",
	parameter	port_clkena2 = "PORT_CONNECTIVITY",
	parameter	port_clkena3 = "PORT_CONNECTIVITY",
	parameter	port_clkena4 = "PORT_CONNECTIVITY",
	parameter	port_clkena5 = "PORT_CONNECTIVITY",
	parameter	port_clkloss = "PORT_CONNECTIVITY",
	parameter	port_clkswitch = "PORT_CONNECTIVITY",
	parameter	port_configupdate = "PORT_CONNECTIVITY",
	parameter	port_enable0 = "PORT_CONNECTIVITY",
	parameter	port_enable1 = "PORT_CONNECTIVITY",
	parameter	port_extclk0 = "PORT_CONNECTIVITY",
	parameter	port_extclk1 = "PORT_CONNECTIVITY",
	parameter	port_extclk2 = "PORT_CONNECTIVITY",
	parameter	port_extclk3 = "PORT_CONNECTIVITY",
	parameter	port_extclkena0 = "PORT_CONNECTIVITY",
	parameter	port_extclkena1 = "PORT_CONNECTIVITY",
	parameter	port_extclkena2 = "PORT_CONNECTIVITY",
	parameter	port_extclkena3 = "PORT_CONNECTIVITY",
	parameter	port_fbin = "PORT_CONNECTIVITY",
	parameter	port_fbout = "PORT_CONNECTIVITY",
	parameter	port_inclk0 = "PORT_CONNECTIVITY",
	parameter	port_inclk1 = "PORT_CONNECTIVITY",
	parameter	port_locked = "PORT_CONNECTIVITY",
	parameter	port_pfdena = "PORT_CONNECTIVITY",
	parameter	port_phasecounterselect = "PORT_CONNECTIVITY",
	parameter	port_phasedone = "PORT_CONNECTIVITY",
	parameter	port_phasestep = "PORT_CONNECTIVITY",
	parameter	port_phaseupdown = "PORT_CONNECTIVITY",
	parameter	port_pllena = "PORT_CONNECTIVITY",
	parameter	port_scanaclr = "PORT_CONNECTIVITY",
	parameter	port_scanclk = "PORT_CONNECTIVITY",
	parameter	port_scanclkena = "PORT_CONNECTIVITY",
	parameter	port_scandata = "PORT_CONNECTIVITY",
	parameter	port_scandataout = "PORT_CONNECTIVITY",
	parameter	port_scandone = "PORT_CONNECTIVITY",
	parameter	port_scanread = "PORT_CONNECTIVITY",
	parameter	port_scanwrite = "PORT_CONNECTIVITY",
	parameter	port_sclkout0 = "PORT_CONNECTIVITY",
	parameter	port_sclkout1 = "PORT_CONNECTIVITY",
	parameter	port_vcooverrange = "PORT_CONNECTIVITY",
	parameter	port_vcounderrange = "PORT_CONNECTIVITY",
	parameter	primary_clock = "INCLK0",
	parameter	qualify_conf_done = "OFF",
	parameter	scan_chain = "LONG",
	parameter	scan_chain_mif_file = "UNUSED",
	parameter	sclkout0_phase_shift = "0",
	parameter	sclkout1_phase_shift = "0",
	parameter	self_reset_on_gated_loss_lock = "OFF",
	parameter	self_reset_on_loss_lock = "OFF",
	parameter	sim_gate_lock_device_behavior = "OFF",
	parameter	skip_vco = "OFF",
	parameter	spread_frequency = 0,
	parameter	ss = 1,
	parameter	switch_over_counter = 0,
	parameter	switch_over_on_gated_lock = "OFF",
	parameter	switch_over_on_lossclk = "OFF",
	parameter	switch_over_type = "AUTO",
	parameter	using_fbmimicbidir_port = "OFF",
	parameter	valid_lock_multiplier = 1,
	parameter	vco_center = 0,
	parameter	vco_divide_by = 0,
	parameter	vco_frequency_control = "AUTO",
	parameter	vco_max = 0,
	parameter	vco_min = 0,
	parameter	vco_multiply_by = 0,
	parameter	vco_phase_shift_step = 0,
	parameter	vco_post_scale = 0,
	parameter	vco_range_detector_high_bits = "UNUSED",
	parameter	vco_range_detector_low_bits = "UNUSED",
	parameter	width_clock = 6,
	parameter	width_phasecounterselect = 4)
(	output	wire	activeclock,
	input	wire	areset,
	output	wire	[width_clock-1:0]	clk,
	output	wire	[1:0]	clkbad,
	input	wire	[5:0]	clkena,
	output	wire	clkloss,
	input	wire	clkswitch,
	input	wire	configupdate,
	output	wire	enable0,
	output	wire	enable1,
	output	wire	[3:0]	extclk,
	input	wire	[3:0]	extclkena,
	input	wire	fbin,
	inout	wire	fbmimicbidir,
	output	wire	fbout,
	output	wire	fref,
	output	wire	icdrclk,
	input	wire	[1:0]	inclk,
	output	wire	locked,
	input	wire	pfdena,
	input	wire	[width_phasecounterselect-1:0]	phasecounterselect,
	output	wire	phasedone,
	input	wire	phasestep,
	input	wire	phaseupdown,
	input	wire	pllena,
	input	wire	scanaclr,
	input	wire	scanclk,
	input	wire	scanclkena,
	input	wire	scandata,
	output	wire	scandataout,
	output	wire	scandone,
	input	wire	scanread,
	input	wire	scanwrite,
	output	wire	sclkout0,
	output	wire	sclkout1,
	output	wire	vcooverrange,
	output	wire	vcounderrange) /* synthesis syn_black_box=1 */;
endmodule // altpll