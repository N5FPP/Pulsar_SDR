��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY��UYO�[<8�;�G�@��5۩\lD���~��D���S
�)�$)�'�гtW�Yu%_J�S�&&���d��/T=9�y���R�+N2����o������E��=�08V�������`�q	"]+�G�[����H�$@iw��������K�	�_�C�DUw볛6z��wR.~����jcZ-��o�{(�G<�	���B���\�_	־ߋV%:/y8�J$x8յ,s��߇��OI�����\�r�:u�ks��Y&���Su��+����cX]��WP�z�a��6�+���]�����eB|�2߯Z���9#���C�~t��x����1��ঋ�) �'`�	.����*�L^�cD�A�	".Fn�t�ĳu�J�S#�|ǔ|{���Ɛ�k����8t������v������,�~H��0Ra��{�I�2_���9:��1\.�m�rn+eE��e�#7�W�у�m�W���Ϙ�	�:|�T�&�ԏ���u�f�\��j�ZP�.e�Ϭ�RJ�g��5�b5!��۬�)��8X�9��eJ�&w��e���ᮾM������L}r_}�Y�7��S�s�!qڠFT�ԡ�������S�z'}��<�I���,o)L��5�W�U�����c����<F�=�pU�;h�'���Y����F�!u���C��l�%��so�DI��ul��跶�kp�D/��@��+��/�|���'+�;���n�et2��I��V��fb&�K�2�l[ �V�;Ѡ�;���Ɩ75m^����=�e���ъW���h�-!����q(� s�3ߢ�ȵ%\�z�zĬ��: � �f���������K��4��(�f�X��gՎ�WJv۩�W�31��k���&�9���m�������3�쩌m�;�0���/��	�PQ\��Zҗo��d��P��1��{�z����-�Jwߺ ���\KX�p�V�d"C<H9(z���:=ͻ62�1�N�B��AQ�$'������Y�PS�i����79,�	�7���[R�NV���A�o}�@����徊���禱���w�U'2��ȌX���,W�5��2��	�ڲ-�3��: �V��V��̽�Y� a��`�q�.U5A�@(����S��YIp�,���:�����ퟚ�np!�<�Oa�'���#��M֛i9ӱ�rB(��.��1���HoF�T6�����mé��E�@Z��'T\�����O^VZһ����<�F8�TM`ȫAK�\�G?�l�<�T��D��L窔���=���|��.%�^�V���z�"�Q*��]l�]�l	���%��b_  ,r"ٯ,�(������a,��y(�n�$\�p����mIĊ�L�@��(l�$Btj-��Tl` ��c�u��IAòݔ�7�٪�hʚ�,=�h%Q�\�Vij �ޔ�<�B�/~�#F}�W�l�|:�^,h3��8�93�hGgN,��^B�t�81�k�\u�Vb@l
����f�ଁqE��
�{���.I�S3HiK�5�2������؈�󩸻�b>U��?��|pj��K�3�15Ҽ�}�_��YX���l8so��"�w�8ϿX��:�l��G�3G�R�Tj����3IF�@����Ҵ~�f:1΍b�Z
ܿ&�IF����8"5��@h�����
<�Gh�R ������-5v��2�2���z�.PSb�n�VE�F�_��8�K��� �+kn����A���J6�J��+��	�t9�AJ4�q�6]��63���B��r��҆��V���ύx�����x|�S��)t��p�Y�ճ	A�
xԟ�j|D�t����ZI�(nu�HR��0�v);�(�������GH��b��Q	]���*�J���gYSJ��ݽd��n�%��$qb�	!k-\Xr���R%�7����.�k4��|����� zϻ ��I���P�b{	-e�MK�F��i�O�%j'�n{��]]�4�0h�=��T�����`�[0�r��|��tT�t�b�7㤖\�4���Ec��2R�T������'�2|6q�،�A�N���O�mA:s[�@��a�x6G?#Ǜ�x�6�N�����c��؟Qߪ�$�	*�q
,��ЛH�c�%�L��QB�7R/J/��F�k3�N�Z�4���4#4*��p�j�'%9�i��?'�����U��uQ;��

N>E�����Y�1�^��d9�����.���x�t�S�R.�Q�9T���h9����gW��c:n�]��T|$!�o����kp�0��F�'~�9&2�������S2���܍��5���M���c�^-��������~��e��X>���]R���O�{,�)�\�K�g3c������J���V�QUA�!l2�	��ȩ�G�ɼ���1���=tn���{39���c���[��F����[�ծKDZ������IxTa@_`%�#�J�R"�rlDG�'��`��D��6yJiq����y'�|� 1]z�a���>�pZ�8K7p&��O_�i�x����l�]����n��i3R׾�ZnI4�[�;�����B�`+���<I�圍��n�鞑Y�хo���/8V�ї�~��� R��9��&�{�VNI�얢�D�A\���o(^U�.��G�_��	Q��_1X]WL=��t-n�D��A�̙��,�@�z3|�V���V��\5���IV���d9An��ѱ� �T�H#&{��{��/��A�4R�����<��j'��~
FEpD��
��Y?�.8�?�����or�`v�.K�"d����|�\�c;Uo��*�Vw5�`���vP�]�_�`��9�Q9�����h��+� ��+�JB���U���̊'�G�K���8�	�Gz.�F1�j{��Ʃ��4_�����W��|ќ�;��h�Up�����ճ�\��<��?6����|GYoFn�0��r�A��MCM��07%���8��Gt��{5����!x'50�N�,���@ aqd�\\��)�3P"�����<�#��E6�����
ţ��G!
$C���Ty�%���TO��I,�X���v�?�ȷ�*�l�)!|#y�����D�1@��T|���x�T�v;b��j�x���-��Qd@+m�\MzNF?v�����1`{M�0|Yڷ�kh�m�*>�x�9Cy�t�ti�Ȗ�[��Xɤ���}Q(N��K�DJNF�a�e�1��*=t�o�4�*���؄�+�a�\A���R�K���/^9��M�Y���k��f�О�������n]Nf-7!t�}�����cθ��
Yh�]�j��Ȏ���\g�@f��a}~1�c ��Np��_��8p(��~4:<[�x�p�#35��������e��Ϟ����`^/�+
��Ю����L+�I�(,As{�qV��=����SR'�=����F?�')�κ���������^꿇2 �zS�Q��*b+�l��|#:�m�{�U��f�J#�栁���1l1e.7���BDQ�s��4�+�|��-�y����z��!H� B���v/�}o��sD4����[ƿ�t�)� Ɣ.Q12�Ѡebk=bR����EV!���F6܉]E������֐��ђ����u<�x�ʕO��O(�ѿ�����؍!"8�X^��b���1�F���v��OX<����F�tr>Ԑa�p1�zY�/(����{�e/�X'�v�Q�uV��"=I"(�,a�̼SH��O�/�֬�*�����Z��(_�X����%�tY/"GO.��Zܝ�+������w���m�j��@�F��I����_��C�W�^YÞ(;w\�A���n�d��5�;Ѭq�wr@o�9�!��g�V��.��D8��%	&���l��g��cէqo^��7=�6RY���/+���a~�ݳ�Z*����tV ��_�գ ���r�@���DJ�)(q��TCJ]�$1����ĞX���T, ��� >#�P8���ei��dC,f��dQ�m�A��A�[t^I�DN��%���Q�H.k�*���0/���/�D5������wY1�W�7�B趉���)�o�w�s
��EQo�sJ6��`D��t?�ĉ��b�<�	i���t��G5]-��8�z| ����u�{B,`��_A�ѩ��߃��'����٬�GR���m��n��m�w�EyB�ܖ�L*a�s�)I����r�jLr9]�:��@�	)��3r��<z�ǭ�0r~�M���t)���:Rm�k9�����ΎsvP�R�N�n ���.���&iz�xфc��E����h�i*	���i`�4�ë�7w;�3��`�4�.�0���G��3y���x�8/��j)��c��0J
�l�gfy��� x�%�4[��QD%�[�սL�8�3	���eżݓ޿u��qh�n;�T>Ǭ���6�X��$?SYRK����ۓ���	o�B��� 4:� @3!H/֕���	��ѭ��~�	����优2'��<e��"Kx��x �2��G��T��͆B��-<����~�	�+x4�B������z�bի��L�I�F�I-\9(bv������j	�0˟��!p�T���wNZ�v)���"@Uz�z�*��f��� �rve��|(��oܛ������ʿ|A��~
�=�?>��W�N9/�c��Af?q������T?}?�ͣ�R������W��_��Sw��#��IG=����O�U�/_8�\���E�7;�w�IH	��4a��v���e����yn�����k�w3����"�FJ�X&7�QA������`
d��hc�=nI� ��Y_�I��&�{g��R�h
2�t?^��Ҷ��{Lq��B^��[�W4���������g�)�xx�q���{e/�[�DX�wd�*�.���*�qp �p޺Sp_9=Y���Fy�ȵ��T/�@�@��	�����0�-���h2P�Xy� � ϳЭ<���Nu�˄�ѤB�I�%`�$M�������Ơ>���� ;�1��%<�|7	Y(�5"�'�zy \���d�R�	��QFl�m|k��"�����a�NC�7��
���0k%��ّ�D�����,�#S��y���ռ���`�a�#��x��^ �hB�R�Q8QK�����
q# �ݒ�Uf�s��I�\
�t]�\�$���]8w7S\��J6f;[����<.����`�F�*>f{���k���.T�28�����i�-�^�D��m�nۀP����q�(�g@<*�X��$����׆sp�b�:h9���q���P���>;��,ϭ3WJ�n���O�6�I[�'�mN�:��9��X��B"
z�pfdtؗ��M�x��`2,�F� W�Υ;�r��dxfM��v�l� ���Ѿ��;�2Y�~�B����&��NS"���:�|y�s���'{�Q��y��Ϡ����Hj�X7WЅ����˔���`��˃I������f��c�XZճ��_t��aM�C�1���o���6T��O��7��ӰE|Hu��М�|���Q��[�mP�1*�"�~��c��;@�^Pp�v��`�Ό�Dk�_^��"I�>N���������(ڻ��Y��98Cٔ\�8L6�k�A�E��̂��a��;�%08�ɻ��E�2�,�W�xi�3|�vi.m侫m_&�Սhx�9����D2i|��\~U��g����n� F����߸�B33{1����w9�N(M�v�9��$(5I����F�˄Z\h~�2��n�Ӵ(����7�V�7�lbaY���� ���4�4�!˖���=o�#�����w�Q|S�;jCӦ�/�nVC����ݳ��a��s!aC���P���܂	�pؠ�xB}��e�m
���8O��֑��`y�CzD��	�"�(O��q�Ƚe*����SVH���c�Ce.�����U�\�A��)�a�#��k�M����6�r�B�%Hq��#�*X �p]�Yo�I��ח��U\识�]S�AeFoMO{qDD\UXp�H.N�z�GM����~�@o��{����1W�)e�?
�ܘI�M/�]P�Dl��Ē�$@��(j-!��a��^�ʨ_Q�����׽�
�K}4JJo�F-�F8^�V�s	w#qR��u�m�يv��\;k��o����w���"�4*qNj0��a.9�=/ "K�S"�Qt��Sήoמ��q�9��:�ʲz���7��#��'	��Wa�ZO<k�u��j�v�y�2�ON�3�����
��}b'9mX.t���^�讬}���)K�;H�+�ЖN�Mg =.���D�?>����&@	-��)�8!�|!�P�0�|�	��#����ј!y���i�ul��D9\�Ke*���[O�=;/�jK��j}��W�A?�WL��O�}�n�5vN��Uc^D����_}E�>�Ï:h�},�O��se��!/�|t+��gMo�>�++<QS��)�c�ȅz����y%A��*�VLK�X���)�"E)���ȿ^H�8�s���j Չ���
�W<��2��sz�������z�����������x�F{$f;cX�íP��l������e�fka?��*V�W7��
<���@~�D0������ɾ��oV<�W4���2d$g��6��7ۦ��K	��@N|w�C��+'￫��O�fc"�U��Կ��C�{� Є�n-�_����I�]��A/j��ݘ�Z�2!5�O!��e��$�6+<�u(�#������@�,�lk��WfJ����YHL+�!�ɳVN���~�#͡ٹ���p[J��b��R�R�u�1�S��G�E��!��v�M�4�DM�Q�l�O}�k�qP7v̉!1�H4��=ǒ��xjOP�*�=e��iӐ�(�.?7G+B��ɹ�2��Jt������U�8GtX�8ߎ�Ep�Bt{�]vw\[,�Oz��zy�W���O�q=�P�a�c�W)���(�ض2M�o�?��mS�)f��)��Ѓ�V����rQ���˱t}tg
�r ��gu�/<�_ ���=����,Y�^a�]�U��lOG�e�v|�XD��%�;�
�ɭ5 ���ӡ��,���$�n� ���dP�F�Mi*��M�je�wR��0�}^���c/4�r�.b#�/.'�`h�R
p�n�y��G���[)���EU~?�%�
�c$��e_��J��C��i��j�kl椟�z���g��<�͋�E�貛lO8�,���ŧ\�?t+��=3
�:ҴC��[���ca���*Zx4#��N��<C<9[�~u��1on�1�-
j_O�V�lۓ�]ؓt�r:8�G��R���L��� �ք A�"�~��F3���=o�ڄ��� 4��i�s�Ck�R�+�����mޣ��q�����T<d����p�F�7���W$@�z�q(%G�S�-���P�?:z�����	l���RM����M��K���"3Ьp��
V�L��'~D L���tT�3rlw�g���IKQ�K�~AY^7�V����WPl����爮s�类��JI2��"��ny�ȳl�`�|v���%F�zi]rq	�0&����g�0}��Yb=NB;:�[���.��>��_���cy�<���{�fPD�Gjn!���.���+ܬֻ��ӊ�D�-�#�Xc��ǕSu�F��_�r���BO4N�kbj�p����A�OndI��n~�k��]�Ԫ�"lv�KNGp��ɔ���VҬ��n1���yŲ�E��q��ۍ����À� yC���|�>s:�|ACp�[P�j�ӳ����JгɎ�[#���Mȯ{��7i6`꾸*�����ˆGI%&��r�[;�[���ο�Ga���S���S`\h$6�  
�l"b�k�P������KS�x�ʋ��R��7彭-r��"Ɂ��Ҭ�x��	8��F������.\1�E�ne~���R�j�X�V�γ߱'2�P��A����r��j��_D�2-B�X/~�E�b�ѕ�n�KE�6��;ٙ%ƒ�*Q[x=�^��hE��k-�d
