��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY[U4\}�(`	�5�p�n�b�b'�+�J\Q���bV<yҴ+�a��!�y���U��_1A�4�Z�'�:&ۣ�s��C�o��no߯��/KtAU�j�2J��"^J:3SHD��2 3�{����6,ud��h.���.��ء,�tB�=I��n��� �^��Sj��p���K���pҩt>����A	�T]�~�a�3�qu�Ac�t�]�b�<����f�S��6�bK�P|_��!	��&�_%$
��s0e� jG+��5	�iA>�-���j�Cuh3ےy��؃e^y�o��|�j��G��é������wjV2�0�}p�F��E���$ּ�'Ar�Z�b���K�w��?OiJb\e#�h�!+����qG��txu�^6՟��_�S#�ǧ�����9V�5	��>FC��^~�.���7�-�5T�8�z7P"�m�h ��S3)��6��@~]h������sI>Q�r��}�
�n���潡���`���%��- p�N��>��k���"C띖W�-Q�Qr���#�~i�G�5k����(r�[���m����s+V��e&��3���ݤ�� +��4[Vx�iv�GMi�9�P^e=pE�:A�m2���G�<y���1�N|^/V�x;�-n&�zs��l��*�� .|���W�F�6�EZn �to�;14S����g��1:	�X���8�|�	��!�9����5 ��Ӻ�\V�N� &Jx��k���)��1��Lπ��m{ԛLz��˨��TI�^�����E�-hO ��b-�:f�M���{^ư#5�t��M\�YU�:8�[�CqZ:AF)�3���7�Q� �Df�
K��k}
%�p98P�XTV���1���d��<p>U_Y���	HC������~�LL����g����J�%
R�'�O<�3���ą-`��Ҵ��7`i���т��j5 ��:�f,�c��^D	����F! �Z���Xƌw�1��a��ce˼���u��I���z?�,R���D���9�$|l���ܯh���fk�ڙ��yX[��I>}�Vn7��{~��Ž}����B�T��+�*�����W�Nٻ
̾�Sl���	9V2\{���K����s�(:p��\��I��ק�
�g�����Nzyj3GY��q�&���A��V>��\;����� �r�a�[a������VaZ~8�1X�(���0F��۴\��&4rx��ie��z�����)g��"??W�c����Efp��0 8�j�Þ�1�����KWB�����8P��c6�P����o�<fq%�Vq�:dm3e@���=����K��SD���)^�	q[�N���ZIΆ����ъV��`�A�Ө)7>I�}
JA�5�jX�"���C��&�}�6��������HQ�zBPa���R-(�ԋ�,��j�E�L��P!��	�� R�o2�{ܻ�����בqU�2� L���ȥl2��`Ā�iQ��4k\����o����B��.�fq,��rDf���#@�K���l���G����?��+A ��lR�O��ύj�'��F�?�1�û�S�8�zR��ūT��c�@"[�/k$s/�k�c��p�6�ˎu�W5P���r���[-?}y�4������
}�~�}P������#&c��\�rU�`��m��&"��.�Z�e4xL�*޹}OA��L�l����%:ط��&?Vt%�,��J�Ɉ�R�zW�����t����!�:t��	 �rP�M�ž�,侊�p�eA�T0M�P\�nJ>Y����~�$�0�]�]�-����n��_?�D���>���V.9E&�����L^fv~	�zA�� �~�����y�L�&=aGw;u:�Ŵ�k��#�V�A�������.�ߺ �)X�SH\�gMY�`��F��gK�q��@�@!�_�آ���s��O���ۤ6�^�Fnw=����2��]��Eavd|�o�o���j�(B���>;ٲ�"	1�aM#Q�,k�a����z�9�i�s�+V����(Pl����~d�<C��	nA!�C�1Tw,N����b�b�����-�Բ��e;�~���|~����6`��� 0��?�+YF1��Q�n!
�6T����O�P�96��	4�
����cL���l��qn(F
�t�zW �?ٞ�y��̤{E���|`���@���`oFa=� �:�B��,�xZp	��;ƕC?�I��Fuc)>>��ߓT!;��]l���.!�*.p6�LL:Pv/�}���,��s�"�6�/r��\��:r[�]��Ȉ0O�����jz�@��sy�xb
�O�� &^20��}��+\W*�s�ÀY��=�a{��גHcko3���&�M�,�&���A�:���͸�<}��I:1� �:Wc�}�R���l��n �HAWZw�f��nڳw�k��� �������nm�+>}Ãk�}}�t���Y������󮸛H�>?��\S 3���¨���K�
���������H�Rz�D��k����� ��\	�L�K��_#���X�	�D��w�F�E
�m���i���}o�a��*Kp�e�&n;�t> �S9�a@�&O�S K�,��*�� ���X��	�CК���c�ݛ|�t��Z �����.������������=��a�gI������䡒��~�m��2��b�w�[a̛��I�4�;]�˄P�˔��׸2������<����Y���Hn6�B*�[H�)2L\���?�"C���50�����Q���-(������]�	�%���(J̭H\w�<�]� �>}sD�����I���8�N>��r/_��U�}1�@�~�n`+yDL�P�g����Y��JU��Ys�g=���	TL�)������� Wé d�ȗub��'�WJ|�Dr�m�?��<��deޛY�{���)� �0_�_g�ݵapdy@E'�Dc�\a!s���p�_�&�Zų�[����q~�тU4�[17�m� ���������^��GJ�]���$�X�.L���9�0��(g��C��z`��֕�����ܼ�B��(�
|h����X[���>���Ч4T����%�z<#v��KaE
sl?�;������%�V���,`.�$��l����A�y�!g�%i��U\c;FN5����(�o����f{���5o�˲J�����1���?�'Ä
�v>W����D��G�����C.h�9g��ґ�՝)�U�Gb�O��!���g+��[]��,'́ETL��T���1nK��y>�Zm]Y��r����],J����������ũ�2VkM���JCtyO��������c��]��ЬػE!��������{[��J��m*�%a�]��#o�HB��A��;�F�n�<���%HFT"Ӥ{��	k�D~�1L�Lsuޘ�6�J������x�ۃ��b�p	��e���C��{)	��-���𒅮�N.m_&D.���6�� �V\  ��vB��N�e���˥�E�
�'�㡤�m���Ԕ�M\Ͽo+b����^	�=6�4�x�� ���@8>��LZ,�@$�`׉Mf���dA�����mT]=���Z��Ú:�Tx�9R-��}hd��]��SJ�.Ł�&���e�=�-#���;D���0��1�4����읱F��T��ZI!�T�rm`��1GfE�fb���Z��8�:�cD9'|��iƇ�=j ~��y3���NL���/�����3��Ӎ��p�X~g��A��5B��| �q;؍��,�i=�2��uC�j�f�	Y��	{:|)f� �"<W�"� �?�����I[�xz����XG��}�c�N
�Q�dM�!	����*�Ƚ�άH�Ӓ���f#�3���Ivw�;M�bB8�@��0�\Y���k1�؜�2i���t�2옕�|�H���| �U��Y����q�K*z#���Y�ׇ4�����H������<g�/�}гz���D��(;���Vt�7y�\���W���:R�z�H���������$1x�H�l�z�%��0�~�) �O�dqg����y@�"���ӓ�>����U��b�Z��j���S��=6|#��yF�m���3����0p�j����W��+��P�)�-?����ܾ�#+�E�}1����y�2�9B&3�&�epa+�I���#��ŀ��Z	��/ ��)ٛt�d��a�mS��3L^V��@A��S�?�-%)���Ļf���U�\v�$sF}@���<	��"���q���I�TcI��k��ݮ��C�9�	)��u���Ǭe��E�CKhk�m&@�U�+T�.貄u���m���	�(=H�J��]�P�p�xM@�dXϥ�u/� ���Rڼ�p�b/%ZP7�y�����e�}�,sUwmg��UF��Xs~�siB�U��V�
�Qh�gxG`��z<�4�j$X*���#�!��W)1���*h���k�N�Cg���V����ۅꬤ�|9�*�J����Q�rk���C�j�U�
��vN&�y%
 -l�"�~C~�T��?��w���Lscrـ/U.�4VP��f@���[��E���(��+r�a�\��n8߀�B��i���Nq8ʓ|$WX>��e�-�4ѵ�tY�d��h�[��n�����g
9�x�k�ź��z'H�4Q�"F�[t��ٌ��]u�����?\�� !ؤ��4�*H]�l�����t���=Կ����a������0\@��q�c��<�w�oL���9�if�Y����	v�c��MX��h���wư4O�7q��Y����P ��{��x�\8�;^�^���nYf,B{�0�c�f�:�~�r�Z?Ϝ2��迎�֗��!S�j��?����]/����C`�	mj�^�':k
('Ofdq}�Yڀ!���i��fO�1�� �Ȋ����/�QOY��sc=S�L��Rs�,F�O��'��� 2���y�~횶5�Ͱ�0�?�vh}Nڏ)ؾ}��op�x��u��5����7�+���/1�;��{8��p��x�;���M��n�Oo�?i�����x]�_����X{��ɻy3�Y�� ��yi�Vd�U"��f�6��3�U�<��?;�q��ٺD�4rZS���	q)<쏷�zy�񯢷@�b�I��Z>�3����j��v���][*Έ�ne�� j���L@��3�;'�j[��h�p�O�b�c|����D�ٛؽ�G�|2_U��TCۡ���׳�"2Z5��Ńś6u�z����<��V��H�����^��#x�ͯ��,�e�+(�gzΊ7����6������|HpT��G0/�{J�nn��K��0�)�|�$�]�z��i�ˌ�3#�j�����Pa���Dk-��1���h/�^؏�B���*kVOZ��<��F��>j%��h������o���Q}�Q`�q�g��\��E<�?vrp�M���׀�CN:h�E�4j�t3uޞz�Rk*'W��.v2��V�g�7,y���q����t�Ꝍj�:�7|��
m��G���=,��Q0r�톸R1�`
P�ȋ�0'j���K;-[��ˍ����k�DΤ�|R����'�P%��g��7��6�{��%�Jՠ��>{y��	�f���	H��'ͽ/XKv��?�ux7<����*�{��F�0��4Ž�g
U�Ւ����νX�OF��5M�8��?��A���7D�o�BÆ:�ٗ��)�2CdkOo�f�f@;��HYK��	�=	�E06�]"���ex�r2"*̊�j�#��g@���%��µ9؟�������懩tHv���h'L�>����%YD�A��%�i.��t�P}�e��a9�Zs�v��0g��	�=�_K� ��o6�CL4Kƃ�	�_�0	�l3VEU�,RBp�X��(X]$��T*xS�Y0yu�c������q9W2xVF]�}t<c���l{�_�1�w�s��Gzp/0�,sW<�'�Kgn��>2Do�}i��R
���/��J�/���G��7B^�ma�G�P�yk���;�e,Ѥ}X꟢���E6Y;�9!�9�h���곬��w'���T�E���ւq�h�n�6�􎒁?_7��\k�E@-o��VXo�������萜��\���xekq/Fp���M�b��c>�d��x !�*�K\�w)�G����o#�\-�4�(�u�I���c�ދ�Rd�h�'m'�0.\�������I�ަ�ǃ��\%��>܄�`��	���\2��i��VB;+Tk��v��m ;!�y��v�m��� +���D@��gB�4�Yn���D��8Yƶ�X����a��[��=����/M������k)EsME�ז[���J�M	!����j�#݀��ʻ��9p���=�1�������"d'%���˜�u%~�`0�x�%M��x���;�ʹ��>-\BX*e�	7��x���m�PN���BN k@5�h�d����c5l"���Ď�����Ij��e篲�Fm*:�W��(��Q��|��������OۡI@����5��/(�(G��=@� �1�g�,�쌟�YU�o��
�%�h�\�����*�ִ��4�܅I�t�Nt�qHP�	B�>u��h������c�6�Ö�T�l-�_�dsl�1�[s�-���z�Fv�c�I.�@��|�2|������3��������:�4�˛�ݵ)6�Em]xi{�y��X����V���	��2��fe����4�l�I����~�h��h���������l��ϽC��1g+���v��م��pP#��$��F�&����V�<Jw��숿�J