��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VYjf�>ρ�f �r�º�-"�|���k3�	��DέMy㿠"e}��oS��kc�'f��v��0;zt�+�_�.2r�#K�%�yE�����[Ֆ����2�����7��E��<�!�`R�kut�����i����d-UZj���ч�(�8����|xTH�	��!�ַ��z1l�s1���@�En-�>�~���$��W	�v��Z�~�q=g29B.!�(����n@�D"ݿ9��@�1g�D���j�vW��^}&{w)��<u{#ApW?I�3m�)9��<�ڱ�-�ɹj�ߡ�e�x�Q��i�՜���9�{�\�����AAS5=�{�;\Z��y�&k�~���ݟ3��$@��M�4ֽ�������8�P}��B�/ND�D�B�q1��T�M��T\��O�<4�pP����frDam��!��$���W���_��g���$�!������*�zŶ4՟4Q(%hǉS��+��ڹ+dPW�[å?�7n� Z��t��G�e����"��/����q��S�"��Nh���ˡ{����\:.��5�|5�
�!����L�r�%, ��~���W�˂�/�k��O�Yy�O���l<X4è�>M� �����ju��{��y��ز��� d�km�w�k㩴� �!�>žd��:��kW���M����;]���d&����:M�f�!w�U��qױ�f�F\�K���B�dȊ���"_�k+ �jl]X6���h����^�87y:$?�����!���_��4�4������ԧ�gK��N�^�Q�.;����e��0i�.�;��Y.����Lƞ�E�U���#�;��M���vb�9;���1p��9&�>+/�	���z�Y5SȾ�T�pܧWY+�S�p�=�y�N��L��$��]2�Y�i���9��*��Ҵ�(W�i��?=�	�^���N�k̸I�E�W,ɚ���v�zs�j|G}Babګk�#��5mO5� R�dX��@ܕ���+P�1��G��8Mn�}
�>����I�x#s����zЂ���zA�x{	c���$�J4���{&�wR�Loqn�{C�8նs���!]DZh��z��<�j�j����r��ڇ��������n�i��� 4>���h��	"�0��7�;�`ct��u�h��M�Ղ��KXq��j�w����i��[5l��^������L��_���.��+T+�A����O�Ad"��Na�z�J�5�4��%*e�����N7�P�j�V�%{�X-�D�Y3�&��\x7�Ny��~D9�ob�.�\(E(PYL;�Jj���X��2-�R�a�`罧���h�'5��`C��`VA#Q��2�>Xb�<�E�^Y��۟��5��r�X����N�ɵ��$����4��0
�P7�j���7�.�1�Ixz�)�Nc��� ߯�f��T�U��1��·7~�v�H�:���'dг|��װ<#e%Q*�M�(�!+�YT)��uנ�
�ҳI��ލ�ΟX��	z��LNlS	�Ň��V������B�6�"�x	�̥�W����d�^�m�7��ҥ�%�יu�;�/i8���f3X�Љn�,��¼Nc�d�¥~���tJ��O�Iqe&Zo%͍N�ó+Q����i�on4��n1�����q���{�	��I�I;`���+*���ܲ���5C��9�ۤsQ�V֚偱�l�8.�Q��!F��ͮ�Jα�`�������á�obM$��y0f$G"������>��O/-�T}p����.�@)��`�O��]���^"�D�%0�,�����L
�/��3FMb��kj��1"c<�J�|^=�N���I6w�2�0����iO̽r[c�
��0k���V���\�����b��y��vP��(z5T��˺��f
'����R	<k�k���ⱪ�"r�ժ����՜*.��V �,��T� $�#�~��@1�������UP_�^a�ys)qr�����o�J�v���GP�B����tB-�y`#��Z�a@h-8@^y�@�9�KF$������Vi�*~��^r�f$*o���o�j_CPk�!��"��Ѐ��fP��qK����"��*��:n2�Ni0p�K�����V`��7yy��MZ%��(�г5���qs;rrg{�^�@^D~D��^y#3�o��t�&j�>���0���[�H���7ˮ���(�2�����䩕����� =�ͦ�(eG&�я�=:>�@�E1��^�p�C�X"D�&�/E8��j�K�̸p�Kc����O2��>$.S�t�����2���4���S1a&��t7�_cXE��An-���M���^=8q(�4���x~VZ��K��#���@�dy�.��M�㔌��w-�ɀ�"9
���r�a�ǻ(B�Ghr�1v8�q����=�^�<gկ}���Z���P���P�LFж,edY#<�搯���X�KniCbQf�{�^���&��#�};�G}e�/�|�t� 0�.6,�K�$���,
W�G�:���3�5�Ļ����K����v������c��#M�W��kasb�[���NF��~�3�<%z*X�W��3E��Y3Q�w?j����&�j���l	�{-w��ø�5�.Š�F����u�m��	4��`M��ڤ��S�)9�wa����r5s/�&�z��mVY�:ls�{!_v����~�X���t��5�:	Zz�Oh� �K�hB:$�򋪵��!�1}ʏb���$n��ip��d)J�.Q������[�ї���~�iĤ?�)t�m����q)�fC�o���01�x�����,�R��K{�tq�Q3f@���n�!��W����O6�s���d�׶V;��p��O</����Sp��bp|l�A�x���Dj�7;B�Tg� 	$������=��Bf�hȄ�Aw�x������gТĝ�}f@ �����Ӊ3��hke}�I~ԛ"혘�[�f��.��S ԁʸYP�v����.lw�)+h�~���"MCn9�s�r-��Q���̛�GS;��1��q��n|}�t�?��T�MO+ոk���h��ײ�z��%�(0F��ꩺ!V�yv5\6�;�I�ݡ fp��h|p(�#�ӫ�l�\j�������#vK0���h��Y����K��<_�� u
�#%����j�P��=%�CM:GC
�gz S	M��Ɒ��F�l-�٦��47f�s�� �d��o�E�ߴp[�"�q�G��Xu�2g~�R%XQ<N����0����gF���)hFH8�xY���ģ���*<� �^�M�/9��JI	�aap�JNt^2&1��Vׇ����АeVg�����n�� x!t
7���߮ӈ�v1t�)�N�)1q|3$�p����Sf��L;��*}���x���N:<�^���N��:�,���%aڣ����|H���;2�ׁJ��& ���˧٠�L%�y>�7>�
�&��������M�z�uu�	 I������ "�+/5��Xɋu5���\�#�������5[2>�BK���HJm�@���Z�l��YDtm�2���� �~��G֖ M:��	���mFT��/�`��n�v��t%6z_��9���~�@p���+^��(���H�Mi�/��E��Bd�(d�<��&	��9��8~�W�&����^�i`�:˓93�ôF:�$�[ˀt����B�	S�_ɏP�Éщ��ĩ�-%HJ*�����,)�ҵ^�۴,c��hP�V�� �aL�Νt��4�p�6'��Zvq�ؤ	���ڑJ+�@>����Ɣ��k.V��$��w&QR$r*?2)���60�?���x��ϑ��#�G�G	��i_�)���;RM)0@������7�Ȓ	N�B��E�4wU�ce��Bl���%���٦~�5[�Rz�Z�`J��I`@�:�gH%��%��U��]_;	�It�;�J!H�Fl+炒&.��2��s�G�l�+�qS� -��ɜO�<�I.`)����лdY�EX���R95�,�T�^G�����=cM��J���w͆\��׻�4�^�2-�!��R�>ߗF���zE�r�zl)A.���_?2�lXE���9��Q�����h� kG0�.U�\/ձ+:��=R�J��_ѬOO���7Zy�t��e���Su������Hc ��|���r�λ�=�����Ι��l�	���>э�{m�ӁW���	�7��B��d�����O�
�p��	])���o���JY�wa���9$L�r���<����z�+[lLzɸ����G<�t�\���-d��^~$���$�Y^n�&���-�k�b1A������+�y1��-`mꅿ�^���=��j��c8;�	a��,楬�B�~�<�XI=\���(�j��	J�)ѓ�~�{�Y���p�
C��b5��/I��t��V�M�OdJ��h��ԡ2C)��ݥ[��B��]�����782�^�z�+A�I����M����E�]:��ꏑ@b��Za�G�R)���L���ʧu�gm�d]�� �h�"O/1����!Y�iBO�k����G̍ho��|ڨ�y�A��j8 ��{�dIoE�"ǄP�����{s���1��w�􌓽�~�1���M��WwR�U�j"�μ�Q0ߗ�s��k���Da�W!*�K� ��4P���GT�)�w�d�Ȣn�F߬?W^���>Gu��Ѳ^����gE��r�4=6�̧8݀kf��H�6�j��)B��qn�	`�>����;���	���?����P��"�r\�FE�-=�L���iߑ�i]�Ų��Y5~<9g}�B�9�͔.1�DD�V�,�1C��~d���a�d���ߋ�<��0hG�����<���:%�7P*g��,���^�������<(��?��n���P�#�8=���,�#�o�vB�ĺ��r�� ���N��R��r���2]�;����a��Ti
v�u�}���a�w!�?�і�?{R>T�b<�F�n/y3.�|������-4o9=7|":~@i���X�]o�3=���Q(6P�hp����ą@��`>�>�E#j��!�� ��fH\�a�3�n.�g��QnB��.=�u=�K�a��lV��2���[ӹ_�&�q~M��9�k0M��VC� _ӳ��gQ���a^>��,���(�:I�@42�i����|�P`�Î,)p�g��w�o(&����Z�ĩ*~�l���z�8v�.}�T�cg1�K���`|�x��6����Q�~S¹����!6��?&��x�Z�b�l3��,�(w�v���~�����ƞ���o���չ���z���o^K�m�Xݎ�N�8��M�י3��S��qblc	�*�0�g��9�a�>cn4��Y��d�l-�+��X(�fq����Ϋ'� F��@N�J�G��2�2���b�A%-��hb��H��}&2�_ߧ�F-��VԈ �Gy'd�oa4ۆ�	�nzE�ܾ|�7m��C+J�vU�Rn�����բ�1��Β�	�bQ��^DcAԭ��/�<R~;6��4�F�,Mڂf�i2��S�X���O�4�4��|��83�-� ��˗$�����Ģ��Y��ڱ1�:k�4@��0cEq�s���1���jSD�aS�.��܅2�����8>�N�A���(�v���E����'nܗȨA�U�H������G^j�j���݄�\�����Q�t�Ӕ�?JO�Zf�R.W�N��gY:7�Ɔ���w}/bE]����?��w�3e�9L܌'\d�)u�
U\r�\����e$:kG��4k��������V��$�� �\a���(�3��}-�%$���ܯ�����>���U IN��������%�m������>�yi`!�2����]͏��+%s�r7�EXP���X�~�*X{��-���"�БVu)@`$���H�FJ,<׉9��4�G�˯2/�8����u��R�V!�*�D	�J����k�y�\�LD�'����E܉������PqY������Dc<�wh���䲈���x�K]�Ռ��}���v�Ԙ&1,�� ���ϲ�0A���@�MG��b���EpT8�ߨ:Cb��
S�Q���\�[�7U�Rl����
��N��sg}��H`��Q��N�d��P���	����O��i���l�E����{�BG�����L�,3�g���k�I�ʭ��##P�d"� AK|�0/Cݰ&�u��~t�n7*N���W`��6�,�p�����lOֻ`��#_7������5ٿ�I���4I�x�_�KP����E�H��J�U��_��.T��+s��a;T!4]d�q���'�]�o0������T/�j�5�Ɓ�l󒶪�a\�w���*$���_|y�wK���?�jr����`O�Û�2�y׸�5��q�+M0+z���W4b�iQ�zd]�_���#�[�Р��,���Z� 7�V��.qZ�$$��F@�^9�K	^z�?`��d@T���!��@;\���zH�w���p�@D�2V��)���g��2y�X�X�n�·��QC�c�u���>'T��]�l�ޞ69�>����M�w(�i���tX�Ap>����I3��	�b�T%�<�n�`�Q	|�'-��s�"�g���H�ǯ���W�wQH����U��U��,��Z(Jyyr�D_��g2�<�f-�Q�R�P�砭|��k߰�Ƅ� 1 �i���&�[�lN�}�Ӏ|�����a��^��[�b\�Ϛ����m=u�W��H�>쉢K���I�L�Zo���+���^�*`%O�46��.�!x�qX���V�]��(�e�6�N0�LU)Ι-N�![(��ʩ��h���xHý��E0�(}�Z��X��~[�j��c��Q��p-�&��{OK��̎(��a��W��͢�Q��t5[b't1�	Y�m��zu�y�y.�@����.2 ��oz/V���H��nT�e��2Ov��iǃ�@���	��e�ǇJ�O�Щ��q�i�t��	�z�#���z[D �A\���~K��2;�6�,RX�XV���VP�ۯ��_�jY3�+��5cӟ���n��*�3����.���oXbR�E�KbxQ	'|a_�, D�ᓆ0���`�*���^��-�Y5t�ˇr&f��w*Z[�8�� �]�S�w�1�b@_��Q�x�R{j��8���:�i�>�j���,y4���'+�E��88��w�U\�ry㩪R��%hR��q�ȫ&o�@�+ꒊG���w����e��vhQR��{�.�!�����S�~����R�:X���<�[r-��=�|W�=��h*��U�k�t����K�՚��&%r����8t;J�����<����u�5e�g�v�r�R@�3u	��b ��|�)$�dbb-����Bӫa*��vF�ǅ�X��/�����b���e�G��^���H�(y�
Edl����#�A�]c�]�)*�eA�ǫ,>�Hy�:�j��d��	������ �^������XS�	���f�F:Rז��*sbR�t�#<���PK5���d�ǆ�Yl�ᢘ�� �_��O�
�^ *n�=u��9��0�{2��uC�0M�)�QEE�.� E�	2��z3�ty�e}4�ΩGZ�4��� �p/ 9ctS���v>�6�I�S�(��CRs�}�ܤ����E�*��2/��
0�斎��e��{6O2�%7V�����g���e�.���޺$_�(i�1*��Z��N�F�Ӭ���R"Jf�?�<���t�oY3(���%��쟓n���b�'��It��{������M��[2��b�}c,Tdg��$U��Ӱ����?q��0�M��%�e�m.
�h��97d����砈?Ө;܇)f7��I��v7Fٛ��5�mK�����,wf��̽pr��4T�/��Up��>��?f���������}�ԭ�����wϣ<}���Jcٻ��R�.Q��t��#j�c(6�����Mrd���t��w�,��9���.O�w�7���LY'��>1A+�a��5G<�D4���^��s�3-a�͉���@��._HU4�S��"����;S��]0��7T�7Z�ҏ��9fꋰ	a�~d�	���
KβƂ�hO�2�d7@�v5=�h��Y{Q�a�ń�kq����"�A}�����}-���oтO;ό�Gz!��mq�:o��S*z�rF7Kt*4.��5KnѯH	0N�v;h�aHrX�!����of>]s�#E��i�K;boT�e�9��7�A�%F.�bH��9�J҄W����i���������6�h�<nm{Q�7:�.��W�����y��p
Ú05���
2D7��0�{>c�������}�N�ZE�cB���̓(���Y�d�>ʞ��s*���M)�l5�O�b�4P#�_+�9SP�w��L*�p���-��+�.���E�kU�?�A���*��}EU:�$l;��W	@�?���rE	W4n�f��H�H��o��k�M$#qo���!$R�	�6��� ���~��d�Ӈ0�{�{�]�ҝ��jz�w>���In��.u���D�Y�0t�v"q�`��޻�-�o���Ӥ��2`iQkG��)&VA׻��d�T�I����	�ּ<����NA�P��E�T&���Y{ �%�+"q;��ÛT���L���!Z�TR�	�G2xH�a^
)g3���A��:��;�FR+H���PMC�܀�{�wd���B�&�d�N!}ˠu���;���㾖ٔr��G�f�/d�B( *D�=�b�x�L���V3�8��njf�I �/)7�c&ڰnN�Q���ua�,�<&Z�b��F��BJ�hՕ|N�*�?B������G���0^)�^��)��Ȇ���%�ts�+��1u~��6g7��:�C�f�rDfxғ^^�ׁ�!�ꃊt��1F
6w�ĳt|̭�Y����%C�-{�����=�%���j����O�J��i��b����on�p�usi�����)����U�|�B�'��ە������]G�r��O�p�2ˡ���?!�ԓ��w�A�K����kd�jK���=v-��T��Y�ZX�^��[��<��[�Q@O�m.}f6��}َԵ�s��u�\e���2M'YPD�4z���
���X����sЍ?�?y�;9R
��AL��]V�ԯE�b8�%����prA��ž9�⛲�M�p��)��8дBl�au�#Axڡd�����A�n�3��\X�n����8��{OK�A#��m8?�2�(Qn�����p�r+*�� �s)ܾ)�M�W^����V�,on��şlfq%�0�^���	26ΎfB�~L{N�ՆV)Tc���d�A�kF�%c���2)�u�d��_n\2g�7T4"��j��X�,?���|Y��,JI�,'��	\���\���!c���R[A\��l���g�C肓���`�%D�E��k
b�G��ZvQ}��@I%�)�1�χ��yi�c^K��ya�[(��D�A��w,���;y���w78:y@ߝ�r�D���1�/����|�;��PV#]ēA���g�6<���Jy3:##�)Ү�e�3��]҈ѥV��o /��y�+V�������^��6`+D�x6	����e�:\�)�UY�@�T���N��Ɇ�[6�u��� h2�$X �{��l!N(��}-�� �/e��TZ�q�4���������s���I�j�z=�AM��.l]E��V��|����4�?)����6hx
���Y��˥��b���]@�p�aa�ahц:pH ���p�!>੖���uI�#��hL��>��Km;ՠUV�����>��z�Ml*wʽTo���!��Fn���3�eqE��x##(�&�Q��N!3�
XLJ����ɉ"3��68�{��X�W|�SV۽^��~O*=��SDE~����\��{1Zy��[���?�Ē,m��3�r���/�H�Yv�A����P�#�W'CY��[1[i�T�5 M��ܼu�dl\xQ�͗��Ӕ����-H<����@�c��y�>��H���^��b���C��7	�D�4���e��m��&s�p�N%��S�5
-��z
������΅=r$�;����=*D�I��&�R�7��сx����*id���Q��5r��,(`����O��9P�bZ�7<���m�����w���ƕ��4-M8�rTVϷ�8g�#�xV�2���<N���������
!zPj�B�g���GTZ���o�1��!�1����=��]bC.�e��{`A$z�d?��e!K�̨S�-z�U�g[¶�~����� 1�u�
OSgt�E���[N0�K�%�2��M��O� ��(j<�C�#0T�@�#��V��N���J��O��� : 0�Մ~v��As�+�<ɽ�b5�����d�zk	�-��(�?����,Tdp���p+}n����E�%�2��tP�5L��>�/낓,,��i:a�wK.9nr�B�cjr�u7�]|\
[c-�c��Z��
�qS�-0L�,р�JK�r�e����.Ǫ�T����VǄAb$~��:uz\e�����P�'5M ʢ����ZsR���qs�,��I�M������+`��}1��5��K����"�����x��U����=��\��l�t�-ǲ/qU�7tU��J���˭�#O��L�d��92�D^�=a���Q�q�0��׍#�L�u��="�Ѡq��zY�U�7�q����0��(��P���bF��O	{ۿ�菪���r�9�Q���uKRMZ�/$��s��y{x\�\�ES�w�*}��f/��\����	��y�-���=�G�k�Qm9qʄT����5��Ώ��`������
 ��u��#&��\Z���؂~�X�mP�L�����8C_��Dw ��*�����o���\֕��?7V�l�ى�cpAO �ڿF���_�\ύP��{�Iq$�~$�}�LK�;-��C #xs:v��n�Y�Q�֠�qgΩ����,�j_U$�՞�_a|�7f@�wYa��78���u��<a�LZ�1a5%Ea����,y�Q>����<^pq�q���,3�g
�Bof2�1k��K���%}���!����T�?R�Z����42{�F�g��� ��J@�_������Qh��B�mi��:�:��iC���zJ3-��@Ɋ/\�G֕�nW]�q�U�1�Δ�4�?2�+��={m�_[��r�^�c�[��
�e�A�eWݛ���*:,�WH���̫�t�8u*�yg����ʦ�A�G�|:��B�.ע#��^g�橦����Q���?+� 2G��:nd@�jgNz}�X����c.[�M�8��ȣ���1�$f����]fS�N�z�jEA�p�08ncqG^��#�h��+}��<�l85��婈�]��9g���Rkg�7�F6�c<*�=|19�$eb:\6���8��R.�����o�I�M��N������UD�`���]ן�x1�߿M]�O^����Q�l\�O�����$�|7cs���G��)	�0��ߟ��'a�hh�f7(���
)(�A^%7�j����<3Sd�F��߃��g������n�{΄�˼VL>�����ޅ������Z�7�(�C���<Ǵ�4��!�o�,�)~��I��R�#��S@x������\l�l�]e�逊���%<z��rw_�Y�~���#����(������=|���+��5D�O�
v�r2őT(�+US�y�4�Wekn92����x��=;X	��fJA���W7\��|��'�K���k�*�����3�t��Ia^�>�	�~�l6v�g=�y�P����m�]J7���U�����w%{�CxB�vV��'�z���R`�\Q[�g9(.+C�e+��/
�Iy-��lRkg��$�i�[N��Ƅc�غ-��3!UxOh�vuRޣS���^�=��z�QլO�dCR�`K��*����(�G6������_���/�G��k�����܉��ͽ�����K,JE���Oo�%�Z!v$���{������Y�	�B�Շu� _���%uSZ��'5��^�fs_�?@X�Z�<�n�[y�U��%
���'H�:]�Rට��eM�T:����t���.�<��8@S�Mر����Sk�liڝ�(�U~�䭟��S5�o�]��sj'Δ��&����&�nA �Tܖѿ_�io?�F�/���
�Qo��:��s�+����'��AX?dIzM�n�3[���;7�:��L� �����45
m7�a����k�֨��ؑ���EY��p���r c#;���_���P~W������ʅ�ZZ��\:��8E�c�t_�̎bTLv�,��(��2צ 1�	�����i�ㆮ^�S�>�|TҲ��`bd�i�t!�$K~h��6��V�w��Q/#��#�
�}�0x�:��@|B_���=�2(�'*��t��?�p�������%��fޒK�o��Ҳ��#����*�Bg`N��.�J��Ci����VBW	�R�;�D6>k��*+�\�˦����q��0�N"ЇՒ�=M�-0"s��#�F��tE�eE��`Sj��.���7�YD�õ@݆B�4%Q	^V)b\U��?�m�9$k+��Oܤ��% �B�����P�8 <���x1�nk���ԛ�����a���Q�X���WK9,I�m����?��U�*5X[�J�Ssi
L��Z��&��j�j�%���	��n��]e��#E��S����VΝ>��i�����G���s_Q�sӸ����Ɛ:�Ibn^+Ghi��������bcR>X�vlTڣEn��� �I���K�^04	�d�#�{�F�̅��S��c����浶wrq��K/$��9�OF����(/Ob��y�c���Mr�\R�J������t�����  K6;S�:��e�.�\6&I]@�[�&Z � ��jtK|�x�^gF��
e����Z+�~�ڌ���<��42���y`c
,���Ρ���9��������� �CX�B\��Y0DU��8�:.��n���pY;%
~.Ă����n����!;��y-�!�s������Y���2��w�>�Ե� +�|�-��3�S
���w�� ��\��T�f�2?苎�K>r��\ĈHkqw�6:�q�s�11H��߆�)��>6�!�c��$^ ��a�����j��Nq�C�}@he� �n�(*����v
���s� �]�w�>��I���j{䠝p�ˌ5쇠G#n�(�^@:���+:�����KC�Z��n�;���)ޡ�2������9(s,j�¡�?J ��/�oyR�D�jt�i�Ł>��ݍ����y���juH_�p�m5�� �R)֑�q4A?�a�p$mR@�慕��vrt�ґ/%�[���od��|Y�֤����+�Ǜ��T G�)m	|4X�wM�Ww�����|�P�5��%A[�o��4{������XZ�T����
���U����fC&�CEK��"g��kC�t�`�K'�/�{fK��{t?�gn��
@5���v)Ϋ쭜���3V׭�o(o�6��aG�F ��)Ӎ�(BB�rr^�)o��.3<z���l�!"�q#s:qH4��Rp�P���'ܣ(g���}��w�|�͟�r��1��9vb[�&C��ϢO~�;�?.1����lzEW���^�N���i�Lgp:��#]�]u�|lI�T�~���u���')Y@|�¿t�+]��T�����7�%�۠p�c+�K�Ϟ�G�=`zpQ��[��m?�)%��nu�!�ojS��`,Ũم����7��!���깰OGŻ��~(��J��N�3���[^�"�.�I����@�w�$��dϗ̾gk��-YЯ�'�"��6��߫�innp�2�����Fn���(� 4(����k15����m�Ge��pC f�~r�3�1�4
��3V� SP�k�<(].�Q��W)�J���NY�
j1�_|�z?�8�m$�Ǜ/1$��t�����p6	���'h�T�b��Y�����&[�u�h���Hޕ�w���i*m��n�p�3[�آ�����D���
-
˲��dP���~�g;	��~E��=�r�<�by�Pm5Hk��ͽu#\s�l��5��Ami��y2�P#��6�t�U"-�.���~�s>G[w�9�jK,��C�)�=��>O��Q���M@/��|�%�p��m�v}77�E��/4���ō��3���y��1���_:����v�"���c����:�����H�:�"/*E7��C�9C���_.�/Qb����u�F���{�^�|�G̅�$�Ct��N`����4*����JD{V��� ��c��y��<�h�i���7 ����Δ�Y ?��&�F��Ӕ��¨��}�S�^�Jʕ�k�l3���\.��/Ձq�lJP�rg��������Qe�J��g~+�o��� xUf0�{I9D����g����>�TB��X����A�����kB���g�;�s�y���=֯�O+X����˔��_-�>�X������X�UZ��z������B��8m�Y�02{2��w�P�oX��8uA�Ce�̒�Jz��!~����̩��mc�Ee�G\¨��Q�!��:_Yb{G�|�{:�����#��2�9Z��*�n��8��x5x^��"��ĉH����X�em�2:���`��^�:�>��*�*>���XO\+Q����h�'���ih�0�����[����U�����7���nu	�{[���d�Y���?���(�"��Y:p�D1�Kw�t� 	�����C�2cm7�2�����N���^:�_�=��v�'��i�C���I��r�8����;_�,�fE�ޔ�I�K�:�,1�A>��E�4���b9���)�6�6�\]���C|z��uo,��=!{Y�i�Y
�<�0����|D�LO��	P2_'����V?5A$D�e[�A:��ҍ�������S�-.�z���\�1���^�>�Wl��``���R�PV'Գ��H�	��ӂt�>4|A� Y
��nTI	�M�2�r�)��5~e�����2��������7�}����.�׋��#.�<pUΔ7�g����� �&��B������2#(�f_\�J��)�ڐ�h�m��At�q�n7���<Ҍn�VP@�l�� _���(�5�2bs�<y/�ƠL_�=�#�0��,}��g���|����T`��f���Α�3$���~��KikF{@����!���Tu���$����-}u���T����R=��>!jU�
��~@��ad`��x�.�i�h�����,A1[��T�Q�Jn�A��7ĪB�v�e�
Lj8����RsF��,#�Ao;vTW+g��q"��P��"�X��K �۹K��X�'O�^���V�m�R�^�7W�ˑ϶�'c�,&�9R�K����DZ�4��֚)��1w!<T���h�&n)��5��?�`y1](���J��)$?�]�!�W�K-t=��rJ�d=�!����H��R67����?���2:�qn�v�F�ٛ�Ť�4�wt��K���E�Y!��$��/$<;������s�M.���Yb���	�T�Sݿ�#��UA����l/efU~�"�F�^5Uf�
©uEG���
h�4�kY�0�5ȳh h�R�[�%t >�{
hb �/�]��2�v�y3A�~�!��AE�BE6l���Q�|I*e7R%#@��)�N������ӱ�*�Y�! ߍeY��"�Ar�x_�<1� %lA���bA6�����*]`&v��I?;I���:vtR�Ή��䍨����YM��}-��җ�h�rRך�U6y���?@��f-i����{2F�$�b�?S�5"��Yu������+� '�����9ڴ.���CI�ı�+�Ȧ"8����Mm�kKe��<PA����� �� �P�|ot�����o�I�=Y^�8�]�w[�n8R�ͳ�r� �%Q3�?B�FԌ1%��i.!�;�/W�i�ջ����O���>yw�dC+��v�O��Z�ux��_M�+ҳx�GjA�-Zf�_ib�EI髮�a�^��fƫ��+b��C@�}�I��SE��aJ4�ZtE��-U��?IU[r����X$�u�2i��EZd����y�T�ւٮ����ٍ$��$�L쉊lu��쥔��S.��v�������s��B�4�u19L�ʦ��ڡ�1�fb(��F�������@�)>y�غ�3�x�ɃF]c�Z�Cw�oٶ�x��|i \��M�R^�ɞ��L=W�GiV�U�M�>�%��J[D
�2P֊>���#��4�V�tǹSSj���.���E�	��0�Z;=�8��素1�hoEڲ�({ֈ����4�[S0��DU�"ẚ�)�M��藑�9��'O5 g��"�)�)�����7�IpY-ǇpNK_O��N��vYKP��~�N�� g������Z�'��X�����:3��K ������q�A����F�Ca���U͉MN��Z����Ό|�n7�s��ug�خ;�p�J�O"��8���pAegv"
R� �̬%E��W1AU��VhCͥ��A�q|�IZ�gHú��g�d�ĥ�g�#>��->꿍�zkHx��O��["� ��{�gc�Ĺ�d)���&�䟫$ECT8E��Y�R~/��2#���x\1��3�4Ct��Ui���vj�����D�وUځNA�P�y��=Lj�4��1ֻ����M�Vl��p����M���K�G2�z����4XG��&Ć��N�R�AY\�D��L@g�B+��S�:��H���)�C����U�SE��`Pk��J���>nO��<��y�̲��l�s-��H�Q��%�'6	���A��N��L<q`��3Vw5��<�P.�5�W�$!sr]��Mb�#4Q�LP?g��(�A8�S��S��ө���N��~��2م!����j���u-B� Ji��dB���(���r0�O���A�{9�Dif��-�ׯ��(�5k�T��D6��.Z�&3��-v�X��t�O��Q�U�B�t�$����^as`N�ts8a��\2F�»�Ys-}Ho�k���-<y)�z�?�(�=�9��[�Օ��櫛D�ˌ(��<�	�=~ai)(��'h�+;w���1�ʻ��U�'�>�*iS��<�����cH�o�ú^g��"C����Y���#����_qfnv��Ig����G��Yۈܼ����$���A*Y�R�o	uO���X{��t�WU!�����4B���=@O	��w�FTF��Zuw�$�{�D�	S�Fb������<T���,Z�}�o?S���5g�=M=�EQm0Y���|%�Е����K�)���E��Y�{���LX�f�5�[���ה��;�@��0"m/Q��Le���64�$۫�`{FdY��@Xd���D��*����Ad[��j݉&>�&4T�?��j�'���f%��S�?�R�E�O�u.�$#������W����B'��G�A���td���Y�\�!�4+� �}z>�p3JcSHk1�V><��"Y��`�0"� �,^��ɫg���MJ�Ao�+����P�P�q��&|ǆ�6�NՌ�(@~V��VcU������e�q�ˍ�6�T�,���v̍.6UU��7����1/����M�h�4:�u^Uł�;(%OCd`��=�$-�&���0�uʊ�a�i�#t��6��I����y�;s���
(�{���簢�*$3)�Q����5�.�������"�P1��*��2�7qU��Y0rAj��Na���U�m�*���yRbE+�x����ڰX���!]g���q��u�q|�B~��ͱO�D�9�)61�G�Մ��e*=U<��lE���^���q�]{���&��i�G��Fd=�� 3���N=/Ѥ�4x��@�_�BC6>ؿ�H;-#�s�G	4��Iz�w���cN3�J���#Z�Q�0��>�� Ci���g����[������ѧU�x眀�.L�G"_�����KC<�<�B��wN���&7�Q��c�Yś����lo��O�W��}�$�����-Z��� �U�@^��a*b�N��H#&m�9(I�s��d.P<Tv�_�o�q�L^�E�ܚ�ĪȂw ��ʬ~�6�������,��CPS��8u�$9��P�{,bb�!LJo��C����%��A��E!�7^(`�$x|��D����+SCX��w���Ӟ�z�PN��FDK����=Ц}2�X3T�2��+���@�J�uK������р�T��CI�x�rd}�I3.�uT[a����l�F�s��U�����uu1��O�Ԩk3 �U1� �H������\��MX$��`?7���2��ALC!�V����Ul�n�&��P�����/��pd�XzS��<�Rˠ0�e���߮��I�+v�FA	�W	1]�i����|��A�ő`��,s��U�D�/����V�Vᴨ�S�>	�V��$`bMe�0J�r.����8�{�3m�t��o+	K���|i���N����|܅]ňGcBy�ݕ�ts�@�U\�Y"v:�K7�ɰ�8����3� BE������G�}�������NRA�@Q�&�Ti�3H��T��NĻ�\�>c\RB������F�N��cq���3�g@u�����Ϸc���w��pVD;x��8��m�v�7\��_���\C�s���Ys���r�ӂx�"`�Ua���%lo�6;�\��Ǧ����"�fh�$:���hq����PI��	5������t���}�4"EH��ޙ8��AR��-���>��t�d�f�ݪ��cF��&-�[l&W+�Q:���k	z�M�0[^�m�3��D��O��Ǯ`�5\��B�M�R�,�)��Q!�-wB�OaE�v��0]���9�Ly�ث-�]@x_�N��/uʈcE1�Nr	�F��w9V:_�C��� �<�@ޭ7�ָ�p���aH���hB1#6R�_�e�&B�ٺ��AgR�\��޳19�}��� C ��:	�6_d�g�����P+�X@+ڧ���1�+�p����KgQ3مDY����`������{!�z���g",J�k���]�
�
/�s���qS:�I�堨'�%�����r��0_ؓэ��9#[�}��S?���"�r[���,������.rjÒ�3��-io{��Yh?�q�q	@�B�"n校up+�\�R;㳔�x���A����Oj�;Y�4j�Q�'�1���S(�2��F ��������@?���;�0�L te�B�I��N���@�ࡀ �Υ�c�d�(5�6$bH�v��c���Eۿ��^ph��?l kgh'K#������ȩ ��6�MR�����$Ȱn|�tƏ��,E��'̈�^A(l �Q5�?�g��|Wϩ��$AE�Wxl�`w� '�QPj;W������������$f�_Q����?~r�t�Ŀ�(gq��	{̳%e2�I��E2-�ȸ_�1<T�x�=EW��N���>�F<{�@P$ yH;������Glh����a^f����N\��RX��p���xSd�aVL˃^AEaQԏq��scg+QВ�W�l�%��
��O"e,�BOi�>�=H�@�@8Q��&A�?a��JU�����^��in�\�t�*�� �iѮ��M���2�]~�~.�\�k�����<�Fv:�i���{�ca����v��ҳRR=��/r(ڎ1O<�?+�{�E�?���n�@�?���(	��<�҃Y��B��P�:�M���A낡��1M�Pa��B�7 v���7�T2ڔ�kϬ�a����ޠ2�~>ӥO��T �k���"@_3������ ���Ђ�j��Y�oS��Ww�N�xA� m(���˒�����!�����C��;��.��b���GU�v�x���N��
�~���J}9�Z�t ڕt!a �s<$��l�aEW98$����JT��4d$2��H��i�ΰ�]7&F���Ύ'8�I��n�;`}��.�,���O���Dh��SAKRs(�^S|�/0S��"P.v�H������N5��Z	飠#n�p8S��^�]f��,Dd���]�lMA�t��D~A�a���#؈٢�4�GJ�;;��a�k�%aSi}����\��tnC�*a��Q��ۤny 9g�5���{ة�J��R��(ס�G� H�}E��(��F�X��/�����&a-�ڥ��"}'<����lPs�T�c��X�:�)�,6�Y��I��z��#',��c�T�"Gb���Q �kf.��:��J6��@w_1<��%]��im��w(Y��`�5#�h(X~k;�����NZ8��g�9�G�,����1B������-�~E8�/oN��Zݽ� .���(¡!�ɻ���Md�Y=X]��xan"b��mQ�5>��-��gT`.���f��<��Hѕ�>r��}w'A	���}tݵ�x��_}��/�B<�w^A��1��k[��M>��v�Jhk,�02�,��gc��rߐ��OL.XZ���5�c�BЂ�d�z�R�=r��;H��6~��kp��)��m�ɡ
Q���x����D�&��3�)b�bB)���8�54*��y.�M��vd���q���4��qW];����Ou�qe��4"&�DO�-Ӕ�\g����$`oL�d��`V鷂�#�F�������v�̓����E�kL���7T��<��^ϳ��
�����i�n>�w3*Y�����?������?�������:��I�iz�C�K�l⅏�j7��P z�㵂��45��P��]�@�i�;v��"����`F]k��;^#�k2߼�~����~�ɚ�k�8��1_������\�mn�fo��D,Is\:��/~I�]����/���M���׍U�qa�݊`xoY������ď�p�/��[�fe�=)��M�1�8��J7�
�v���k���%��*��2�CS��(�w�<Z��_Z�-��M�����B+{|y��PVl�1'_��2 �����:�W����P�U��ꮟ�%.Ӌ&�*����n�ac[v$#]�'�fS�����K�Z�|��=#�c��$�y밻���E5؅W����yPL�˽G��±���-����Hǈ_~�Y�h��������)E[4�ꆘ����,I�Xv���v�1'�d��§|6�=�}��r��E�}���\G�u������«{����/U����La.�]M6��X�Yj֍pP����Ӧ�LOQdU��y��O�ho�(��ҊN퍧�Z�i�$7��<������߬��)$�F��rz�6�D�q�?���B��w�^j.ҍ S�?�A�*���W6^�&X���+� @|�I����xFBᓪJDg�S������"o%����Wk�&�؁���U�n&M�\`�Lz:�)��9���ښ����W)��c�j�[�#�w�],o�,�J7W�x��u��)�քY9��.�tR���-T\�t��3&�:�$	���������s$ƣ�e��Rh�j��>s���0_�����K�h�M�	ȁ�-��DV�~�SE��
/}�-��bJ���u�a`�ԯ69��=����)���^�Ѻ[�'�,+�v��?m�v��ls�l�o��k�r ua��t�L��\{e�bل"*W��l����݃��V"�\�4�=�a����K�]��������!~��?�e}��?+[����a�dg�X�u�x�^�������#B�
�؛Iy����ne�\o�M I�GR�)��)͊'��9��۝��7dn�����c�.jM���l�ca>V;C��ҺV,�:�	����a2/��%<B~�a�D�|g%Y��0�:#��M�@X�f,�}ʼ�(�D�R߸+>�����-C�(f_��`�\v�ˈ���4�V�|+&MC�Y2Z	9.5M@��՜�9k����[1mP�����諽��h��Y4�����!�GC�eV:b��l~�s�ٵ	�U��?�}q��_	4j���`j�@�w��B�J:��el�%tዅ&�\)�/y]cT�=��h ��F�H��׫�t2R����˅���I"�Wp�B6����E��q�*������wik�6ɹ�*��o�QU�O���^��
�d�є�\�v�gx�=FM�w��fJ3�^�/H���Y�X�I�2��%ШT������q�Ri���E+���k���`1�i �qY�;�e�I��HMp�Gl �*�\��%�r"���-S\�7����/�����c��m;�Q5@�����Av��b14��r[s�=T͔���7��-�M3^�Q�q'g����qz��Y��7_�=�2��4�5�4t�P+�o�(*p��4Cl�� c�K�����I(�_��a�&�8��z|��f{PD��rZK}Su��A/n�b	��΁*;�|77�ż2�8��k��0���4���Pk�!2|������YY���:J���y��F�S�=H���.T���04��f����L8j��(��$���j��5x,3�Ν�'���7�����鳇�2+9�n`'[���ʤ�uf�H�������D>�E��Bo���5v�?��c�˝��L~����A ��@�s�(��ˈu����K{���s��.Ã���~�wa��,-Փr�YY����f�3,� ��fP��5�.���L������;���y%���3���v@�=ͤ�����f�)Ĝ�'�,j�f0�a׃2��¿��غ����iFl�!ڪ��qw[�����rn2?mNP�+8�B�\�!~�]�N��sYm��݄���nJ���3s;C"��k���Ӆ�;_ę��x�Ő�r@���ܗ�/G�)s6;�D��g8���Κ�9g%%kRfXHN�����$�Ć]��؊X\��A�Q�F�4�Ȝ��ҽ|%P��.���;�S�'��w�^�!��z�����W���
8_Ho^˼'r5gZ�� �:~9�Q�8L�U��(�P}��l i��������?U4�m���z�1W"$oDc~���~Q�l(�茇Nu�/�-�%lwf�'y�,�jz'��vl��%]1�~+�u�2ek0�m֮����R�<Z���Z�
��s�?�V>�r��XZú�Ķ>�p�}����}m���)���!��
�$|���L���D���:��f��#��m��`ш��֔��$�"�}�z��ᷗ\U�9�!���UO��F2s��_���8+�!AֆY�K�`7��B
�}���@j��P��>bN.�!��?���M�?٤N�#Q��:�4��6FKV�a ӷ8m��e)�(!�{oY�ԟs��	_A�y�|/D�G�(.�W�mp�G��cEa^�[yF�+ �v�л�����l!֩x�����T��4�ʈ]��f��Q��\���A�����h�����v�g��$��Z�Bxe�M ��Lm���x=oͪx��VO�\V�� n@�b� �=yvΤ�N����8�\�����M>������0}��\qzk�B��"� i���Y��3]�J�f#�TǴ�#���IBɚ�z+(�K���f��%��?�IJ��ZL9��# :��z!~�F}y�b���;�f\"5
Pv�_6`���W�Q��UJ�ƀ4�Ֆn�^�=�l<_����k�
���c{�2�X	S[�p[/��g}��p��oΞg���7Qr:����Tg_o����'��%Ѡ5��JZ	Y� �o�M�p��r�b|�-ȋB�A��u�\�`�I��^�H۷�tU�B�䉡�Y��/ g��[���^� ��Ȏ� ��)I�OժͺD���;r=���n 玨I~�@r��"�Qx��oA'N8�.��8�s�����}�p��ȕb�ymy��I�p�їvZ�	>ja��%��av[rT���X\�xD��=�)��;ܡ5���)T���~n����]�n�e�g$�?I���D�&�n�(�ȱ$�Ļ�r1J&3N!��
�i�䰒�J(��n�����4�d����k8>��/]zP�:��.��P��8k�e�`Z����x�H�DXü��ކ�#��?o-�O�[ ���q�/q��{�iˎ����;��]?���A.�����D䶋b\��G�XXӘ9 ?6Q��Z������էR�P)��9^bb�@�C@.�/X���A�����O_���W �X�Jp/�ֆ�
|c	m@���?8(ҁRfW�0Ϛ)h���X��OMa�,i�����	Qe��H��^0�P�\�� ��J�'�97���^1��[������ya��6�b���-p�6�J
bA�	��s�D �Γt.W�� n���	�z8�]�g���{���?&�Dd�$�����;�}���VW��6�׀�i��F{�su�p0����m�o���d�!AE5�s���(��	�6d��d9{���.�Q�a�'�Ͼq7���x�,���z��vC�ȣq��إl{���L���K��nҘ�/]��Ӳ�wq���m�Y*�	,� ���4a�`A��������dS���J��jh�s�HON5'�Oa=�/]5�	���&��x)�- _&?�s��ش`��n�w}��G�f�Q� M�)�x�}�9��|҆R����11�#�F$]Jѐ8�mMٞQc�L'Ҿ�����h��bf -�`@�좔l��{	>�R�~����x�q_���s9,_ZuO��G�y��$�H��@ ��a���11*.g̽6� cv��Tt!��~����h��N�kxm7�P��n��>;�*��b�G'��]	�,Q<�����<��*�~�n��2#��[�CJJ�J��f���H<��o���!A:�SE����H��lk�� ���K�|�\nޤ��6�2�ީ䲟f�?����m�5�f�0[t���Z��h8��l���2� ��V -��4nB�y�&���3�����	3D`WӘ�#N���3�����:
b�Btoj��������\��<�u�hi�g5����C	u����K�j����U0V�]�[��s+v�ւ\���ٔ=;�yU���>��T˽.Ŷۋ`�@���2�o'7	D�u�9 �&Q�ĵ"7,JM,��V@@ۧ���6��[G��l�$v;�T��Gd�'l[��L�坿!���TXR��=�������,��%f$�SbJ�kw����5Q��ӱu,��wAQ!�H��$Y�y�'3t�,8��ƗY��d@Ԩf?z�ur��u[���e׊Pu��b*����_�%���*���s����v�*	K�:�»򼰟z��ݣV�zJ�\����̻	�l{M�Z�)�P�.Df|*�Uxj����L���ʷ�9!��*��[f�Qc��TmJ˷�F�a,�E�(W ��9��ְ�3����N)�u*����wEge���������RR����6THvi7��Г��{,�%F��3=�_j�_z9C�iO"���f�A�I��P�2H��lz@�����,o�j�0�g꧓���q���YV~jXޖ��%�N�6�=��c�wey�I�(t�AJh�CZ�aE���6 �u�$a/.�О+K�į��i|��� S��w`%R?�	�Ɉ��%f���-χ�B�C�s˰�"�����0���;���~$�W���)6ZE������_#����鷳�Y�0�"|�'�$��b��6�OP���=v� m��$�N� �������UΆ�1��e��b���jɛ�i?�U��d�v������A<I�?ђ��i(�m�_��A�ݪ�Я[�g�O�hg��Y$!WXf��1Łި�Ag`�A]� P:���5c��0Ԥԡ��օ�&�=m�gw!4���i�Ć��Me�ApUΫ9���� �(����L�\�`0�k���7�wK%|8��"~���8j_���u���%@�s�	��Y�=N�ɢmȁ�2uqބ}���_`�=;_��x�Z4�ڛj�j�ViY��W�{N3�!�YKQ����j��eXƱ'%��Rk"T���� �Dh)��=P$.V8�
�#�K�N�ǙpIU��Z�Y�Ro^+�V�${p��0��T�3}��a��x�/7��"C����J)��c�6���[��MBI1c�rI��I/v`�T�����-vl��Ila\M��F����SI���a��6x���}�K��1e=lxM������X���=^�3Tpl6�]�_���tm;�̇c�?��-T,�j�U���A����x_e�6�Ê�b�rq���b����:���Ž�^�9�ƾ�\���� ����X����Hp�x��ǳT`1Z:'��1a�t��^�2�ܴϑ�CRȮ��jQ��<��s�i��I
�/�z
�fbk�=Rn��ig�ˏ�#b����QД��nͣd:��i���#�[MY<���P���5!>�{R��h�Mh�	!"�jm�1K<�%I�-�#���<�R�Ň� Τ+�aS��A^�����y`{zbw�A�cu��M�
Ӵ(���[=hd���ݑ��Q��
�=���lrc����(�צ���~gG���k���]J�����8c��쟍�ׁ�#�J���ΘSg�p�y�O�n�~aѪ��Z��vwҩ�t~�YO��"���N���V{Y�ǗO��^�jC�KJ�������~2If^~�4����ǟ�������F��i�j�u��m�(�q)�:ͪ��Q�:�R7�*��h����4[��.���PN#��GK�A�o���N��sz&�Ȇd�@g�E��X}NR�r*�++�];��Uѯ�FE^�
��nWpArF�%/W�YX\r�;8H#8�2�ì���}׊����k����L9,�����iu
MIk܅���r�D �,�S���h����\7�^��AI��lĚ#B���Α�eğ�Q�Z�L�G�,�@|�>м⤒�A �|t�1���̇d��V;�}�|����=6'j৞��\Y�@���)tv�P�Ѩ�`U'��ιE~Qg���֠�����5�Ʒ;PV㜪�����A�$-^�����F��Խ�V�\Ϩ.9�ӮZĒ+�$X�X1
m_��lZc�p��Uk�������ҮߕC?��;��&A�*�on�Q\�nf�J:��~[���P��:&4@���532?�z��&)?���9k�C��xr��3m#�>�$�)A�����
%_i˪����p�,B)Gn'el`��~}D�_ �t��D�q/�Q(g�T,0ĜX�*������G4Ù�r�����3Jc#��SI�ɑ~#Mo�@Z�^�ۖ���~|����EݞU>`+qǘU(�aGk�hu�[�L��� �<
H�B�S;��
��	���e�f�sJ���nq21L�lZl����-g��X.��J��<ϊ1֭j'���Ĉ8&Id��0�m��x�Q}�s�����+���"��{�	=�&{�g*����:�����)pWT��Gc�+�*GM�i�<�9�3�����D[�S@AL?R�-�P�#�a떋�⊞��L$@FCׯ�0�hk���F�E�v^���K��z���B�لD,�r��g��;.�[�,�va�\���STkV��R	���������a���I6�ݏ�ͥ��@&�6�#���u�E���+��R=~��Z}��8f�8ӡ1�(:����s��7 
w��@�B	r�}wY
���$����7j�}uR�W ��c$ċó�n�_�[0�*[�	+~����Y�ӳz�y�4��x<Vo"v7��j
+��S��~mx���Vєۛ��
�1�zp`��
����ҍ�wԫ�I���,|����$�oB(�� r�oUJ��^� �*�$*yF�°>K��D8Kc:�|�٪�ڣ:�;��Z�A�=6���j�^�g�L{�א��&��H��d���ݚ^�^�,��ud6�0������Kcч~�."V�L��ݵ^(�����Cs/B,�f�=Be�.�[�͉�z��?�nÇ5~$Z�A%TI!����ho݌�������&�ɝ�\��mP~��Фƺ����	�~&�Ӟ�s_
tV�	����I��	Ի.m?%fΟ�� �d���-�ߝi�j����·S�6 Ni|�lK".z�3>���.�A�O%^^_-�����J;h��<�d _�r���I$����w&8��l�C�k!�TI��H_���x��-(W��ǐ�K��y�󤢕.��6
ިB{Vk�8GG��y~�Y ,B]=/�E��8�@����WT�L\�
E�
�  S�� '��?8��E��ծ���R���Z�T�|�r�uΰ?A)*gш�rZ�\W��K�pm[x �͍m�d�q@݄��V��ʶ��snl�0�D��V���K�Β~�(xd��Ro��@�
�v�/;�;�k�ߘ�+>{1!P���*d)����D� ��5O�<�����t�?jE��3�r�
�u\)�V5����5�)-��vMR�=!-؜^�1�3f���%w�:1�Ղ��[W~�C����-�HeL����=J�"cَ�K�R7�d'T���:�H�5/�7n�B��5����c+�^���@���ؑs��	�b����M�5"�3G>�xw\T�}~��%�|n��/��W���Kr#Bd��e�.�6��U��_��(u�69�b����6n'���V,b �@As�g?[�kQ�����Ŵ��l}H~*	df�dI#��0�#zgg}�o50������S��д��`Y ��"e�<�Oz���u��1y+����7��ٶ���
�>�V��Ē�!4�)�`g�,l�i���$���}���ձ!�9D��3H�]C�-�ƍ����A7 �r�dCo�i6�Mt�'�X���b6|�RH�q�z�^�F^@}�r)^9��ͦ���Ukr/g$� -C�Cm�iB�W�n��%LiY��C��³��U�ws�o����U�o���bwl�m����W�d����z�SD`���z�ϋ�m@�ٝed�������s6�@B��ZnK5�ҳ�*H���vy]{�'ųm���ALG]��s�R�c�w��]+�~U'��R�5����t�Hx<sO��s?u��"��������Hvg���k��{"�/!ג�׵Ƌ���X$*oC/���IU�A�r��*�0b��$K;�R3���ò�sGD�>p�(E�h�	�v�ÎvF=GK����]+"��<��.����]�v�P�M�:����>��s��c�u[N.�sW��-���E(ډ�֥�Ҁf&tB/O)���v����2b�0*<�#,�X�d�탠��h���,8C���B��)bq���l)��F��VV�k�qZ3z��#�r�_q=��������u�Fd�
ס�W��\�7_l���V݆%�>��+�=��ِ�d'nmU���x�#-a�dr��Zq� �l�'�����Z��43[H���e�@�*w��r�b�0X.f\����,:��M�s5���K�3DzǠ�ޯ��:F��=��2b���-^���E�aIC�F_C%�5�8p6��tZD���l<����ƥ�q���Ƒ!��>y�c@��筊�G~!N�;zA��c�4<R���ȉL�.쿑��N���L����l���:�E�	��d[o�'������	����g̒�]��)f��EE����!I���u"�|�h�^Z8!�����vE/���!*%e �X��t~.��L��qз�O9�� C�F��)v&z�Eϸ�㤉������3���w�5��{xw�A��^���}������&����L.�{���*���#=�Va�}�I��D�H�ʫ/1��$�n&c�`�?��N/�!���Z��&UE鄼s�$�y�X���**��%n��v�E�*@�YyLd�����8��	 R�Q���vnl��	��5H�I����_����V�5���+)2��a�%#`�W���E3���h~Л��t��c߇�,�UPf:2��7tKGrv�m��!�$�#���\��1�w�G��)kK�r�R�f�]��J���H�	N�j���<�2luc;���v}!�R��'��R��e�4�y��3U<�5ZeoUB78"&/n6\�ӡg��+N�����p�b��혱3���Ex�#�H|�n}�ySU��[�L\h�E���Ŷ^�x���_Joc��Z�ӌ~��A�I2�n����`WdL��9��!9����5�:6
����#6��Y��fb�s�N3&���q�'
ܿTK���w*XvEv]�5ՙ�4Ű���S��i(���i,m'�q���r'C!�t�г*4�V�+�7�yCM��E)�?�4�B�+)h��J鵧�ܤA�[#[�P�k�Aԣ�����e���yW��u@@��z@�-Ձ���eB��g� �7wP�Ͼ��c�9C�_C�5%M�\S#x����k�z���=.6kIf7�e_�]�MS;�'_�!y��h�`����L(�67I�s3�Ԙ��B��濱�$m�&�a�N! �A�a�I����Đh�=�;k]���cT�f2�Ÿ� ��tm���*�ف��۩�E�HK{&C�
�3�]��E	���	v�<el!#>ˉ����'y�4�	U�yyL�41�:QU7E�2.���k�cE����oK��XP}�X��]�4�oz�!��v��U�m��=M]d�%�+[����Z2<pu��h�+��Q�,E�\��'=Y�<�y�Pl�
6zJ���٨>�g�п�co�$a�nO_>��Ë�w�}�[YɊ�ec â�.�֏;2�[v��  �X3��o#NO��)�iB���"R��}�m�����8'�m�	^b!I�%��Tp��֏�l6Z"=Z��Cm�GWY�Ȟ���Ga�8H�An��&�?1�-��"�o�ܸ*')���H�`��Z6�38�C�b�|_��X!�Xy�sTI� ���-��2xv��������"���]P�w��wñ�?������9����S1՘��'Q)��5� fC��j#�����ּ��#o&Z�����ùe���<U%{�S�8i8~�6�`�y���P���)q^A4ܛ�8fا�B���`nd擞m碈�����|2Y�	~pD���:�-���V�kU�6��
'o�)��7�'6�y�߀�fa1f�ޟ�]���6�AE}X��ib��"S�X8IW�8'�H��'���We�Ĺ��; ���~e�W�XTG�G�0<�#�>E:��%���v  >���h&2S��Hbԗ�L�Y`Z���� ��F�©��^΃�O�BK6��} �ԙ�s��'��D�K�U�fO�ܻ�kl���f@�:�:C������CI2
��C��'���ZG���`T��h��_�Ĭ���(�&4�L-D�Ǟ� S��x�MOd������ıvI�vfC���K\e��I��x�δn7Y�����0PK񡄧o&��D������F��BE�Ea�B/�-r��wdc����@������z"9ޢ�c�p�+a-���R���j���3����V�=DV5o�KQ�&\Gzk:��]�o|]�sP�X{��h'�^xlY�
�������b���㪻��D1����	!4�F#�����B��������;�� ���t�����V�dBH�!��f���ț�9�g��\���D`�?v��Rr-���ڝY��Ϩ��r��u��i���?n��&i��v
�8��pr�]�3jLX�*���p�cf�jUڶ���R'�F[Hz~J�I��|3�3���β���oӎ�������h�'|F�|�x�:ˎ({�[��y'M��`?�� j��OO�}��#4uI���憜�l��Ģ(�}WCF�{��=�ڈ j�W%4+�L�G�VߗUh?3wLυ�����aOnړ�K<G
,Y�4�1|rׅ�.-�ۚ�L��U�����	������S���Ǳj���ҢV ���I�':�Ov!K�%責Ϸz�G�,oF���J���_U�A�.i�����A��x
���S^�3��P�w<*����<�#��/tEكk���L��m�X��#rU}��E��5���|��˷�B����PHG"n�Š�`[Q��%ıچ7_T
��?�|�_��mn��f�$��{}���8Wl�b8�m8І%$|�X���yq��L	�v�K����B[�M^�{f��(�~��jT��AM~��U1#4��juN�#�q���/�������]�&0��K�#yF,�PF|��.uq�"G�����:ט�$y�Č������6��)��fM2:	�pѕ#���l<������w/���	���r��H �PN��	U��m���R]�F�,�!�g���v1�����z���I�&�K�����e�}a��5c_�a!.��tF���r�����V���k���Pz<���Y���@���.n\[����e,�{�ȉ.�{~=���r\!ن�뱿�����3�`�)�MHU�dL��2P���\ �v{���N6F����
{2��?t����^|�
��L��/�Zu���#��-2M�6	Y��Q�CM���a�x{tm%gEƝ�_�%č��WV��6��j5���S������]�rY6��-���O�E2�Z�v`l��1:�ҁ���D�IX�E�}*i��f�W�+�ь�?��>�,��t0����M��D��7��<��;���;�d�
n_���Ʊ#�u)�M�He?�ĳA˴P�L\����E1�s�'�E �6��-�������W	�C�=�̽ ��w9z6Wc�\��:V���Y%*kEޖV�NC
�=���:g�����}x�������x ���_YR�Պ�<v� ��=��ȘC����+��>1Nk�)�h:�h�DK���IO�$�%��0$�  .^Cc5^<>��Ɵ����Фn��� �|͸�����+��7h�ʞ�j����y%C���!3�u��	��M	j�ֶ���ΰeD���� �e��޺�	WVO���_�n}1�c�$�F�(�Q��yi�)-�d��*�������\.�'�P�鸟G���q`�����L�ǥ&5^zXM�ۊ�J�"Z@i<���b��,!TV�	�}M�����S�y8|f�&�gٺ{�mD�%I��t =�O>�t19��7�$s���m��ߓ��i+e9wO�"��jM���/�v�!��8k.��&��#��+��3�
j��q24@S����[���h��h
%;PA~D��(�8Y��[��w�/��Gq]���Q��+�;�2-E�zʹ�%"�N��瘥�m�������i��q	lz
��®.�4��%��tl�R��s��)Z[�S����gn������0з�@R��%�����K)*����@��$�Zy���;�X��g\��P�o8�g<� �JUy�;4 e��N�H1�Pq����ya�[̀H��]Y�D" �y�Vz0�F�T���a��̈��V"�ư�-|C������z�� ^)���c��ԡ���ڭ)���T��empyv����>+��T����s��owƬ�(u�(��æw�u-�)p(p-�4��Ӳ"m�g�7���9x1��ݏ�P�/y�ۯOݕB�c�7Lq.)&�"{:<P9��@���B��N�¿�֜�+X>��$��H�ā}%�`i6�l$�p�{US�?�Σ��z��1HN��}�T�
N��L�d��9�� �Z��M�*�,����uc5;�ЁL�[���2����#�0#��\�-�g��V���Hr`�B���$��ǌ�����GE��.��inE�1�B_���&�\v�(�q�|�w|`�+"&��R��$�,bC�Ż��^��i��aٷ�Γ�ͣ��Oϓ��챦���t$o�^���c �UG��&M�a�ّ^t��%�g:7���d!t���p<�2��ƛ"��*}��onF���ץ��{�H�1S^���6�ȝ�/��-~�?�����+����E���Ȯ�ѧ���a����6TPu�ϕP��Պ֥��Z��,������K��n2F�j^�A�;M���N�+�9���rE�8��=���ơ���a7���Qo5�����;�u�*��������Ev�?���1-���F�9k���; uCi����������rO
��C�������
���#�ZLZ�m�U�ab�ȅP���+͝WtLfd�E�[��L�y�N��G��Et^2,l}x�Y�d\�|�F'䗈��'њ#q5)
��IL�'���!}�j��̌7�62y����D��x�%��ay�}�͑G@�6�^���R/�;g�b��4�Dڟ��
^�l����G0�#P�I7�����"�^�$Fk&lNd�+뢯`�;�Y��h�Y�� ��M��n[Ϗ�d������Y&"�4ρh�w��|6�92ʩ�I%�Ϊ���+ $(ʤ�8�?��y@O�L����hSU�$�KI��bc$6�z$K���Y]@�/�ȔT�k}5R�H�ݖ#���k�G�����}�7��}�	\GT������G��r�~�$�Z�7�qa{'X1�}K`���+��5�3����51�������2�G�:N��w������W@A[	��I��0D8�Y���q) ��I�XG���ۍ���&N�=W��`^����%e��1{��,ޱ���Inq%ޫ@5�cz��n~���2E9|�;��>��Bkp�M�Km?i����3x�W�m�$ګ��_�aO՗���G�}ᰩ���H4��7In� �6�]�ǂ�W����J��
���s>�z������	�:d(^�|x=]=;Z�6��{.c�J��8�s@[�x�t͈ݦ,%�"9���%�,��ƍbb�cW������=&M��{o�`�Z��C5K�ԥ5�ޱ]�ڳ��3>���������a�$��$&@�h20��rf�e���<Qb��T� �0�YgIړ�C��s�8�JNZ-?	�]юl�-!�S_bQ��G�ÿg >���s�,���V�t:�j����.���U/��ķ���XM4��;*��|��b7��?����o�&��޽���4��E�e���s�/Ҡ���g��"1y�V����߭�17O_;m�f����'���N�(�V�k�Y��.����6����^�ܨZ63�o,s|"�`��G�N:��KH2n��ý������WpJ}�ͮq4!11	=KpE���J�Of��=?A��$�^D����Y(���a�@�ڜj9�74�YBA�_��̘�<� �Cm���/6	�"�I8XN���H��M��ޘ�n7��m��'��۳��8��>�@��H��K��E.�1��}�ט�?
�ڻ�0�m#�p�^T5',iZ瘗8&��hf��2L�@�2�����n B�#AY2��F���%Q��W5P�)k2�������`���I2oHĲ�CyC܇�:���w���[��5Є����9���W:_r��71��	��8J\$]kE��:�U��J6�3���G�2�0�1A�,�'"��qi�FP��Ԟ��	�,�erjA_1��7��P�9iD�$ӿ�.U�Ώ(3M4�~v��O�����x�p��6��٩��']��V���Ƭ]���:�������c"�4�ɺsSY�;���FuzڧC8Ast�o���Q4GVv�oWo�C�����X�x'�����`� ��<�P�E	�
p_~�M�ӏ�+̃��;y��+W��.����~�����ف�.�-�<��d�<-�1e�F�d�II�J	�Me��	�u�cH�����3.�tx݌���˳�R�X��(A<1��v(=�"T���Y)~A2	��2�#&[����d���c���D~�ryjA����	����:�/�5�����E�kGԨ���%���.�,1c0z�:������	JQP��WؗtV\���gebYw��#?��ޥ������jߺ3�����/Mw���x҃��o������]�/��RF�ט�7Z5�Zw�+��]hp�ap�#�|W�7��g_3���f�D8��e��Uۣ�ڜpBS@�{!�j���6�e|��Ǿ*f;��Dʿ�@O�x-�B�Bw����r�ɫz��3
�p����.Ϲ�7�]3��U/��t�,�l�-$T���Yx8-��c�`x��o/Nd��c�	zG�7��16�_@�e׼� ��3���	�L�YPO�$gӇe��W.�;#�\�Q�U�ܛ!��3��@�>����W�E��1�/Ȼ�&J�eM�6B-��Ey�vC��?�&#�!����s1b�5
�4ǯ���V��!�p��]c�'�M(�N�J?�`�j�U������d5�z����
�HkY�4�{��?b�� �����K>�!�w���lL��QjWYO ���L.�׀V�mI&Ȁ�c�����լ��3]�^ �F�2\�h;��e�_�%���*�IOIa���<��h�I�1�7�U~�=����`la�2���AQ�j���~I�ގN�J�a����o���'m��;�b�'�Ȳj{A^W��F���BU��$ L�<Nk ĤCyE\�[��P1��T���a�5nL����[0�BA�B�ժn��&62o�v��S����u� �4���M��u?¢�ƿ[X��-}�����Nm �#6 =�N��5����st�D�H�������v�*5��#��ճ,�8>G���n]�䞠,�Fe�e�`���#XxTH,�g0v?Q�q'`��~ƿ29�&B:�p_�d1�"�x�-0oL����gE;���x�"IT�Q3~	�,ɬE��z���4��+�0�j��F�E��Taj�+�����cI�͕�ںj F�G���'����G?l1������$�����V�Ԧ�-n�D����gQ��|��R6$�Ö��M�Ѻ�y����߀��i�;�B8RБ�ǻUC��+2��4���%%�6�$��ipM~�������0�y��H˦���t��//.�aM[o�~,PK��� ����h\v���!�ؠЖg�m�˲ӵ�7
�O�y�������U�V�F�`c@z��@��|��Ӗ�ae�W��9���QHQƮ���6�}��}�o�Q��>��#����$�v[�j#uPxj�@ߔ��v$jXx��GuBks�)�lR���vQ
!,�c@g��o#m>p| RԞ�d����#,.?�گ�3|���?h�R	~v���pE�B���l�*��Ws �:�W�Ia����F�&/N�#PN�e*��A�]��vw�'��FO�:2��dw^rd��5�?Ƭ�Np�(ڜ��ܓ�C]�4�v'���-%��Qτ�D(�GjY��2y�Iem3IE���{Ѝ>"���Ԃ&@�,���0�y��s�X��B��V�V�-����8n̠����֛G�+�ZNOA�\��DV������^3[?����X��!q�<��5�3�}B�T��,�t:[�����-?�%���=��V}_C�;����]��Y�����<lb�C0& ik���F�^(R�uΣ��\	x����E���w�oI�ճ��:�� +W���Χ�t!��a!����Ӄ�� �3r~0[x�h�h���ޏV�z:J�ۡ0-x���r(�gy����Ϡ���F+�)f9���t�c�N$�#����%���	U�_��"�d~�";�{WN���~,cs&��Vb~�?���-��/���p��c�rƪvF�i�-o�?��%z�p�������^�ǹ��3>Cn'���Q��S�+Ws�j�������Q��=��,ҮF��X]�[$�3�.M�n�Q�p8�� � ;�.*`�Q>�w�Z���F���"�ґ��I�"ͩT��^�q�H��a�0���(i}a�L7�U�2�eDVrΌm�q����%��r��M����2r)�w5�#��b��\�=�?>�� �P�͌���^��:F�P�҇Q�)v�z%^�䊢b4~�0oR���)ie����{��k�W��;�,�;���N�����P��V�|qNQ�X<|�3X��Wc��^���^i�F�����V�S�a�me,��I�i��� ���9���A�9hߟd��]N�J|�������-b�3���<�|@�:��@��7B�Z�T��P�z��X�j����q���/�ps؀F$�.z��q�����ht�0�N��P�,�xL<4��ƽ~Л��#�ʎ�7pUĔ���3��<���_��Vk>ҫ�����Iy����2}�$.'�Ï����\ϸ�K�/��{��OA�&�k�a��@Z����h�Gf�ȟ��}���$�5x���� %M��H(��Ǽx�j_j�?$��=���K�8)�س{��yp:�
����{�]q[�%�����_�=���<ŸM|i=Si���Q��yy��$
�U�S������D�n��� @�:�
b�w�O�Z�W��Y�<},��7��%�u�U����B�k����뎢���9J��[iqTZ ��Il����V����!aB^X��|�-��3� �YQo��>���3��T�F7"cǖ,]���.XUA*V1�k���+��G>vnBG��yi�o\�o�LS�J����|��P�$�z�n݂qVu+m>p��#�TZN�܇�|��=���5u�s<�A�$�:7"�c ��%����L3ďF �]1o��eC�Nh�]7�mޘ#J6�no慵�<"�?7�6?2`�|��"����Ϙ�@�v<#��w��3�=cR�p���y�ڈG�|:^'d��ޡW��;I #��6��l�w���N�|N20rr�	?�߿%��C���2wKe�G�xd�h:0����%�	1��!�o��&����|T���~�N&3�3�~�Ǧ.�G����G�lx]��̬�Wy<6b\��z�Eq�=;�q��X<V=�gZ2l�I1g<t9� b3h�\����Ѣ5��K�
�e�Q��+��K�.��k�'	pY-�j7l�D�;
�*��v쏊⦞� ����\���v�K���ZK���X���	fJ�E�R�|�؜�]Q�B
�A��s�L7�Rl�����k|ѮR��A�=�U�|	��F�\����*�����- ���n��
K���3��R�@6]�����Vh
3�}���V�L>��v·� >D�so����UŪX	���b��h9����	��?AL&�*r�vdĹ����IfJ�<���n�Py#qQ}�0��21�8A�P��[0W8��]�:s�O��w�:6�Sʤ>5I)w���j*�_V�Wl`�o�.��>¯.��о�F�3�=L��EkP^f�.�v��9��K��0��>�|`����������)xr����PIܪ2�k����'aut�ڷ�<
����؏�z�7%�Dܐ�f8MH>g�SOVR�����o�k{=�&1�x��X����@�!ﱀC�F8[�g�����sE3b�jq��q�1�K3�oW	t��q��ݎfխ�����a�] f��J>���k���}`�]�5�bh�Wx��@���F�p�cǰ��~bC��^K��ސ�3J,i�|Ī@�	�:���F0Y��h�?Q
�� Hp�,.@.�}����O�P�h¡�
W�-��DC};w� 
T�Ԧ�����P�C�.���w )X����$�C�h�;�0iͪ8SV�،��|B�)����3p�t�O2G��JUt���?��Z����*��G��s�����䀏�)��8�s�\-�q��S�v��#]���Ɂ�X�Tf$8\�s��	�<$���w� A��q�~Q����z�>�?!��u�ΰN��	p��5�o�9��Y�P���8����!Q�3K�5��)98�@������.X��6�Y�Skۣ��~}Ed�`p ���}��;�ˡ�j����!*]�ƹZ��q])��^����� a��V!}�.J��q��i�$s�sMƨe/��K��WA�&#)��8Dq�S����j�.*���v{n���l�����$�kq%<d�Ą���	����4|��R,����_��Rt�
�,��D����e����p�����+���^�����b��= 8"){;���P�Mԁ���MG�`�s�����u�p	(>��Ϙ[k�p\Zz0U�,$�c�	w��W:� ��;���tG�K�Ypܺ��|�I`�	��ι�A�%j}�j{~xC��n���C������vW�r>��"�\΋b)���ͭ�w���t(5TK��]�ecL����á��h�?!�4f��Oӑh��e2����0�]x��$T��L7�Τ���ݏ�������0�7��h����o����#�2�$���:�p�K{�H*He�0q֚u=��S_����.�͓�-:�d�T���a;A0-MA��b�	���/�}�����K���L�gʹ"^��l
��Q� �vS�M����pi��%�?����=���TG��	/8/>< EI����������� x���^g���.6�{����)�(�����c��5dqoɮ)�s֝_k�	��P"9
]&�F� *%(
�)Z�Cd�`�O6�Ԫ5��T,82�-��t�K%��+�Z݅*��u7�UrY���kYv��F�&��O:�âj�k�^�G� �Lk]^����c����ז��=�[�`'���]U�r�ߞ{n1�\�a�}�i{���_Ȋ4#+�Y%��W\�zتӧ����N,��5/�@Pb`�i�s/}>��� pL	ޯ&;�e�-dR< 2O��o��[?����F8�N}�~ p��w �)b�	�+��]�T����4 d�������ݠ?1� �o�G@�s�}�@��VJ{�Ϙ�>�w��t	� c񳞗{�R�[���/�p��Nl )1�qq��m庭��.(I/sP��1��%�*�M���/�����gc�]jl�J�3�?�z�&���d�S�Xi�τ�wed��[�M0+�-��]���[�4;7I[>+cͪ��oI�������nB�m��SB�eeJ���p2�̳42�|L�A��2�\8��I�f���a5��z������1�A��Uy�^2|��-R�!k��ʼ 7��s�"1(�h�/R��v5�2�S��q
���."L�KƵG2�
�^���v���(�e�ڝ���.����� N���.߀�H���w��.��՝j�FB�d}
k�"��#�-U]���v��k�)iVk(l��7�/���D2Hd�~�Z�r<T>^�����B��҃��(��bp"����&��q��ʚ�jr>-���0���%(����TR�|�k$6w��vAC@��U�#���.X��5'�+�V��[����Kic�%�n^{�܉ov�J��*�*<�L�i7#HreΌ���z��2�Fi�*f�۰8�'݋N�$ K�������� ��=�?'� @(�L��<�e�!�P�@y����,�>�ZΪ�)��c�����f+�����a`1л��HS,��)3�o0W���^�V��Ob�eV��RȌ\��Y#��fs���D�o����"����x��c�Rn�ǐn^��*���M�<�2�@���Ӊ�����ګ�a�]y�����A>�9C3ӿί�V���	[۶�Q�T�iɓ�R�Z�����K����gyHڡĚc��;�^����A��}���o;퇤��"l$lC�G}��y��8g~�zj�����C���� �+���Y�z��s�C�|�ȴl��&���UDn��s�5J?h)�Y��蝕�s��l�*��e��҇�v-����\JK��H?\7N�X��8|���u�8���UJ�q�+�g5�o��X��[�u���]$�!g�'�pT'z�+qU�� �̛<��
|<�� ��@�toZ��փ�@1��c0���<V՞�b�5@c�JY4��[OG|�f���}[�'�&%!a������^#~�<���I��Y��Uf���0��}�/f	*0�MIBu����N\e �K~I�r�80'�Ng� ��@;�e�cp�R��qFh�ҩŷ��Nv ^3��t��� z4k,Yb��c畧�`����ȕŹ|��c@C �2��Q$l�'4j��4ξ+׏���*��� ���V���H�b��Ĭb��V�ap�-!}�h�|�O
&+wl����W?L�X��y�w�9��V����D;���5eLU���I�H5��Xn��N�'�H`�l����uWbX�>���}w�뿚����铿�g/���y�s8�g���
r^�WN ����l���ʖ1;��D�t^u ȑ#2e�>�� EY-|��xǮ��-sK�����\�LԲ���ӷ?�0�25/G� � ��ЛЕ�5*��Էm�&�NxZ��L=h)u�v��O�c���B+1��⏶�\ZAƪS}���y��������3gT-�X���5|��xl<�I�K5��y�T��g�I���N��y�����p= +�:?mĿB�W���^%ePC�8s��)l�������y&�_�
��X@����ʫ��9���U� �������2�K�9��c���֔+��FfP�� g1 �`%3�L�̧J�>H�Oy�G��t�饶L���yK@~9�
�����T���EUу��7��n���f� 3�K�?\����?銷�����;�i�֠3ET#�H���M�,��\C�������c���!C�
$܀J�!ﭔ�H6�4䘂+�t�(���DR�#B���:�d&�I�x��`3��9�3A_`�,�xS٘p�b!�3:����������F�ms���x�Nf����I��j���X��6+�	��XUlZ�v�IM�U5�����a@bNW�A�N!x�'Y�a ����Dԙ&][6�� �U�z���$��W4��܂���0��3_X���srw�Z&�;ϜA��n�(P��/�7�QN�Ò>���:�V�� U�ʞ#c�w�^8�~ߐ݂�4�M���ו5��/1��V��_d���t��<I�ҍ��:է��u��"�B/D<\�B�
U(k�L��S��n]'�Q�QO��y�҂$�Dy$˃n��X���_Զ�����aY�P&>�=��kzY��	�����ǻ�4`<<
�c@���t�� vI��T�?�t8�q���v!S@�)�R8�kk9�b_@�qZ[��\4�d�U��%`(4��_��g�zN��[��hɏ���WW�]�9����ts_�� �Ӹ�� Lg'����oqG��B6�bz�����*��5UN~�Hud��w�껹�8+{��e�&����̣�oD:�}E]��'�l&�*b���F<��=7�f��pE��}�)��7����<X�7�!	�[+��mi�k�qzs��H_?n��y??`hP��0l�c��Zn9��Ğf�%�ئ��:R�H�����}�>��I�����5���ى�Z�ե0�%����)9�����ԞL�����Rem�4�-c�d5Op�J�b�l���R��D����Ai��+_��|1�w�.Y�U|0j7���?����c`��N�b����6j0���D|��� ���} ��&p�iB���P:9��@M����V�)-
�lAZ8ºiuP.���k;�7U�T#)aߜ���t�Ԇ��B��&?C4�솖,+9�c����2�:5"ϗ8�l�
��eC \��S���n4�Y>�;���')���N��������Ӎ;%\n��:�(� ��|fz����[r���RÑ7$ ��<4j��}�Ӆ�\�qI�����P�`ql ���#�U{=[��>� �����!h#t��El4+�fj?lG�0g�ΚPT��b� �uՅMp��+�w��	�6D�4.�ٔy�lLfD~�s�`�hr��$�b���W�M�$3�jK z��?�}\�3ke1��@�[5Ʌ��+qhg���d���Y6�q�����=C@w�v�WoΑ������<�ny'��Q���q�<�Q��e�v隝%��q��s��%�������lBJϵ\.�-����t#��X���Ɉby�x��d�i�n���T1T�mid��7��j�����B�(�k8�!�O�-�ABO�%L�;n�����bg�S���8%yxq�l���'��,�'>�I�,�e��M�:���=��V�s���4>tows�m��5d�ѐW߁k��uo����ͳB�U�+BJP�ғay�d)�Ŵd���v���߄stKS����Fpt���-�8�O/���k{.H]E���gG"�K0��YO�ۊt2�:�LE�O�kL���qXV�l��*1|�I��KG��Wa;�#�/i���¤�v�!
E�>���h�2Om`��8�m��R�� ��C�җ��F�*�L\E���B��E���G�
,�)?�I�?#Dl�
tUzO�����-�0�Z8�(�� 2(C[�s�Wi:���{���L鏗Y���N�4��n"[���1�G�řni*� 8su�3T?P��H#�WwZ&҄3��H�J��rZ9>'Q7I_�d`��0�LX�
����^0��.����|1Y�QsK���rH����
t0G7�x��lT/\��r�-�!N���<�lDۼO �OLю
�
 �%hb�%�̄�Ԛs� ��0�|[�6�����4[��P�u-�;��[�J���8N�ZAz�dy���OU�<4��$�HP'�ty#iU���S}*C�a,�3��[��Aʒ����i���]8�σ�������ʡ��w"a�̝����K�n�m�'jv#:�Yby�@�S��B��`�nb���gF9����J�c���R��U���|ٝ�v���A���r+E���y��}��}S���	ejuAR� -|sʶ0[��޷Ui�z#s�|Bv0I?�3�5/^��?|�����KK�-��	#!��2E.l���\����Z��n� 4�c�o�����ƻ`c�0��҇����������s��{��+��,�N�J7��*��F@Ϡ�v?;�0�rt�c��r���z$��׿��3�s�O�Ř���8@}�a��F�1+�bω}*�HS+9�b���ef��hƀL{k �W��?��8����3�t )x]�����Z��
lbb&i!��Ѕ���⋭��~ds�N��Me�^� �G-�;��M[���J�H����:� /���~��+��"x�g��+��M�G�YXz�pd˞y����}�0���K�7oq"y7QD��NY��bF{�̖�	Ϻ��4��-�*wb��k�]1!���RDH(��DFLyCe��{��+�M����7�����'ӭ2��(��ť.�K�l�����BI�oU ��褮�<�fu�D���g��O� _}~�|����$]ȆI�
��}=@b(ڄ����3=N� ��7�b�"moy{c?e`tT�h?��E:Gq1�\�`�r�}���m���TJ�ȡ	�a}ʗt�EL��Ӟ� 9���!�m%��c��M-���HhGNE������P��i_�v��5�@��\�a�!}��7޲=���_�li� �N�����J�n[:X���.ϲX���2P$��v�P�JA�_![�Wۦ̱/0�B1k.߭�pt-��{0�t0���v䰋�ge0h�1s�T�H�V�����V��T����VM�+Q�;U�S	�|�i�;����t��`1l 4�I���,6,lfr��'�1ՙ5ê�F� t��]�nQ��P`��1�����e��bsa��	�&��"zp�<��UӦw�,b����RK�Y��o��/#�D9���
du�_L�F�x���PJ.1E;S�J��{ɐ����l*g��0�'���+�Ŝ,���1ձI�Q�{���.c%�8@��*"��6�����g :�r��c�Ka��X��+rڢ��z����U`�uI�(.�(6ĺ���VK��D��[tQ�$}K�vMI��H0X��ʟ�T�q�<��ї�%��n䒶�R���}�h~�.�!�:��?OO�p�d7ٻ�\�.F���6����J2;S4��r�Px�CAq�,�j��2�N�X�ن�2r!.b:��̱'7���y�$������uUď`�-X�e_��;�4�L�t�;׃��z�~ƀ@�直M��/
�݊~��.���&R�/�vG��dXO�Є��[�ǠK�\~,u�V�"��3��1��$����V����=m~uciK����p��{��빢h)�{zл�o�B�q��ӎ7��\$�T�i�k}��&*���˓@n'����"�S􇆒�3�LC>(�g^�!E<{��Yv�4sdyuᨲXG���~�o�nQ���s
����\��{|�M�Ī����j�>���~��Q���+\���&xP��>�	O�/�<�p/�M�gF�P��.~�=�2�AL=H\���،_w������w91���b�yp�ɧ֔�w�d��"�ϲj>6X_-a��%�nP���^�&�c�v�o�ճ%# ��&\�if�<~t4�>������Z�2Mh��#�]i���2Iɵ�ŏ.���j����������{ё��&QPE�W��ːp ��3��2��U]QUh:t��VpN�P�rm,e4�l�Š��0x���5�}��0y���0�l��.�(M#�H����.>s��P�i�@��lQ?o9E���[���/э��d���f7i���q|��y�U]5�@�5,�:��7S7@s�4K®�C���w�`�nت(��6����~>G2�c+���ZXG`���z��e�^�6��[T�Ā͚�H��	6��C��(��9^�E��7�S)��,�:���փ����%Ĩ��jL��؁0�?H/#�G��g�)?e�|5'�d^.|g�l=�#ZiF58��,����lh�[�ۨ�^�c[ �i=��'��a�ELE,٬>)��?�f���OQ�߃@Ō{m�= �i�����Y�M��yZ�QO�']<���*�����r6:m�k̬��
.�Ԭ��������´R[��h^k!��q_�̃����T��k����ӡ�r�FtA�ъ�:�;���!>�.��P:pTd�so	3��uJ5i=7�r�&��@(K���&���)���M�جj/l��� ���Un��YNV�2���|�zu.WN.�W�H}w�쪊����3w~F��4�z�.,t)�9'pi'�B�zE�~��bi;����B���w+Y>���|lIys/�f}���.��,�yp;{[�Z8=�Ʃn�Nt�q1'(�_W���G%s�����v�'h���`&c�r���΄3���B!l"�vXLÖ�
�q�j�y�֡�O_P�)�(�	{6��%����i�~���_R�~)�g{S�Gv���n��ƴ~&] � �6��l�?���n����o
��*�Tȣyɕ�a�y��P�ѓ#yٗ�7Fǯ��[1>Td��ܲ¯�B� 	}K��Rs�͜�:	C�$ʓ��E��F�M��,npEz�����`�T����z�Ξw���ɞ֟���M*�MB��9���N�E��������� �&t���̯Ø}og]�cB־Ad�v/\�0�}u4�?_`��N��R{�&��oR�W/<4� �\n%A#�VHvMOt� ^`Ga{7�7��-e����v&�i1���2�y%���;�e��ns7� �N`���{*F��8�:F��o��e�A��p��
1_�����VK�s�nl*gB��])���¦D0cA�����܉��	D�[��Mt&�Ӣ��2�r޲^G\��_���:G0w�QՋ8zhy�F�h��>+M��Y?��6o�^�>V4�����|y{��,��s!O~	+@H���-��d���'�Uo&K�ך9E�����^�zF�o9�ʎt`n[x�r��X������Ew�ޡ��Пs[�ݰhv�k/�ћ�>��¤�^�O	�yGL���ow��G����N>c\U �	)WZ�	
JƔ1_�==���`�=��N��8��!���F�^_>-䟠�m��L� ܅��4T}���y�;���;*����^����pAY�T����Shl�mw�X!�$N�]5sqg������ٶ�h�������T�"�c|�YV�Z4a�S)����@��xK;�P�K�&镛��F�o��Ӛ����VE�:�+C]��.dؖ����#��9�뫦�$$	kw��E�s��h�<��yQ�?����N���Ә�b�O�Lo}_��@'9���:�X��~�����I�M�!ȸ��nG�@��Z�&�JɝE��P&voG�v6
�6WD�d�nFK��CG,�GF����Ԧ�Tta%"����Ġ(��S���\�e���(D��u^|���{b�@�.�!�PT/q�8�9�����n�,��X'ph�w]F%��O�� �*�����ͥP�#�R�^��l��{�%a~�~X�B�#���u*IvS����3���%a��00����լ��{�Oԣ�+}ӛ�Ж":s�|-W 2������؁�4A���|�X�"����	k/���V���kKk�AW�P��N��J�9��¤������O�H�wz���2l�OIK#�n�%��q�����h�]���,�K;-�J��ɀ�Lr���r}, �P�M���Z�n�%j��6C�g��
ƈ<�t5y�~Ǡ��`��H�&�ԯ�Oi���tL���G�!�h�lA�����xN�K��i����q+㧍��hb�У����7�U7��	���u�� -Q�@tzH=���umby��/��Z)�~���n��쁅�} aB���g�]��!z�[��W�րdA��!�<�%���D�]p��bS���V�� .���(@f��4��4����uj Hz��{�ŉ}0v�QW����f,��q9����OG	b��6��DDg^���rr{K'@��o�6�%����ڬ� .B�n��"!dOuU�*��byO�"��]4�V��KJ0pR�Mn�k�K�\BH��]b�=A��pD6p�Ԋ�蜏�x�6q�`�.}\�XnC�e7-`�!�|�ȥe��v�n���0��HZ���k}y��?���ir�7�l�b��1�u���d�o;o�Rە'����h��;v�3w�} ҥ�6�t�ֈ�c"��4���Q85A8!�)��y-*�ݽ�`�G�k�
F�i�.&�z�5����Ia�ԩ��r>���)�,�caOv�X�v'1��j�ê���Fq�����@�Ay�juF���W�MӸ�F����Lq}��m�l�Ў7Bh қ���`(U��?�bǘ�`Ý�<C#�]�C������֯�4
i���^nVD���:`�=@�ޭFk`�d�����D�Ąv�׫���\O˔�d� �6�k����/�k]��<���(lk&�PA61_�&3�4
GD�h0�����;%����io�{��׎���	��2Y:��/���9'��E4Buր^l�O㋮C�U���dc*��l'<N|��9
v\Xfhf�(ZÜ��~1���k	��lm�5&���pr��9���|�����&t��	2�p{���}�$�����z�j�W����iTw	����;?_�������D������6lI߁�D9��Ci8��~�1%K�����[�E|���r+(���4�@�`��PB"b�:�N�KY*#��<�$Tt�58V�*S�8>���j�Ik+7^�`�������eˆ�I�����A�e[ߍ~��=#t��OW�K��f���r��9��Iؒ²��4۩�W�o���*���l̴�js8L=�՚x�S�eKĴLCޟ�)a�qrqj��D[P�/�T|D��������O U��3�B����V7�b�w���ֲnĴ�FO<��,�",)��y��ƪ�l�a�=m�-�t�܁!��.w550|�N��v�Φo�+]h�𐘘���0��r RMl��B{7)��Mc��`6sa�6{Ȉ������2l*�)�v���w���) ��T:���U�g�هz������V�q�#ᰓ
�g��7DZji(g.7�gOm|��7;1������ӵؐ��9���\���P�=О@������֙���q�t{7�w�����x:,% �'y���9�i`��X�ȹ�P����x��$ƙ�Vz�MUq�4Z8�w�"�=%!�'�Jz�"��Ҏ�dnz���8]���Pp����b�I�ʗ<:@Ϣ��(1�×�7hb��E�bz� ܙ�����1���&�Xa��I苎�KU?���Ƿ��E�xª�G���D�"`Dʹ?9C��T�}|�>���[��n��NHh˚��r�jF,1�ˉ�(4p���ƨe�Q��|B/dh�f���?�su�l�9���k�������VBqQ����ti���v��b���"1	.D_�s����ќ�A����ͯǲ��q��_@�d°(��Y�����s��dj���@��6f�d}u^�����d[4��2�k�#��|;"���Y+��{w��M�Y7����0��PxNqdgW�������YK�6�l�C��?��w�r�س��ʜWN�f	(y���[����4�! �4�m��z$=��?�[�X��]׉�	[ma����ɉ��^��)��N�\ź4���q5���؎�`���Ъ��Ư{>Iu ���	0�Wm�޿G��e6�����-(3Űx��
��d�7`1�JB�῭;��U�`��	�x܌󷂫"�L���|��$����K���6Ɖ����S9�?��H����lrK.c�pD"p[g������qh�F턃B����8��o!�������́׏��cy��[]����u���G�����K�ZϚ�\�n�V�\n߽u��q� 2<{Y��:F�ΐ�f[��W_����~���/��T���%�o'���K�॑3, |*
�(M �`
�L7ŏv}�	�t�+.�՞gC�a���@�ǖ��Ҋ|�Ol���
���ބ��w�~n�h�O��C/�
Hg�����n��U�8K2��t���� �aS����96.q~�?�f��,l-H�0v�	��-�8�������!_�h�#�RI�v�:��/�8@�����ן��{A�Y�C�
F$#����2x��_6,ݬL":df�Z����@�Ý><~���\�*	�*�G�Z;춗f�X����
�Y��t+��9 ۞U݋�4��!��-��Ⱦn�ͽ[J�&�b+s�2�]��s"� ��1J��IDi������g�
����C��R�?"�֮?�f��YC>	��YbE�p޸j�	3/R -j���I6H�_��J\��Q[���"HB��G&`�g�B�ϿQ���/�	e� �@��E&��6���a�a���k ��Z����w�tk>�r(y-C�ޚvuP٠=�q0���%Z!�a�G�H*���(���[Ȝլ��B�FN�-z�N!tHI�����9][�0��{>Uc~&��/M�ļ)i�^�B��	b9�{��]����6�.�\FF�y�h�9�3h5�V�l*��9((�z�Brc%ޏpd/�yA�� ���G�2��kD`��NQd���1/����[:��J`��v~ه��}wn3�IAG�yL�М몂�>��սI�+*����T�s�nO	D j?"�ǌ�O��a�d�w�:K�\�i����1�n��������n&��)�uSlG��~�)�L9LpG��0þR�ݩ����&@��O��#�|��~Q����q�����e�B�Z�H�+�����u���׳��M����nb��z��lnن�.�� �����3��GU��%���J�,$8�#Չ�0�W`�
�q{����V�)M���K�?Y��Ƈ{��j�fY��+�]�#�ܜfSd��Ŗ�����s�(y�;����0�1<7����+�$>�Ev���3O$d>��Jz�B�zC0 ^g)mE.�����s�W�5��T�/̽k���D���{X1�I��}]�+f��cN�`Q��fKE�B��b����{�C��?	:�-t�(�r�+�9X�{Q�ҭ�@��Q�ˊ���Sľ!R.;�ɟ���/6T����Twu���y�+�/#�x���Vr���k�+}�_��a�A*)�PC \f'�kۻ�:%�ll��Z�nWJ�Ԥ�<�<��<����Α�F��Y�|l��v0{�z�-��Pŏi � ��Y&4�kIf��pQ�n����;�ߢբ�K�R�ڨq���3�����w�OB��U�+���	E E�W�����w�ښJ����36N��)K`rM��JM�s�h?����ẛ,�R���3�ѨQ�M��gGJ_
��3��䩞a��l��1,�a�(���Y����)=�O���Ꙏ��S��Ͱ�� CC�#�G���2l��O>�)��~j�ɥ艤[�kS�Im8�|B�T�Q��k�
���j���a����H�lp�yF]V�:�z5E��7�Sɮ���-�p��S�\t?���SR���=AP��1(z�v��;!��ܞ��ܓ@�m�����(��- ,]���ڶ�U8E,��L���]�]=��]H��'i�v��+�t����x���H��Q6�"˫*A�Iq���&SeB��J$�Y�׮���'���s\�3�Ƈ=���3˟�, �T�~d�S}ӗ���-�>�kZ�D���rf��Q����Wa��ӓ=OHb�V��E�6�uQ��E� P`f�G���`/P5#��F�3=�(.�%��С�m>�S-^�:VvxTCM�)�s��B�؂7N+�v����W����L>�9�M�7��D�jY��hHk�t��8����Ј�xu�k�Q�svwo׵��-��	q����v/�����(��X��V�,�1(��}%JK/�H�����#���	`-V��Y�*kxOyKT��+?��:��ވ��4��D@1�#XljO%IsH�2E$�ژ��G>q<��8��U�^{�o�'���@e��c����,\�mV��r���,��.�y�����_�B�LUi@������t�i�����,B�J����I�� {$�Q��ʀ��xۓk���w�9��`�����s(<�)�G6d���.���!��ֆ����>�xE�!�2��
3�*٫]�h�~T&�Q��ضq'K��nx�^ţ�%�g鞤���ǎP�*��󏮃�f5PyH��IΧ�_뺻�X�~ �qyx�T9�'��%���t�y洠y�77�9lfxʒ;�.l�L�uMڙAA_���qGٮ��0��n>/P�5�����ׂ�@�1z�∅�K]n��l$7��@ĕR&�}0ժ�4v��d�qTi��G�����9�eVGj��@ĉ�? L�wj�6u�c��� X�Rm>s�4>�4���H�.��_ ��ʑl&������s����f��x�jB����x���4o�
/+N�s�S��*���h��b�U����澳õzԙA����vX&u��$�O �&:��Ʉ��m7Ϲb�J�q<	�ع9�T}g�e�����*��U1jYx�9����
���^���#[^�N_��w��C+��K辰 1>Yj�+�IK���vχ��&��H��X�`Ic\���Npq[v�pb���������w�ga��@3{3kՁ�ە��=�)7R�#`AT��2�A���Kn��ߺ̼�o�70�����_z#����C���)���ŊC"������(�$FA����Q٠@Ck���SJ�j��)m
E��� Q�у�����ve~�k�P�-|OiF�?�q�~�\�6�Juht`��YC&�t���>9�/��&�ˠ�,�b�����FM�δCg�B�^����C�@Є�"��c�/J��)�l��B�ň���]��{\���!�n�$�����P�4I�;���
�H���d�M�v$'��+��[HJ�Œ0Ołc����!Pn"�����wƿ�\�l�vT��i�eI��<�.D�%"���=k2�����O��=��KhED[�@�z���w��u�R�.VQz`Z��G�Y^����ppL��v��N�L�3�'y�{�?Ī�$�6^��Yb�E�BI�����S��s��ii�M��Z��(�7�����5����l�i��`�x�:]L�������h|��z��vY�Y�q�����d|.�$r4�l`U`�'0E�@+�i�N�&��k*�w�o�L����I�ã�vK]X�z�w��GA��Z�,܂���zBR� ���ԞiX� ��-��Cm*������5�X��P�&�n}�88��G���F$\�H�
��ȃ��;&�����#�vg&�1�7:9����o-�R�8�J�)��l�s\�qh�eIk�w��'�G�����U���w��-$bB���j��hP��G�E�+��_ڣ�q���f��yZe���ۗ}B�Y`]�b&�j�R䂰:�҆٥�3(�>���?��6e)m��,��@_�L�ZM����S�\.���yN؋۸w� ���!�X�x�_�o��Bk�hTڻA�	o)��Q����r*Cdͬ�.�dS)���GfX0&x�lٔ4�15��A*�����ߑ�5�x�dBϷ� �2	����	1GլH;E�ĩO�]&̥�QZ��J+������=��(Is���x Ⱦ�9�7��Lg�h�ɧbg��n�^�%]6�#��_y1�ڬ�([&�	af�X�"${��Q �s���������Kۘ3�gg��z�� 3PjvZ*��jK��K�g5j[������%Z�o~��sM?x����͵,^bm������{��*c2�RD����LX���_/��\�4�2� �QI�r��^���+��F>>µ� 
��.�x�Nq��U�5�䖅'��A�K��"����wٽ�)V<A��j�K�\Zs��[	�c�b�Hp/O�Hp���5W��=�򁖳C8�W��#3��7��T��%����i����x���Db<�q�`��xE��x}ɗp��fѦ�?ۓ�6�1e�����1 �/E��R�������	+����)���	�<_ũ��³IX\gC(~#c|-Za������l�<�-
t2���8�ŧ.����P��Ԫ�J���i$��x�
���)eMT�]��X�!>��ؚBK���S[ߚ���c0�1!����@�%e.y�pa9�����
����HF��Y���"�oS���Ix�]C{F?I�<�� 5����~��L*}� #��Ck�����u�{��~�xBȿUr�����&qQ��h���Ϸ�R�s]k5@�{��J�`�S҄z��yO�Z�xUY.X5#���z�B�>
ͭ�D8D>{D�z��V���'aμؤ`�B�c����amS��X�p�~w��ʢAp��h�-�߸`��(�QMuQ_�ʏt��n!Vs=�}��Wz71�,������Q���-�	B+-VA�S��zpR��9�^>9>����OI��9	e���c���ܶ4�ˋ����m�R�G$PW[i���S���" ^DZ6�N���/��;4u'��J�*zx�)��#N���i/���tB8pkϋ ����ƹ�_.���K�&�5�%?�,lЗ�uOL|i�׸�����v��ܘ6+�|�,
%�/�Ck��7�̳*�O|!��� ��BbFf׫�e��xS�>&��*��i�����ey*��O�aT���<�K6�]䢼���.O�o��k�g��e�>��F�w�y�rT�F���#�:Ql �uO;��+E0��+�{^���[+R&h����p�sy��`Ջ����p ��n�d�MF�&4�m�s���B�g�b�ெ��_J�[~4F�Vjx���H�����G{�ckQ��w��ࢎ��(���e.M��PiX��^ǚ������q'�.�77f����3�(e�w����uW�ӡ ��Dukr�� ���n4��L�V� ��,����N��/��'#�g�rQ8f ���
rݹhF���y�\bg������S�x���7$u�Dڤ�����@,/�������zvI+�y���C�W<+��	vT�72�������uJ�ө"���O���1\��b�;$G��9���|ۚ~�bFe#x�����Ǒԕ����F�ol����G[ �0*��FZЃzӼ�Z�tԤ*�UQ��Ì� f�%Ȧ�� �E��4����*N�I&�� ,�0A����1��c/��Q��"�N�F��л�M �����s�qZ@��|4C�ʊ�$���b.�ފ�����%����Vd�`2҇g��2b#�
>sd�x��$-,����԰@���g8"	Q�ö��hu�V��j��ҋ���و~���&p����-i�0���.ً �٩n�\�ʲ��e����v�ڰ(���&B��s�jǳ��(�"�-��ϖ�D$q"sh�w��k�M�nrp=� h��t��L@�v�����QnX����z���������!�H��νA>��?��+��鈐���.���/<�gڽhEx��C��K��@��7h�MRd-Rw��K�@���y �5�-m�ߴ1�3�(�O��K���1б���2wkb%��Lqv�C�Nu��-��׮/����!����(�K=Q�\�B/��p�a��V˃~�2��6si0K�y��O��Qxlf��T�ENsP<Q	���!�a�Jn���ދ�YJ��=���J�B"]a�Ej��y7�T� (����~��v��SK�{}ʳ����dw1r��+����Mt#�i2�qi��Vx��=�^���g쇙�����A|e���%q;��A0ۇ:�2ra���ې���U���;�����U��P���<���ѵ��E5{v �I��D��(|ˬQ��n�Ҡ���Q��1�ͮ��
`�^���}�;���(�qK�@��t*��k����+�t�v����!ҧ)Ew"i���E��E������`L�u<�S���&	��[v�'�LO��ג{S��6 $V�Y���d���g����S;±	��ÿ��9xn�+�0��l=��6҇P�&���@�0#������GrDػ2��8���w�[�0�������H��O�,R�9IY�s�w��~�j��0��׌�T�z��n�N���R٘�w��{q��
�p6��	�(g�\�Ģxv����z��v�����3Sp��f�ѪЇk��E�e�v`���1�şzok��@<R��2��ik����_���T؈�L����Q�|2������h%86�����B�e��e0���A�UG#qU>c�>6&�b��ϔ�T��L��n�>7ބ�ŘH��=�|q���lQ`�WQ���<�4����o�uv�^���+a��ʨ�`�v=Q|�EO`,��ʤ@;��ưp���s���B��>>�<{q��Jf�ɐ���.k����Vߛ�Wg���l"��Ua\��44v;(մ��6cy��SJ.
��٪����SAaQK�Ċys���G����܃�i�+���6Ԯn��83�b���>-������Ά�1��_h���͋���g��eU�i��E�v���KIp*�APC�CRD�֬����g�W�!Al��|���4S�s�'5"`�>754�i׷O�"#z�t��eXJ7��e5Q[ 	JM|t��~�q$d8��&,e�5T���}�0�H��?����;�$�~�I	�~��^=Flw.*~��x�k 0��(�hIˊ��m��"�����E�[��a��Q�h�`����[�3aI���P0j�t_{Bi�|�̓mRpc�%5�SKg`�A��[���\4��@��Y�kT�4f���ސ�v�d^]mc��Ԑ3h~�s(�ɏ\\Wydm��r¯@l&��%9�Q��*�:߮�P�G����J��9� &����w�g�P���$ 0�F��b�w^'�ǀ�(��見�U��J���u[2P���Ȇ�Z{J $����U޿����\�[��G� ��RF(����:Qc��#����˵�q9}u�&���Ktf�'h�I���&��*p�a]�� �,�̡���/U�v�m�6��7,�TQ�E�ƣ�}��@{��d6@f.�ZQt�?���h���b�؜JU�I��C�{6��?�ʚh��{����_�����i�|��֭�3=��Zb���~sWF��:��"%1�ܬtv�[aA�t�^�SH}��N>����p��|��sl�t�b��q�D�`U���^�/��?&t��9z���*9{a�E�Vz�\J�J�xB"��]E	��~���Í���MP������H�O@m����9�X�h�z�49���Љ�
�Q�1Ů�ck��[�?�݌i�)�ʲ����1%�`~���5� ,r%j�y����2L�m�
{����z9q�h��_�Oi�	�]��
�����TS�ϒoo+��Kw��W��i��q�Eh�m�|����~Ŵ��
��]����#���#�4�i�O�i�C�}���S���}���CKU]�b���X��ӸL=[�w���d�Z�4J�|[C(�e�!m|KP%�1�+�z�Æ�=xU���`0j�=q���^������TR�#�Z$���\�؊W�@ǋUs9��
�?,��)(���-,BǚM�B��g� Wa~=ĥ+הY����u�y^�~�hf�ĺn{{4U+6��s��vN��H���#Þ��W�Ń&-^𾑧Y���*���Z�DƱ�+���#��[�#�,o����
OG<� �&�S}���r2�0�Tzk��W{�9�_�q%6�O��%S�0���CX=�"����LL��1���d��R&�D	�Q�4�A]����)5
D�X�|ݷ-Wo���<�է�@4�K&���z���h�T :0W.m@Ʃ2�b�9�����8Q��0�\6��P;`�����Y���~���ewsO���f�lԙ@	�%�L����77w�Pq�(���7?��2��ίgV(ڴ�D��ȟ��Y�ʏ�ڴ�J�m�ʃnF���i�vP�ٮ �;��Zi��8�vK(�hD��B�~Qz������*C�����%����יʀ��%����Zq�;5ft��A� ��Ÿ	~�(������=�?\��i�i���Q)`�0�.�_�#Z᮷/��L����f	x"�����v�����!}S۪8D��~�o�.i��/�R`/�ĳ)�������6
�φ�D�~�K����Sӳ���W6�yLE �7h>MgJ�)��J?�Nu\����J�C��nb��/�n����S �
�9�IߌVມK�F��O߾�X.�r\�ʸ���3g8d��#P��,ƹKm��.���ٜ��c��S�"�Ǌ,{��t<ߏ���B�l�bv�R���������`�KZ��7��n?o��u��vm�J�ݱ^�jη㤵^�#ᮁ�@���4����ɶ�Af�#�^���2�������c��WQU쥃�X��h���D/��U/�ˣ_�u�y���AK�^�`n"^C�n@��"�a�^*![܊���n��M시|Ѽk����A�]��ɵ%��jl�{�sa%���_�P��J�B:&���^Ҏ0�F-k�⿢�[��v��o�I�m"Ǩ4�R}��n�'0pX:���>�5�=t;��#w���rڏ)��Lk�iEX�ުI>�����uK|"��z	��n�!�F��JzÒ �)$o��F\�,\^���2NO���d����R�G�|u�b�>�Y���u�����9���-�5�u	T3�� �Q	�I�/�6���R'#��N?���ٱ�e=	2��W��Æo@A&"k	ƭ��.�h�M�r�T�1�AطG�[�X�=��<�j�;aǽ�7MS/[���H�g:A�ٹ/�7����G��`?�Ð{���	s�)�|G�NVY��\��f�1ml�,�4��3.����u��t��sS�����XH�Јw��z�t��ʷ��)Hnmv�����,��ʯHT����9$�Z��l�6�����e�k��y�f�=�`f��&S�O-���w�8R���};���徿AKѵˊ�^��{!���2]��Bʙ$r��24c�.j�a�9{���I�k٤Į�=VU4Sv��2��"[B��`%��A�-2�j����g��Fk�(:%}�����\�'`yYA$�F���HPFI+î��X���������\+�6Q���(��>���p�, �[yK�rٿB���/�ޕA�^:t!��ҚgW!v=[m��ΥㆍDҭ�K��C�B����i.w?]f|A�R�x{lح[v��ͽ����Ff�g*�
�U1��826T)���ޤ+f��+H�(����EC��yK����0�%� �uw>��rƼ�qV�g]�~ḣy~JL���(n����G�O�D:\\�I�_�EFb��������K�C��Ԭ�P�;a݋r|�tV<j��/�k�
V�cg�L�ہxEB�;.��B�-�iܵx��0g�E��V%�;%l W�Mb��^����K]�2�k���В�	O s� (�+��4�-*�#�r�\���\b*cV�x݇?��O �TiMUqc''+����lnfa�2�a�s�G�N��f���/&����f�U�-��[��7��%�ʴ+�sp�YGՓ
EK�z�y�w	�5 �,�(��*�l2��M� D
 ��(S��姻&�3�5�͹5P_Mu2�������'C�c�
�9������7>�R|�,q�XB~T�c��7!W;�(%�F�.Tj �w����1v(:v��8�E7-4���F�i�
�X��DW[A��&��&�@�%g7=��TX�����z�1�B)��C�77Co�7���cp�{�r*��wJ����â�.�zz���{��Pa�,�F��%��0�o�zyEk�[���P��zZ������r�����vw��i ߩ�М$ij%W��Y1;���3��!{�<��S�M�]5��{M"k��e���3�G\����H@��L���);r����־RrZ�h�������o�P�,���|Wj?�/�i�ʄ�T�*��~�+do"-'#�����5QR�N��K~�켩�pG�GM~��Rd�7&�C�"�����q�q>A���T(F�wZȺuĶ`nK���]h�*`��K�lƈ�"5���4 "5��f��A����܈�H��T2�yҏMn�șLW,��ʪ3ɟD7ր�R!H���Z��D��>ͮ9�}��-3��J��%Jwq���D���yuu�����`�ZքC�"�\�[���@���}�=�J�> C�{r8i�V:ZZ��G&��/����	�J��Ԍ�&�xx�:���luI-�Nn͢��HZ���#��쳧�q4;лK�ӵ��ntas�c_��Y��jˮ�E�h>�e��1�y�E�S���1q����}���o^ize����Ŀ�	�����I��Rٺ�^*~I�.�Je��&�t�Sp�mڂ���}��л�������T^�-����Ŷ�w̺�9��#���M���3$�
nSkNaU�'�1�<w�}���[����P��Q1@�G�k]P�/m)<"X�_*���w�@��A��(��&�$=&�?�Ī���[.z��<K����]�f�a�|�'��O٢9&��$��U�����E���>O/)׼��mPq��}�S����v}b=?R�[��Xb��,^��N��m�Q�cCd��
�lf�m���$lI�&���w+Q1QdB!GD��̞�7��y�Z& $c4�_}*z����3u��E����B�8>N}�Eʷm�-��<��)�sٴx�n�i�E޵Ad>/��MW��J�6T�}U~��dh(������^������G�ʃ�Uu�6�蘂�naT��s)aѤgH�Mob��>[5{ڢ���Ѐ���þ��v?��N��5��Jr{[x%�@��Q��Ǳ��&{ܘ"GrJx�l��N�v�q�i?���j�oh�|z���� ��.G�����5��YI��e~��P�6j�Џ�?���	�'t�ZB$yͪ�.xq���S��(-�|�Ð�ߩ���՟��K4�E̞��Ⱥ��-���Tv��gݨgd���a"�/����a���
ԩ����l�p�ҝ6�#Wz3>��z��+��>Uu�6Y˅2�Vk���$�����s����ҷ���&�3��|�n)�|�Ǝ1E��(˔# �&��l���{!��JKP��Uv��L�������'��n�h?khz�m���Ɋ�񛉒�����#�AJ���O�)�u4�R��`�m&]�	��i�c�h�;��=\�Q�L��P�R{t��]1�3�^�~x��؉l�)mw�ܚMف�\�CrF�	��M��P���.��C}F�0��ę���2��J�Zr�����܄���#I2o�L}�Y����?�0o<��R��Y��N���}6{�� ;����d/;���2Qg{>�`B�rfwL�ݮQ�����k�%H��/
*-A�|!�i�&�����nVB�<g�֐x�@
��<
c�Fo������;�%���?[�̔ҿkl��M.�w�a�� UE����7̙�{�W�i�l��p�0�G��5	B���j%Y�3��\��4�וC�4{�9Z�rN�ϧC�
y]T0-�$�� �=�@(y�C���0��ix�!+|�|>}9S��~_�n#�;\K{����p�?��L����ڰ�K���]�&�˺��(#I�K1\8�yC�M���H���@>N�̑��e� �P2'y������I;�4i���?���?��悉�W2�r5�
�)+�t�<Ί3�DE��4�,�俼K.j�PJir�+���:��K�$Ħ�/�2�����+ԲbV��g�6�������hDؔb��F!X4��KE���HX��|6��DW?�k�E�]�Nbp���HsMq����M護q�OP�g��m�|,9Y
n��q�D䧋 y��*��ۀ񍸅)@0ֳ�1jC,�������W�#8���t�R�)�Qj��7����>�?;�NBC������iz�qR��g�->�[Oa'���k��z�!�m���N�l�4+vuH�bcț��Y��hv)�����I3�z��4�E_�Y������Y;�k����rD�ڮ����;y�uCh��
}gK��QW�^ @�	嗥�H�q�
�n�����v�Ԋ�^bc�Y���b�d����h��ȥ !�=�"�I�ʶ�K�Z��H?*rxt���D7��������/�b&H�<��X�
��B��#E8�]�I 1f�S�'�6|��H���;Ɇ�ĔY���[:6��qE�,�p�O]��S{��Q�$�hg:9�*Br�(i-ꐚJS�o_b埓ȶc�����zg~p?+�v���]`��Û�ɦ䝃}���|�ޣ���B�&*H�\lnގ{v�����\�D�}�]7���0t72�I;��,�s�N~����;��,���N������-y�۞�[�aoγ =�M+���;&j��cs����<�0���.~ȃ� #��{I��}�Wv���Tz�>)�6�h�0�rִ>��u�i"�1iׂy��ȝ�j�W۸b�Vgӑ�Bu�=�j�;�h�I�)���p��E�{��#ti8�&����F����gޯ6�Tv?�i��~c8�.y3z����(��h�.�zǏveK���{g��L�	~��V���@� �t�VCNv�^�iM�sh���8,��]x�y�� o��3�X�̺���R�/0p�� b#0I��<����e������FO�"ۇ��`���?}�ppd���Jb�*�`��謗P\�ۥ�i�^��)�� c%<�8��\���$���ظ�ި�%�?�������'h�Uw2�N��V?����<	�B>���(@�0	dM/mN����}���7CJ���L�1TT^�#&w���V�'}����?�q8��rP8�I�so������P�]!��q��Z�NY�œ*Od��6�|���v��QCi OPj���1Zu��ǲ��s
�چ�r��]�1(��?t1�X!�Q�S�5�&M����V#��*�V<�*z�ϚVI��vP�E�,��6m���d�_S6�ZpKT�2/ol�T��U��W�?���mm���,��W!vΈ�^�q�r��a��-�����f�_e�s\V������:I��TaK�a�R�&}���N/;�@�6U2P���9�P�0c���d�B%���p��ǜ&��T�"1�"�O�A�-j�/��x����oy� �.�k�*���
�|�AKIX�x�!��+�(�������hv0�Be�����+@裭"��vW��� 0vTN�ֈ
|!��E$�Vs�1'�P�^�oS�4�D@f����n�������ͻT��ei+	eb"!P0o�1Z�M!���	�$fvN�Rrm���b��\�7�u�Ld���x�%�h ڕ�N��o���JM�u��FgG�l#�z����c6���P=� ���9e:$������CE�Ψ̌��u]�J� �O�^^�%Ǯ�Y��Ӡ 4�6��6��1	�$3пǏ����IF@'�:?�{�箂�e�p�#�^�Q��=���+7ϭ��<{R1�2���\A�?2��~�B(�Ăn��2XpJ�i���ix���G~�o���t<0F1s��ǘ�NL#M�<\����������$��=\�#�ٹ�&� ��S(��T�����:��¦D~�+d��Z����9���O|��}�������'��M�F�G��1q�r�Eě�D�����Qa!�'zHH8z�C����!�����3c�4&�~$�x��G��)��FT�Ȯs��ຖ�Ha^�O1Vcn�pt����;z�C'��M(�^�F�I�%-;ڱ���v�ixq�s�cd�ƪ�~!�c%k���e�&��X�`քօ/:�4�+nͅ����}���ڑ�<!��y��3�!=���Sl���K��;� 
��;om.�ex�z���mq���j�X����j����)����Z.F��5�1������5�>N;Uޅ�t# e{���'�Uj���&�
���9?�F��'gT\[��F���؀%���}R-���(.���;��2����de4Z/�[�նrV5���zkv��6�<�A��=�ˎ�3d4
S����7�V!g�͎�g���@��d���.��j��J��G�����ki�+��~x;t�k�E"���e	³�h��
���ڈu#9t�ndۗ���Z&z��<��$����M$���F�&��&ȴ�^�d��%`�>����C�W}���
v��� ��·�0��C�.yM���R'2D����
������S��um0P�u�$"�a���,ݒeu�?����G��;�T-_n|�M!ٻ�Fp@	�1�&h&�!�dp�\W J@���'�5���eQF~��D�a����ܐ��ǋ����xʰ����"��M����e�����͝Y|�0K��� _�C�t7%n��J(�W[��g�U�!]�v����t��=w�<�mæ>��CY�PD9·��v���ؐ�QP�OYso��cx��f!��i�:�r�c����LH���֥ <"����0+񙰚�T{h������9�7J�y�0���nq{����<'�D�*5@m^6��{�ؾ��gy&�G���K��JIy�IoE7���>����\�@���Zt���h n���O��H�Ot}�Qm�;G�Ԧ t�b���c�Sc�z�Sv9��!��4�Q<���C�e��8�Q��-�2�A�ڳ8��am$�ț�|�x4i���}*��,��|ӾX�=x@�@`{�GE����-�wj���&L�+t)}&/�7)z��}/ſ=��~n�D�!�Բ?���һx`KE ���~�k��a=�`4+�9ff?٩��WU�糨ܾ��Q��M
i>�I�Q�h�ଢ���3���@AwU�y��F�Ѽ`|��w��Wt) �(���9c����>Qv!}��~`P2�܆���b����T��}���g��b%�A�/Z�ݷ
����C�� >Myp��c���`�@���v^�S�"ңB�-�9����r�Ӊy}<����� >�4��E�8<���sd����(y�#���!��Y��e�����A��MGp:���P&�!�t�ۓ�
\�����7�`�ԥK�f�ěr�4K�y簺���7{�Ww���ec��D��n��쿤�^��e4��3TÈd�����YT�^C�!���jGMZ/��� �@iY�r<�}�xB�XO��9�1ei���!j��$	Up6�0\>D���-��L��T�#��b�O_��[�e�s6^YI�k�:PZ��j�Dj������<��"�����ŧ�/PuK�kIW"�iϴ�GP�[�Bg*�&G�v�]�)�۞�7<�bG���s��qg<�O�������g`9m����C
^��)��֑_�c�=�	D,��t8AqYm��OQ��R,�M�O�k�/������[H� 艊n�X�� �^��\���q�P�{�)6���yc���Τ�S1��\�G!L�Oȷ�fO�;���&���s�[���i�!��6���$���ȴCX�u�T�8f���,�.���"��EZ'-@�@�:�a�k���I�䇴�od4����ggԭ����$��M��:bg�pγ.^ZF��ekZ��o�'3�5����}�P%Q<�Mj[n�z�ǅ�����W����y�����w�!�S����Hd�0%���G8�����?��'��k�����Smd!�s�䪈��Q�U�k䅏'�*)�>B�*�\�!�D��װ��U�+��D���Jů蟌_r`�É�[.
e[�V+3x w�}[LϤ����O����d����͝0%^�R�(��tT���R�7���`����^�;��D�d��<�h�l1��[AL]�3��g��l�Pj��93���0�`[��1�"����<�);+	^�Ȉc<�V�繖��j?����W[Kuo��Gp��'e��AZU�������t�9s7p�c6֟?=s� ���F�f�ȷ�r�E��o��j������bϴ/o�]��F���	�IVԇΆ�Tx��u+GN^ۗ���ջ�擹_�SH�nn�G���Y*�1'�D�F��/�����gZ�`�>O���.�~�
�c��êk1�2E\dʾ�Z&��z�tICPt�%�������ZڥŐ�C!F
�əyB!�56��R���]���t��%��L��8l�
Gy.����b��,"Ы�B�{��~<C����Vb7���f��f������YYf��t�(�~V�{�̃�G�1�G�B;���EH-��Pn��*���C�C6������(O�����JA�F���m�)�]}~d��>�z8��8�1\ʳ�1:�� (O��z�:��%���Š�T���u��
K�W�x�rU���#{�d��R1��k[�J�Qhg�B��#�w\��ந�@7�i�k�*jF����!���jT�G�5������;Nݩ
�!۴�C&wQ��B} Z��n�Qa`�.Q���ɰ7� �zޚ�U�����&׸�@�� �°���ތ�zv�Dԣa�|w��U�$Xi���<4�5ʺ����W�ؼl2pB 8��L��@�X�o���S{z?f���9�H�(嘦9^�8���i^���٥@��i�cs�X�WJ�ꓫɋˁ���5P���F"}2 b�~ؿ��G��J�k�g#�Q�������EZuU�,x���a6Y��p:�Zǚu�j.� r�;�ɡ8�ݜӾ���E���Gr�5���٩ޥ����ν5�'/v�|+B���_��]'d��{-_p�][�.@���#��Bč��?'��K��p�YJ��	������3���' ���n
�-��60�����DS�l�-4�"��)�-��ϵB]��d�)B���c���,�odͺw�z*G�Ɵ�c"�|�h��{,��q� UUy��)�Ǵ\�c���em(��ٹ�nӍ�z����-&۫l��2j-ҽW��t�L;[����ߴf���L�85��#
�ڜ�6\���T-糯�h��}��F����:�E���?��O@���m6y3���:̍��ט�\��Е�7�`-��d=|�*��n"n}E��q���v��0Y{_��J:��2���viQ�舘�l�g;�>����ʕ}x��H��W��eV��ӾRO��c �1�H?�!�Ύc%�wP(r�����UŇ|��H�;΢�����%�#aܥ����c�p��<), A����Q��N�(��H ����!,z�p2�+��W��)p��5�uF��3�� Ҽ�t�u�xr;�����x��f�ʃ���m�`�
�@�G���Q�N�簈� m����]�1ۂ��Ce��D��/��߇�R7���:���e�*/@RBσ��$΄�[��K0y�OI���{�j1}b{� L>_�i�s��~.��$� �����c�
���Ů ���v�V~(��BNe��IS��8|(
�#|cKv�L%�1�&b���~�y�\�xM�[�vP��!5�	]���O#G3?b�aS(���-�1�v
�B�`�s���y۲�������~�j�:(�Ƀ�0��[&<�S�Z��	���B�;�x?��̮yXC	���^���a%8��m����hcp����lnUouDY{�-|/BG\��W`�ʏ���LG��kL���	ߞi�8��Be!��������`���=Dor����G�-2�lg �T�J�%?z6�y���s�h��|��X�Q���Q���뺠��:gt� wA)�ϩY�xҢ-L�q��2=3���Ì��i^:O��%��܃��ѝ&�S�R�Gu1\�<<?�-]�-�V9rP+�]�����#ǣ�p9;�M�â6I�4�i2^�C�)��/���8OĈ}��P���>ף�ޡ^ԣ�������~$4�!(t0�$��������o}�8��0�^E�y����h��Q�\8&01,��/��8�J�M��4 g�i��?)��W6�獳�+-�<����8D�-�������99�y�������z����_���?X�&�-��Yd����\K|�{����5��Yܥ*N�6�J8����U�A��Z�@�������}.�;^H�·f�@��6~��V��a�v��g�Y�l��XX5����1�O|����L����^Yz)�f)�a��}[xq�\��ѷ�L���/�_��<��eT�q��3E_��-X�*�Ԕ&��Qm��ua�8Hf(���r{t�Niɹ��O�$.WSi��ۖ�gT��&�/b�F!�܋�~�����J��$T'�Ap�'ܗ_���	%j�����h)�'!]6ί9�"#����LB_P 'ίv[�0��Qqd°�26�i2^���D�����(�_P_U.^��Q�yR��FDm W'�t�V�%QV lI3�����s�n�����4�� ��*�ی��=���פ�ߝ��	Zq���|@|Ln�/F�X�2��D�5Wau���z����Se�gTM7�x�ܝ�n��4)G����R��U��7���Ǉ1�:k]���4�Bכ7��A��˺�VjT�(d�V��dv3yuvwy~\�Ӎ}W���ۚ��HH�D5n�;�|lD`�i���,�ᛛ|P����M���0�@)���,:Q��,I۫�Mu�ͱ����ڇS��:�m:+f�)$�o;%�&�=��!.S>��Rُ��C�b({|QW��Yɪl���ӫ����]�l��į��Ӛz�"+x�����#c`O[�Ls�W@C�D;��%�:9�Ev��E��KNG��Rp΋3@|�@��p�\~Cfb����{�?�<�u������C�ò��������"be�5���k�ǡ���po�E	�����4��'�Uڿ�䀄q��'�E��i�@*
�P��%�0� )ֽ�i��~1hV�+ơ($Ľ�=˷9OeX�HL�x8I��t����Y�E�_s}l�q�j5ω���N�\zK���z�� U�i�6��2����Q2p\g�_��.������=�8y��/��	�i�Q{YeP�ѓ�}Q|q�i�ԅ�t;�h��ҥ�?���=w&�U�[��	;�5������qH���%�a�H����_��צ�n
`�[��}LY�%1"���Oo�"R��+;0��Y�B�7�h�<�|{i��7�}��Q��ィ�D}����X�i�ߖ��(��E�������	���l����� H��1�??/� �i�U��i��?Z� ��u���?Y��y����A�bϕ]G]h��`-�U�n�13�uxϑ�ڱ���Ĕ�l��ޯ	�_�F@��DR���|�l�L�ZA>�h��k���ʷW��`��:o+z�+rE8ij����dCK��L�Ė�u6�;!T ��_�Yʽ1�x0����l��"%P��`��E��q:��6�с�B�H�Y�qmeW���ڙ����E$�4��S	7��������R�|D5%I���~��Iy����2�3&`�����g�k�Q������t�?*���Ȟ���(�������evR@_����+7{�Wcj�����)`h�� �	y��P M�?u��B�3t��9��cV)�ˋ,
3^!�<h���Z��k���l���+"	~�21�$���f;��@�:qʵ{�2t�f���.ڥ�eھ���X6��K��������r)񷼫��v��8�4��0�0AW��l@MF�eh���������!`���:pJT����GM���|[��e��
�o	�ڔ���@K�y�+������5���Z�-���
fs�{����䭾��0X]�N�F�q�<�B�QM`c��Nv�eF��bm�J!�U��'w���������7���'b~��!�N�@�h��Fe�>�~��1/c����a`�_s��j����T@�Bl���8�^_�%�/%Hqj1ekP�'R}mQ��"Y���#�~�}��}q�K��$Fj�F_�����߁���N���`�����E����j��lE~sqa��em\�8)��bǥ1�� ��Iߐ+��ھ��պ|�2��9ߠɘn���jیj >�V]o#Vµ���OE���=� �bY*i����TI�Os�Eq�H��t"!+��r�4D��qؒ4��jM��<5z�wu0�����y�w[��X�O�u`�vӄ�j�;*1��ȧ�t���ݪQ�:��
�h�66q��\j�ܟ�m���gR��n��|��2ۏt��(�����q��@#Ѡ`���/�N��O�&�K�<��O�TR����raw�TV�U�-m�~�/�7��J�.N���i:֑~�`m���s*}����v�����_�+�~�:8��J��:M�#�/�*��	��D[��~J<�Ѱ�(v�a�&	*r��%�K�ܨ���ĺD|�\P��6����4ˏ�O�H��Sk�\3J,]���Mݟ�z	:N~}�0$5Q6��zQRH8��@�x���hid��s/�WF̧�7�\�]i�EG����:~���	[�T�&hj��>��&��ZA�j{�n���	�&*���sW�2a�r�V<U��[��xK
�D��k��]f�Ot�t	�'w�qɊ@�\B,J�:h0gu��XXh����}3;$��?[U�3��/M�1{96:#L5Y�ni]�~��c�p�d�2���A1d��3�^��.H�y�{$��n���5C;@$�ɐ����ȳ����Cp�R����ohܘ�k�GB��8G��[|P1��s�\X�h�����E��d�G�\�{�gg��h8Azד$�J�Ce �9}}��~A� n���aʑʟ~�p���ehEd��K�o��z/!�ɮ:g$���뉪7UQ�EC3�e!���Z��l`<E��#R����y��I��w3w���lW���h?۔>��?�Cl�����'�x�(���YWKH����^ �(6�1n����J�uG7Z�
x,Xآ���n�v4A�N��ā�Ky-��~�%���ٜ�	)^{�.�_���^$�{|�n>G��� ��	L`�>3"�@\wݹ&�8␄�ƿR�5�X�?E���w��G���B�pn&��=޲��i��M	�-ǧˎu�8�$5p�%�K�q�A���&���X��m�4G�W��0tf|k[
����(G�h�|��z��|)�"'�'{����0�"�T�s=���#1n���VGv��
����m?8���4�����j�4m�o��y�b!Bp�[p��I*Z"N.;���!�^r�k'�Ȟȋ�ML��%���ˢu��1���y�S<�9x�r�੼o7v���b}�EN�Ka��
�羴Y�R�Q��ǟ�[�^k��#o�U!Z�2��bά�{VU���O.�b��	Y�48;XA�k{y�xL"����BH�
�#x3�ri�m�!Bܰ�8�KV�	�b����%|����`%nV���d���6�w)$�A�>���HF'��}ًE�BuV��4rȭ!����>��O�|x-���Ȋ�OK&��ߕ��P�0s�#�)���P��"��bc�rͩ8��F�)��r7���2��8�"�����ȷS'�4,N����j;�w��fQT;X�/�[�i;�l/3��uXB��{��6���O1��F���_��b�����ݜ�y� `�M7CDM(�_��w�B�����*p��.�6�]�Q�%����%5�;��[O�dF�����6Q�1�˱
nӦ$�U�.$��w�Ձ.G�Y��o������4�#fJ�J�z�]�Db�iƥe���Eo5
�F+Y���6ȝh��r5j���P5�n������Ϟ�H�r���N;��֚`�O�p�Źۛ�7^�R��@k8���\��*�kM�$	tkg��9K{�8������S�ھ�!ug�n����q �w.uA�4^�����T�Š6�C灡�sܳ�g?����Kg-�>�IB>s����}�H����^`�L�MW.t�U����W�(�~�hG$�"4�Z6��*���� #�SA��l���+/VdQĩ�	i�
Q���$��棼3�if������O���Q�4����ܾ�!�Rړ�!��M�����^��ک�v\
*�-����_�]ir�%d�}�����*����FWm�ӹ$�M�"ꌍ$�Q���fp�V5�_Z��w�Rn]�vR��_�(��Ƙ�m.%>JS�_��h�~Q����>E8����z�i�9��&k�[�mYkH�S��	��SiГ�1�=A|����[��	���XU����%mP��>Qs%�0��Ş���� ��3��e���/�ŝ"`�-H���}U�ޗz,�CZ�a�۫�z�+�m4� �(e
q�~2	�&��c�P�c�&�Uw`+�[4:Kvb��%C���T����e���º��gH�s�hc-��}�8�����t%�Ӣ���GNk1��K��ռ��@@����Nl�-q�I�z���HP6g#N[��4�? m�^�*�6m�@Ԇ��1�cr�K���ЮT�jg�Ǐ����I0���j�//���e�o؟o��w3+x��p2�#��}����4R�2��7�v��"h���C�W�TL�,�Bkx:��9n����ㄞ��+�� UR^BQ�dUC�ZA�E'�Y��e9tj��������3��-"�P^� < �d��D��q�4|���  l?�.$kW,k�O)ų����ֽTl�����g�����|X+@�	����Ls�.����%n@��E�U���ú�g �E���w-T�F<�9�bh;_�x�>�.�A��bƝh=#m�p�t,~'j��I�����\���X[٨�Ĩ��(H�^��� ��%�.�Z����.��i��X��9&��0���t��em���?o���Blgj��Q�#�ʻ���)X�m�&Lq�x�M�ur�[{]#��j=D���8����sj��^��K�B�fG��4Qϙq�s��2GA�vT<϶��ߺ��z�gsZ�S�z��&���]�97 �Hjf�_������s>���Ŋ�f';��tI��:"�]*�QZ$?��<�Of\}��U�v)r��a�68>I3h��E@a�ʹ��a�孨��F`7˴���Q�B�f3�sf�!O�����H&��c)�K��&��t[�<��B��{�V)�N�����y��"�4��,�2� �8����a�3쁸v��$���?������6�,��!��O�D}����wadNXk�3_K3K9�H#(]��G�M�������3�tm���x��[:w���o��FKg�Ru��*t�� ��x��\��A��������;v�������?��(oU�F�d����h�r���u��@E�Z�0�3X�?h#�K����?3z�А8k�� $�+�F�� b��>����tNE!�e[�8h ,xK��!T"n0��Ev�r��9_Ix��0��`b*UKL�eu���?dDQ�,�:E0���X|��d��:P��j^C�p9�I��,
{���5`��?8z5�
H|,�#�ڞ�����`9�L��OBl��pV�o;��'Q�D�����������!�~n2�����m3V
�7""�~�p���������\�-�e�(�\؟�?����ט��D=� �9o�-�1�=II�0mƿÇ����SU>LΫ��;Ȏ����8x �Q"E����sO���q	���Y�=��^n~�4!O#Y�H!Y�ɸꚞ<xrK�	�x5G�P�5�u�7�j�j���DN%`��|���������
�+k,s�ٖ�7O��>��, ��*,w���T^�5��*��bVO����vO-�<�yE������Y |}خ�b�(����U5����m�
*&�$�����*K�m^[���#�8 bF����*�s)tYAF�����Rڽ7pC����(<���{,����8�"xƣ�%�z���[I�#z�Zp"�e�=��[�hS}t�3��})�}�MԻ}����_�9h��Nw��������2}�{�Ǯ��|�S�� ��X9�i��Z�z���c�mgH,]���X8����N�_��!v����X�"&����U*� �b��`�j0�9�$����(��9���:��ت~ ��t�I��I��+e sW��óF���R�ZDw���kP,��Ka��4��w�Ő�I%ld`�����v�Yթ;p�O���n�_"=*�v;t�Z��I�����.UH;f.�$q���W����ܖR��>��X#GX�(G�J�P���q6dϹA�
2C��S���KQ�9����,[��� `��8 *iS��@	�H�Y��]�rD�&D��	[�VGI���J���w�ߘ�($�:�Q^�S��"?����C)��ɛX�2����)�F��ߥ�z'�6��Me�r��_Y7it���a����N(���?�R��"c�>��_�&j�637_����C��i�ꖬb��.1��Y��$����l�,�BƠ�F���:�T�'�	��ΌϏ	*�*��L8C����J�{)�Ծ��N}$J��D� ���'��g�H!/|��$�ٰ��&�B����1�e�oS�_�� ��U� "T�I�>)!���4WI�����^L���P�����P�9��+.�	l��(���D���H+������Y�gǃD�|}�G�WzGsf��D�U����+dyZM*N�-�L͟�U̑�Gș���I�L6�T�a`��� ,-;��0~~,�w?|du1.U�rzz7sN�/��I�� �=���1H�أָ�7@c�ma]1Ľu�t�b2���&��@��t5�烁��"��G���ەtP�뭟�@�;�R����G�u�*Si=�2�ʭsUS�|J��B�u��m�T���uQ�j��s����0
�^��\`M���Ih���-�`]Z�\L=P�&�sӫb{�%�Bz�B�%�Af�op̊L!�a�,R���o�1PHFG���d��°���=T�sX�?s�_:؎�qU�+�h��{/o�\^����޻Z�� �B�&Q�7�e�_�@I�Xߦ���{}����.��D�� CW��t�$���k`��R�gǉ����ݺ� *"=W�3(���pu�F��1$^΂��c�LB�`ּ�Qӟ�cU���$�}T���_���t6����̊hxy5$�mm"��A2�M[lY-4�B��C�2Y�Pqh��w��tC���C����/�"6�=G�[\���B<��Ҕ��0VMB�z���h�B��=�p���J����-��k��t)����_����>9)��,_�;1�dw�7���D�_J��F�ד��҃KSZ^]��-|���ǨL��t�-Q��ޞ\��,�'��lx��\IdK��1�޲5crۣ�q�"�D�YGf���>�#�����
�]w�.>�p{*��Œ͔���}��0�{��A�d�лK�i�����-i����5��	1��=�����g�A7���ė�Ӥ���xx�5,�:o������<��J	�-#���5��*���x p#	���A]'���H-6uP��Y�|jwU?��͵Z��v\����x�j� v�l����(�Rĩ.b8=���e��[��<`t������5M�x��~)�H=`K�88W��%�dU��Y4K����1+QV�Pu�Ӧc��'�L~/��'O�@�?C�0v���b��M�˵J�/��L�5UY�Ik#���sT��B��Fϛ7���g��3�cO�a3���TG�I�Hz!�N3m�c`f��40�:�8�������R�9x�1~d5��	�hP�|��6c~�AT>m5�%�4����#2�V�Cz����k �[�:�T�Η�b3�I�25Z�sE��Q����*.Xa�P�� G��W.���?cG�j⥣Z�,Tj�$���k�K3���Sv\��<-��`<�<������)K
�`Bc��(�e�i�d"�MGB.��ԢU�����<v�`����Γ�6����n��G�g?+��8S�E��:���Zq1�)P΢K��-8��*.�e���O���jB���!v{t�s�|~��7N���7bЛ7��w����1]uf���P�O�'Y%SXɸv;��?�zs�ҭ2�|�h���Z�!�������%�9"P��KVZ�>On�_X3��"�t��V`���jjz�^��cҥ��NE���/ü��~M�p����Dd��hWΙ~[��{��D�EGs:��k"ĬPf��: ��%'���a�2�b��ݑ��~��$��9�e�E0]�r��"=��C�_��}���ଡ଼,��z{(P�L[=@@�V��6"v��P�*FIk|W��Æ=�|�G��*ᛔu�	;���m���뤹��̦�����邹HOH�Rs��`<%JX,�D=^�x~uA��X$���6�E�w���RI�a��ݸ��/�[	]uԧ֙���Gr�.�I�ک�l�M��X��ɨ��|��	��Y���8��A%�ݗ���qý��V��$����m�����)�X󉳱T����&�=Y`�����`����L-�S�v�Vo>\��vi��$��_�����4����D(�)��S.�M� 3_�_[]������M@��Y�/,���L�Bw�&�D@�٫q���g�ozD�J���e!2��07��/O�����1�{���g����|
���=cA�u�JG�|�r@�����Jo--�Q_���$�Չ�^l�/5���d!�md��$�^{�B�����,B'�HH�:┛ߤ�b�ϥS:�NO�|��$˼�E)�����4J<�YE<��lb� �g}�O
��j�AU���%��ʅ	��LzE�OG����/��9]jެb�4W4��<?�.@|=�����j2m"i,����R��C�nPXX?sp������7�F"�a��K��6��|*��7ym��RΓ��E�B�O����F�8��μ���%zC%�bF�:0�N2R�d�t!���~�)����-X�\N�ozb�B��b�*G������L�bW�t�?!o<r�XR�K\ \Js��b�߯���g�9�Z�(1�A��[�G�:�&'(s{�piɰ�_�܋���EK��@b��:h���	�5��%?}KLAM:{�ۭ����j�)��R���B�s���)?��j�rͺ=oy.��rR�Q�^:�� �B�@tI�)��&��#����6�4J�FlM_��y��ؗ�\9�ß��5b�_�����D��b�*�d"�O9K�~fp�!2�m�U�h8"�2p`[����k���^9V;D>�8�v�+��R��P� �9Ϡ�Ϸ��]Z�ƺk�h�BljL�����K|�C@%(���-u��P
A�Z�l�`N�ys�r��e16����!#�]C��Y�'��4իt0EL*�E�&,Y��Y*y*��ST^��x�����p	�����m��`rJ�y���)xҮ��6wq�+���NzY5��ܲ�9n,�c��s}w��mz5N��f��-�ɒˑ�ƍ�Q�TE��8�]�:E@[b�H��:9���yw����w�t`h������U7_gȱa��-�cLDl��3��X�<}�!.����������t1ì�J�˰c�/4Β��8ac��5V�̞L^�[r1#�j�9�r�����Y"� `�Y�MI�w��:��M|�S,��U��y�X�70�E���2���[JJ$>���Cq��@���u ;�W�X.2��vi�ۆ�}O���=�u���(��>kz�F�۷X���Sv֕���ީ-OB��3�O7��7���!VYq=P�pr0��\͋B��gC�2���3G� .&KZL�C#�ܚ �|�|�̺��r����#4��	�#y2u1[�� 0�e�{Z8��Z@³�UJ���a�O!�q\c���T{B�����S��$N~ݰ/��2�V�i���u���E�A'�� ��.���_������%k�M>�s[F��1^������tO��2�(����)o�U<��~��OL8D��W�{����4ɔ��&�匠)�;�R��E!d�fK�̚xn)`�Cu�g'�1ר��o ���G��!�;\�G��E������|����zi#$�6�7���Y�7��~�FI�fa	�q��-T�;��k9(A˴л�T�<�ֿ_&I��z���,Q��0s#P�y4�XQ���~��i�̏EY<:�ȭ�ӎ�����R#'�c=�#ĮHTe�w۰_֣����f�y5�R:[<��BiP��v=�\��&D�	��ɞ�f�:�s�+�o�$PX�'#4����t2̩�ݸ����m�ɪW�c\w<ku��w����w9.��6��zYc��w��xu�2���G�!�����LnK�Q�Q��R�k����0�h7 ���*�;~�GO��a�����e��BH��
>9D��Ҿ��kgu];뻜��AP��)���)S��E�*G:�����sf��y�3��1��'p��J�ώ��ǻ�=����������9�L/C�������&����
L���3�4��t]ǆ�OSq�f��2bE�RZι�J��� �P6�1��Ж?^?��1GZ˯������j/��LA�0:�6��f�J�/�o��}��Q��7y��n�7�1N�ί�=�\��8un�X��������ȳ����k� ��#�^�}��nunjă�2%�#c�,��U`����x\�������>�1z�[�ō:�ܩ!<��>�X��論ķ��hȖ���|�<�ƪ].?�.��9e�ߣ([?��|��U��a�q�ck��N]�� �!��G:<�� r�AI�8<LK���<��T6:�0$�h��y�֨��ɀ!��K���hH����/L�����h�ә�	�aD����Ƙű��t OBu�W'4�LK^�7����z(E�>�P���S����gE�%;�߬�L�*ԩ*	h��!�Mo2���G�_�^���%��?�l���4xZR�h�>����l�2īSN����۸�(LP_��4K��_c����|>����v��b$-P��1�69�1��B�����k��Sd(>!=����9E��쭎r��A�Q�|8��=��5arަ�b7�5�C�L��
�b�����`����}W���$(����N!zs"�;��7�7�˜&`N�|E,�� �O���]%,��^��	�E��YY,�A�w��o���B���`�H�GQz~��8삨�����)f+*7dg�2��$��֞��-y�9��ı�NG�qՉRO_K�poK�`���h��� 3]��D9��/�y��f�D�����Zg�n��-����h�&G�����G�$K�(�����V
�'C��4�S���񯆏�*��n��I$��U2����@4���͐N?<LY+�������4�CKӎ�7�I�򥲬`w��ₖ�$s��᲍:Q
�ȗw�����{Ѡy@��&O�1pw���!�'��S����&ܞ�OD̀����J�fr�j)�D_�#1´�'�'{C?�֒� ��� 8��<o)u;�f�vS_�����>@�gH��:�Q7��N_�/��1K*���!i��z�o�[|K�"[��w���4��x3dnJK�w�c�	�����ఘ_����C�ڽߴ�_�I��ԗ����[�מ!do7���{��#G��`a����gAډ�R3>�f�z����W��хJ�l���� �
ϡG��i]�hÏ"m�彭���j��=��/�Yg_��e�M��48�!�ѹ�M4�VBR#�]�^P�pu��ɩ3b(��BM%�B���m� �6�H*db�Yc����oMcd����٠7	�:�e�ȡ@,����D�pW���<V��ǿ��Ozr/P�����ς��'�iR0�1+����Z9�C��bd���S�;�)d�aRB��[Ã�ͪ{m��Lzyn�f�Q�e��'n�� $��jtl�2U��榢	��N�8�QI7�`��;�h�-�*�Zw1,�UZN|yA�U����6�<���#�CA�Pٺ��h�����`��#�(��:�W��o�>�����d�i��WM��(e�=���{�I&�WWz�gZ�HhIH�M@��A�'σn	r�d2II�����B�@��L��R70�`qD���׳���e�!MF��������+�A<�d�ɋ�3*� ����p��K_s����'��᮶H�8����+j~���0q[1&I�aKw�u���nU���g1`���;�8�I�{=W����A*t������Juj?�(���5��I���7�C��ĉ�h�K�r
YKs��n�	Bj���h��P3 g��e_f����.,���4�|X�D��k)�U���r��g z�:}q��B)�F 񇏇࣋�G
J�M��rq�Z����M�Iϐ'����P�i�3B^�6�d��@���	�/}$���&�W��ߌ�ZB�����T�9�H�)��
d�x�/�]0ز�����Q���+�X�,���`���Y���:f� ������^��m�ۯL��C�m�7��/�@�@�:��]>�ܮw�J�X�Ue����\��H��u"�	���|�Z�����V5�������(��)O�[��}��@�V�K��4dࠧ�n�t��q�1-]�+���X2v��.��e���mL��k��v�;�}$'B�� �e�g^�yI�	�ɍ�1��t�v�6̨#�u����ǅ��d��$�����,��mK^^2����sD%�q�M��̔��'DVk�|�l��hA����g8H=i�t\X��ۛǟ5��̞��.)˩:(�u���0�͘�-_)z���S~�f��dA�ى�ڕxFy�k+�ldF�_��ziJ��ԃ�[3���U!�m͇�YOb�����ܨ�
t�)S,N�_mƈ<����;(��A��
<���Jy��S�8QZN�0��� !�-��_� 
	Jb�]���0��$�՟̱�JU�9�~���^s����Rfk\�yxb,B��9����y%��,�~�a�5�l\7�/��D�%����z_�v�6�i�?�y���Se����tǯ�'
:���g�l�+` ��cn|-(�Ϛ^��v�����u�d�ɳ�,�"J5H��"�σ$_��i�x5�#�ÖJ}�s�4]S\1�M��4{֨���}�Bf��Z�4*i����W�],�v��i�lSqX:��t�$�O�M��ȭMp�N^�v�*��x�]`��;��Ztu��4%�۫%���"9���N�$�����ҧ��`U�s=n$w>�_���x���1�G���@���Da�q=�v��3;g�!hp��fՖ���ʬX�Ϯ�(M�q�sj��	|��aܔ )񠼱c1A�<�v�ƀ�l?>�E~n�ؙL�,Pd��%��`�G�_.gt�R��#"]��ߘ�uCW.�D�N(f'�gvqp�&�S޴����1����gu�3P�L}Hk!)ؚ{f<tV7�'��p���.kٙ��c ��0.�e�	Z]_"���};fq������~	����Qȁ��(Z%�/��,M3R���F��'&���:i�(ۖ��bXK��Xg������e��e��<A)MQ��|V�<ӳ~	P6
�G4S����@�����Yv�y;Ȯ׬'�2Ӏ`��Uށ�o�nЄE�`mo�q��C�j9�J�5KyE�܇4>������Å���G�I	�̤����@��P!����������6yf������[����#ڀBڨE�Y��Fi/�{��ՐΠ�>�i���5��g�W��}v��f'b��9�R����P����=�RWqD�1h�T�ؑ��4گq�b�b�qp�r�������+���9y��}Qh��W�c�������#aݡ�ӗ�@�(�%<>��j�KfKn!���C?M���������8��0���Q=�1o�h���XN��[�r��z���>�&A���i�����@~��+>9\�GoQ���ܻܚv�u="f�#H�C�
�x0fk�����\�Zp&�Wm�̤��vR�?n�gӭ{��6Ԯ��nHI������D�?/�Z�I:��skG�ܹe�C�
,sz�ӹO��L33���at1A�y�e�#`����D��Ub��?z}�C��XC����tՐ�d맣���M����=I+y�b�e���l�+�>hgc��}�~��,\y�]�o�f��j<K�~�m�%h&�$�n{�g�h�0�6�>�k�������-=Xlؚ�;KL����tP����L���F�;���kj@Hjj����w�.��dZi�3������A�u����E��8o}����L��Ɉ�P��� �vreZ<}��>���*>��k�J������^b�����oc��dࢬ�p^v�L�Y}Vx��ꋸWSȃu���Å��;��0�� !�� �W#��27*|Su����bb|��A�sR�k=�ߧ*���zS��Cy>1�dd;'9%���Ui��������X4²�[&9q���⻲E�h��L,�)�P5'���=�Р.i�P�&�5�I��gQ�w��t��l<�ܩ������?����>E��C~o��]��<���3�:ҠX�?�
��tj�))G凉ݽ�9�R�c\���&8�N�6r8ɦjZd�3�MLә��]��b�랱�3�����w2����X{�+j ���D�8��������@]�VCT�-{�UP�2�4°���rgI9A�7��(l3���8@&b8�p�ze�P�7��64W"�c��_rvɸ>C](�3��9��..�����ǰ�7����	�%B�'Kv���@_�`�Nv�\�t�q��c8N%-8o�x���-�y���n�pؿ5%�6H�K��2?[>ő!`c��pz����'�xFj������<��U����e���2�ѫ,io~$-��u���l�S������t�7D�F�G��Md�`r^��&{<k�����~R�����s���>R$īǃ�x� �K?r�P�TI�U�DR�7���_�o�����j#�p��.�G��W��O���� �v�"z�͢��r�e�&�SRw���{���f*�����I�*��3~~�R��������J:�ȽU1�8�}AbԢ���溢��Q��4U0���d�\��H�)�IYo���S��{�����M̢��,�5���uf��B4�aM1�-�Q�L�ShX�JMz����r��������
�+(��=���Bo�����%���`snp�^	6��T�b'�W{,Së�ⷊ�G�[���������� �M���A�)�?'G� ����	K��B`w"��@l�� �D��Y�ml_k�<�@hP�0��ȋ+ؤ�*�	�*�3{�����U{>-?ըݧ"!������!�!7���]�/�L���i�K�j�ZUH,�{�n�S�o=p�J6�N��n ^>
I��("�.��.�a�e�����,�%$�l-$��{��� ���8Q+���2��H&Ecȏ���e���)�gwvTX�@~6���g�{�����ݤ��\���� �=%O�F!�-�X�WZ�t��r8ɨi��]�g����k�'ە�b��V�@r�g��T��!��wO1���D�G�B��nE׼`D�A����=�	w	���W&Pw�\W!@�]S���ޯ(���_*�ނR� p�=8� `�`j�w�Ce��댟�*�,��_�Q��_�VJ�y��6f-����S���ZZ��\^<�3b31�*g������A+O���mȴ4��O��vu:�ҫ����Ұ<jG�Q5mł�چ�u��m\��?!��D���Z�j���v����Nɿ�pR���Cob����$�����,z{���J�e�)�ކ��M��)h�(��Y����M�I�Y=�&�����t$�w��,�� -�g^Dݼ�GI>����f9iB���Yl�Usz�����XP_���$�W���AI��#��z�L��������Lz᳭�
��R��d`��Ǚ͋[lM�e��Ik�*�}�?r�Dۤ4��sI�(�	�o�?�>�;�����:H��TQ��.X������A�m�b$w2O�'��b��=Wz�V(+�䜦`���k������QV;���ɥ_�Z�Btۊ^�BV�JB �B��,�z�	_"��;n�¥�������d��)Pӵ�-V���-��A)ňG���~`�+Y.N���pō�m0�˛_Dfa�r=m����2Ü-;��#��t>|����xH}��E6
E�Z�:�#�u�Ɠ�̃�X%}ٵ��w��i)�ʼ�����D�v�L��	\Hy�0tݲsv�y���V��]!���sj�1<�R>���߭�j���s�$(#�����&�H�K�8F��2�����_P�L�pp��6h����.N�y)S�5�o@��;�q.M d��F{l<�,����q��ْ��g����3x�n�u�լ/n�7Ȼ�Y}�Ѥ�� 3M9�3�"��n�Amb�5���o��<t��~@��}��_�vT�{V��������?ɠ߂FƟP~�L��E����T���度�G���J�"�:c�>�N-`bW�!Ai���W
�>h}Y.?��~��X�.v��y	��w��IH�T�w�F�ѻ��ݙM�B�-�}#��J3�'e�x4���J8Uh;�~cP�w3�BjZ!
�xW�o0��n|��� � ��_Q�ŷ��
B�D��7p�cC��T��UVq��k��ź?J\C�@j�A����y�L���G^���	c��G�=(��������?��~��e��N��g{���K����v����7����C%�YAAy.�@���_tQ淸=�V���?	{7O�0/�GI׈��{���(ѳ�o��ZK���/�i���9��'W^(29 W�~�<k�8]f�G��ό��_;�P��3� �ﰛ�a��26<�7���I~�d��27���h�����XK���!��Dy�c�o��2'm�9*T%H|ɡxyå�� r`�Oi�*F1Qz!�z��'2���ͽ�r�RT�;��8y��"��g jK�}5��n<��%��<���M���Ƨ���V����%��{Z ��}c1�}��*��k�X5;���H�����=�Њ�12�	�L,/�ZF��J(�4�iV�p�:����@訑�����*Ӭn`\�c��RJ"o|dB�;6c�o"�<������Kſg������`Z�x��qb6���1%B�|�c}U*Y��D�|J�þ��9�ζ�Ȝ��7�GёF�Z�Ӽ�D��Uk;՜5*+�Ev{����1�7QZ�˲��Σ_Gj�	���0[���O�8/��9S�� ����yg��͜�乭��3�S�V���N�D������0��A�_u�
H_I��is7�d��͉G�e�5��*M&`[��6j]$Y�j;��3�z��L�r�Q��A@�Q�O{4��o�"�i��7�ـCR[�l���r�@V�ѿ�|X�1:`1�0{l�m��K�9�1pOT��WɃ1�D�0�\��ľ�8覍>��xH���5����o��>�'IO��z�"LM'�����F�%z�~���P�I������yɋ��Ʌ�3=	�laNR��3��9���/c�m��߅�,^3B�g�vp������~�1,8�N*2h�1*��(�
O��Ӟ1��n��W
�B�B^P󧎘5�<���J\f�3���G)�Hjݻ�2�	�7����tyZXY~8���o�ة�j|֙�Y<�T���x@
�'�q�
/�D����}�в���ȉoXh�U/N�wVͧ8i�C>p��{����{������ a�k�F�?Rذ-(����'���<��#�{u���{ y��V;� A*�.�]��wL��F�0�Б,d���{P��I�:Q5�}L���k�5˭����K ��"�1�9��+���%�{9�:9�(H�M$�h����#K�KI���1ג�4d?���r�1t+���T�e��夦ó�;�E�x�e�*�:����츻+�(���{���<��oO8gOdk��̠�G�1���"���]|t!��M�
�<wK����Λ�]anat�\Aw�U��!9����L��F	�/�W�_f����rwZ68b&��.���آ��T��˥��GSU���R,��ZR�q^��u�����˥3�>,>�"� f���w]�����jKb	u9����x��G�8��ϋH�`��D���:���h��C.c`���on�Yx�;���G���! -���R���|dr�O�D�y�����=3���oR-#�|T2su�|���U˽�"gF�(r��/�eѥ�x�K3��8G~#j݋g$嚱&��& ��>���Mc�L(��)�Qp��7-GZ��ezv��t8�_M�Ҵ�p�����g�"�a�a����Cq%���^���M/����e\��sp�m	�PW%}O�D���1J'�Yoiԧ�U��xB�AZ�1r��J�T�EU2�6�I?���\���Heʘ�蝼�C;�w�j,�Z���� �(\|�}K� �R+(��	��iԇ4_3���=�����Oiǳ
�O������ �O�ug���&���O�	�>�:��HE��5\�}���觰�p�t������F��u��j���*����� ����
�XD��K�m,����'##Y�f�;�u ������8�+�]}
�i�>�q���K֑�qkX,$�p���Mً��ɑD���{"n���h����{i49���5��4h�G����wqA��~��w�r�oU*|�:u*N"�c�NM�w�Q��u`����¾�M���^[Bdw�GK�������Tef�0�T��VNL�J~��1�x���SB���S�1L4�:�R����2����4<ɥŦ�[gް�2�}�Oy�<�5���ጝ�gj	��ǋ���Mhp�B���������NoJ��X�N"��9m�حg���~)���O��6_z�i"� d�\Qs��k�`���.j1&HUNL!|���=n^7�Y�Vt��A. F~u�%����r�O�D3a��V,��1r��a�XBޱ��o���u�ߚ5�B ?|�w�+ZmP���-��V�/���Oͱm-<������l\���ʞ�ЌC�����U�x-P�
/<Z�J�#������X����>�w��2�2]l�Ac
�'������?��"?��+�Y�C���^M�����t�Ǳ3+�4���
:5Sx������[�$D!?I���f�?BPF��Q'�����6�h��Vqz�,�z|����B��$��w
[����u��oC�)8���ej�x�#���8���'�����:N�)���C�Sk��k��c��`<��e�a�_�	�1	���狣0>%`�֚��A���ϧ���V�ʪ~�A,H�UI��i�h,m1���:h�����ba��HS$�[��s��Z��C��u�χ�3;>51�F�X>�>Ү�%���TX/���pΌ��R����*�3��F4������iR9��[n]`��m�E��;n�X�ݤPF�ܲaZ��9g�����]�d+}ޮַl{8ڃ�����wIH;���DVX/ӲuZnA;�m�|��`!�y�m�c~�<q����!���-�y����6
b/S9�Mr���~� =�3�-��R��a���/�����
��쵪������51������`���Ss̀x��B�V�
t����C�ou��Du�X��d�Ni�֒�huS�S�N�O�9�;�P2c�ow��I[�(D0�N�_�P�3�-���c�,���5ϵ-�6)KC�o�,���VW�>R���	^M���蟫�H5L� �CM^lg�) �A��Ɇٵ<�ؗy���z�~ۖ- _�[�lI�-.�������R�F����a;��)�ސl*yZ��pPR����yA�(�uL<��KZ�����3"C�<U���wğ�����Xɖ�-���i�Ge_�2N+!&l�v���D&�]/����<v��f��gܐ����L��aJ��z|hn4�<�c`�Z������~�ta���G��LP�L�����>l���KQ�*hܛXo������',��i�?0E/��G�����ߐ{3xm�lB)wJ6�r�O��A�[���'��l/�V�}!&��:�=�.x�E�ry�)�n��	ʍ�{7Q�9��������!�j8��Oz��8�����0�H�2�QF:��Ӻzxn���j������0��Dd��J*�>�4h��"�w/���|!�ҡ�VW��G�rq*˯���ul�V$t�wuU)�t�Z�)Adi�NeI�R�'�C|7�@�'>O�������`���{�0{k.�7����<l��}Pg��j���n6�(��E�y괺�s�/u����1�X*>ID�s�n�]�ýZ��
�
F���E�[[Ò]&�;$���Wz����&3���qʵ�|�ϪΩ��_�}���=�B�F܀؉N�����w^�'Ot7���DH�vV��\p�v����od7%�_K�
(	Y�G[�= ���~��\���Q��)�t錙fM��K
->�8M6�7����N3��uV���3�$�~6�*�1�j�����A�X#�r����@K�]]�������8p+����ǁ>#?�,�*B�$#�,�6Y8-nc�����`{WsR�����zk#�v*����.k��P�N��Y`_�<U� ����㤏�?���$�%�!�5��'�ӛs���S�'�1lG����NH�F܄%r�7N�s�~���yރ�1׹���y|/��T<|H��b=m[�W���\�'�� /S��D`sz�*
����ZF����u_gC�?�@�&)��Am^X�T_��+V$��y5]`�D���ًA�ʙS��id3��3p����op{�o�t�����.w�A��R#��[����tj#Y�h� �'=�\���$fu:[��vP�E'o��pN����U^��X�	��Ǩ����M��pݤ},>Z�*
�:6Ate�~�P��7��3V�V�)�&c1�x08v�}v�1A �A����O�	�u�d����̬ͨ��X�h� ��i[L53���X�M%�R���qj?��R��Ҁ� ��c
�J�k%K��1��k�52i����޿,;�cU�	�-�uF"l����}�h"�>��v��AO?�QPa�@�j7K����r���aa����S��lj8+9�3�Ӥ�Sm$a��<�	V��Pr��yK�5�����p�+ ���K��SLV�ȁ�r������s|dGE:$2dRm�����&	-M�B \��G7�	�d/>f��to�G�����{Q��&��xy_���u�*��l@(]-�0d��U�p�g�*� c=Ytb
PqW�����|�?���T@���w]�eD�C@ckK�-���./Ӌ���|p+�V�ۉZ��!��ɆE�nU�G��] P�����w���]yC��9��!�7��ٻ�}�����̘r$Gq���A7H0YG��0�3y�xB �%.ġO�'Db2��?_��
���f�`�t�歄5f%x�utN�i)�'̦[q�Ȓ���cd�<�b���%d~�G`җTz��?
��F��|+��q�� 1weAV�^ � U��_������	J������ض�h�K-P.��D���(�e[[�[���y�F��{�sUFιm�Vc�m$�q��쪬�b�Ǣq�ZM��v2ˡ.�'%Z�/���.��;�b�?��� ����5��`�x�O�e�Z�ׂ��� ��>){$�έ"�K�I6�xgϾ"��m�aN�Wm�D�'�q��f�":��/�&�u�*@$r�~/�ӽ$۠	�Oe����R������@�/xL�K@gܬ�ȧ
���3ŃFWu.�[,�w�(�)��b�杜����!� ��e����q���G*�B�qG0ӆ�f�|J��7�}⥐�uئ�j%<��z\�^��)j}H)����G'Xֆ����QU`ۇ��y25 ���,�z�4h<�q���w|����N�3�d�R�W�J6�X��v�ek�C�4�m�_�U��\�+��)��3����@��aCj+�vLY[�����67��w"M�ɟG!�e��Ǹ������[@&������ɍ�J����"T����د@�iӕnZ6���,8 �U�	+Ja@&���(�c���Em�De�`٩�_\�ewl�\�[y������]�$
N��������RУ��4,
Q��!b(>�'>�����¼��xGt�'�Nꈑ�9F���0q��r���z%�����8i�q>�>�Y��� �����.ƃy,aw�3���|���F�L�b���vj����eCi�T�m>��g{)����=�QKz�l+IC��͂OJ���3�^�`�G$�jGvvcxnGֲ��`�b��$�_�h�|w)�|�]tp�M�o�Y=�%�R�"��].��PɄC�DQ�4�V�/��c���ҡ��1l��@�aYo��[�:f�(,�}Eܐm\��I��h�*᪙��� 1�0�.�f�r�R����c�%̯��Rp;\��+�L���V]t�V�,���
��z��
dl�t�p.�*3����V.�`�r�v�L1b�֮Km�3�5:�ԉ�Ԝ3{?� F��b����I�K뤨i=���m�r�";ltibc)�
X\n ���/�P�8��I�Wת��}/��\��U�T�%"Y~���D���ɶ�!=����Q0��� �|�\��g�̜x5C���+^��[�;3,CB�/]I5���[F�|J� �n�����rC+�ȧ:�ԣ���.Y;��c�� ����oOXh�ɷ�l�����_r��+S�䃫a�<.���"2��Gj��b��a�"������67�ܡ�Ct��)RE�D�r��^�P�M�;� 7ZI��NeNn�Oj	���v=�,n�I����P6ڶ�Lc��#��@&3-$�1���?� �6��mڒ�>� *�.őr���2l]��
:�����T()�N%g�}�5�Kb �^�1�#�p��,4B>��I?�-x����1q=�#Ns6.g�g>����#� ��8�py3���Eh8[��Cj�<ql��OI�&ޤ�g4%{�'��Bz���x_���Ǣ�G(���@l��l�9�C��Z�������+`;Q��(V��j��Z����~��4f�:QcƧ&�����y_�%2,���O+Ϛ�w1ܖ��j��&�5W�y�]S����������RK���P�Ӡ,����	"���w���!sS�Ӷ�#�Y~&�~�9,��."�6�{�se��FS& }�J'�����(�����p����Y��6H�:.���F'%���b��"8:E��I�J�%�zz�y&L�}ς���|�	_���0a1�.̇%jS������>4 ���ʬ���ʩ��vf���U-IQF��<v]�`���)�S7��E�Ub<��-[�N�^���*���&Y�5�uhޗ�'0��{�L���������H�%�D�Z���~
Y>��D0�an���܊�\ٟ��0  �+N�� ��*qp� F����,(�v���5Jθ��o(;Z����74Q>	���D��	T��dl�<mU$�Y�����r�*{$1�J�bj�M���v.��l�����3�˧�%O���QGs3?<L��͢<��`iJ�Ob�U����U��?,0��%��	�_�Ѫ�����z�#���<�T��{�օ<>d��%�:c���Ҩ��
A��҉٘�a`���,~1K5��|��G�pڳ��ҙR��f�?��0)�̠�1STl�I�̝cD��xK�G3��������fp�	��U�/��Z�>A�Z��ƕQ��_�9(���j4֯O������c�l���T�ف���3Q}�t���o�s )����ua�(���]n7ֹ��s� ȶ�m�����;�]��"�1�qj��.-\�6���K �����?É�q�|��%���%Β},O⣟�-`���� �=9{�6�Տ���� 1
q�����1wvt����v�(�g)M���U=�^�<u�U��%�O�s�$�����n�u��	8����ZeU�Jke�ipF�,T�3�F�N��ǭw9�H!?�C����E/��u=urt큏5�x�����;R��d�`'z4}b\��C�i��F��|�*�yk<GH�(����W�o�G֕/&�+�9�<��.;�{��ӒC-�&�{+���i��R�̔�^>�a���2����g�	B�m0��BP���f]��
wt��ԈֹU�n�kEY�:�q)^���R��@�RL%�Lk������H��M�#^)�I+���<jujbr��t�1�<�"n5S�&��v�N+��"�x��pN�����0(1�t�%b�CP'�Xg���34hX*1��ĺ�(��q��/(U!����/�og�.߳;i\vX J�4�m�(X���l|��?Qk��C���9�QJ�-?ѝs��`�3]�]m!\&��S2^5�]}�n��s����,�NA�g����p�E�a����)/�q�ϑ��A_!������2`gSx}���Z�}V
�����(�t�w��@*u�yy.gW�MGMXƂRܻCB_x��fj)�47�Mwn��q�������Ť�Z�O����Ҿ� R����}�%瑏ش���E}l�6��?O޻�6�HmYB�S2q��ұ��ˠ*�<�� �i8]6�;�"���<I����5>?[���x.�}�$�3��  �y�G��\4ҁ$�f�A):�կuz�����,`�5����B�&�|'{^�zr��*`n��5C��F �P�Ɵ��<0���`�iɸ����d.�yߊ]ϱ&HZ=Yw������h�������3��M8(������G�\OxUR����$Z����>�pK`p�;�WÆb8��n��8j	����	���Q+ˌV�9��B��gi�"o��`���_��=�Ј��|�=�w0�#0��TM�|�Iz���o�xi�ž@�呂��#d~Ig�q���ĥYH�v�������nU�E� ��
�p�
�6��%�����ǐN��n�M������u8�_���vy��a`����e��D~�O�����,�}��Nw��N䰂�E���3�څ��z٭��/9�����q��p��IV&��F�z��>��w���S�3�L�)x١o;�N��e`%*����=�l�>p�S1.��;՝�|��G%�o��k6�����hr}�L��@��Ը�ja��,��S&�`���b._���D4�������\x��H��Z���p��ET��� ����c�j*�qq�:z���Ҧ6t��d3�(��X2��\d "�kѭ��l��՚�N2Lb���7'+�á��a�Xs�K�˾U�AGl��$[a��~��f��癚�c?�?b��������qv�7�RwZ3�7��T]�ׇM�t��ͨ�E��Y�`}��{DK�eB���fF�۬��y��2l�mKJ;tK��"��,�r��y#z�k9�ȃk/H�o�����k���x[�����|��Ȩ7�]�nQ��OY��蚶=�}�3�?0RS�xo��ϲO?"3K�|�+��[Ӫ�%L�h�7@i%fʰ՞��s�qR�,��y���>�k�V�µb�i��B�jv��@��<Ǉ;��r��ڵeQ�W1�p2�1%���V�1�=���K���xVY�XУ������8Ժ�	��!&�c��qc��-�Co��ë{։��%�K|�K:cB5g��>+�<Y߉�
o
��f��P2W��䨿��4-��z^�s(��F3�N��e�0��3�UC�"�EHy,�O$6���;M{�k��g�D�Ӝ�ﮁ,����诵u^�.K���G���W�=a�W��Rb��&��B}t;ؑSF}qW�P;y��F׎��ó�쏓1�� �Ȋ%�z��#�8K|�*I@� ��݆��&�s�'���~T�#�ؤR?�'�z�~&SB�#�w�n�������!�Ȱ��	)̽��56BB��W��H|g9�ll�P=��jzm�xb��bd$��6:#��s�A_�:Ps�����j�WH�A�Ȅ4ݲ'��&"g�m�K�,b&&�ゎں���P�:��|�W!��`���JqIaB>�����~
}#ȶ��25&���C
2͟��>\L/u����Wv򖡅Ŝ�{5:�P��wkW�=�H@���|��q���h�#bB�-����_��,����oβ�wz��v�8e7Xd�����o����D�9=GNQc	�x uc�#��3���_�z���;̹��Ynug�q�W*Ny�՞g��'���P�$M*���RO'�B4㊴ְ`�j2���������-���ﲤoK�t������Wa��W���
��C9�ڵ���k.��P@ =SLv�d/G�M*߬3�Ë|�\N�E&O����`�ae�=���}�{��a�r6���L͈�5>Q��=#�E�X�\*����X�|�,�$�|���{6���z�J>h�;</��y��h�yT�;{_��Z'ֳU���{�#����j(�`��P���fd�:�����F��
��t7�A��y>�~���b�A�ʤf��VVܦ=H��� �,:+���K�=�[�i�O�����]-zMLL!��ܩ�N��R=�8��TН�K���`��z�V�@��C��'�xw`��Id�����:g�
Z��ƘG�Sc�Ќ�s�S����Wס�&FKe�%а�u�> P�ǻ=숚��p�R���������+/m�C���t�?�wK���t��/HQ>H93P睙�=��f@�����DŴ�鉵>鿙�:2�;���zh�A0�LJ�7�[�뮒m��4���7��Z��2�� Χ�+�D�Z��Nj�H$)}���X��j��k���Ƨ�-���Y����Э���1'�ܛ�%	�<�U�H�亨����w*��Y֭� �U�%m^�4%Gr��v����FU��Lnv���/S����x�Uј�n�B���˷p	��4<b��c-�a[>���c6[��0��xČl	��H�-"B�7,+`}]=	�#������?���J�@��؅y8QٽJ���z��9�50;T�-ɫ6\ٛ4��롔�j�
{���n��Lۜ��{�~����<�UI����.\¹3վ��#U|���Ytڍ,)$�C�0�^�o��vڑ�8�X;3!�H��l���(��2w'5aF� ����Ј���U!�V��y����gs��,˻"ܲ�0~�2�T��ޑ6�� 0S�����χ��!��#p�o\�w��z��^4(��#Ա��?l���<לegȻ�I`��X��_<\�?4��ÿr�ɛC��32r&`5w����	�J���^c�1�A>g�KX�!� �JU��o5
���{J$a̿~�|X����ʰ�.�9�"�ۏ��?ƚr��JAf���^�����_�l��&a�?�A����[�v-y�d=�>���4���vh���N�h��A��h!��<���3F'������k���/�5B-%vQIa��!�oJ��S�t߲7)p󾫝R	�x�9ؔEG��r��ԩ�2�:��jT(���O����](4P8̅Q�=������^t`�ʍ"bY�ffdͤ������~-��զ8��=�:�N�9$�B߱���l��j�0�9���C���pu����	��U.�V#++�!��=s��ȜRe���iV���Ei�v�a�!��\JOb̺�m�/zVU��<՞!m>���c��ƺ��u5N��5�����6̷��+���sdH�)�?�4�"�=Ҕ�P�}u��� J��ϻL�f��V���9���HWpvJS��M�)kR,7���h��*��$�M�@�Z~;Һ2��v�%���� ���`hq`ǩl~��W�_�a�o���Ws�*Й��;W�M�TD��8�e��Z.~Fڹ#'�UE�ͫ��,��\��H�zd��/ub(��
��Z�DtA�w���Ҍ~\Þ�2=T��-�,ܒ�EP2}�:�vMrOS�����
:lMަmP9��(�ٸ"T�t��r�Ҍ{�ִ�u �����ب�?��M���ǁ���䗩�@�p��m����l8{�]�9+��vd�Kt�y�����DL���ƥ��T�"�{�]�C�xà˥�����v)�s�4�ň�8ϔ��++���h$1W<CK�1%�C���D8�?sT��g.]8 ���P��������>
 �#� %2՞�����8o;�b�.\������b�����t�}�Yw�Xs6�H�� |��G��Y6Z���I�D��ݩ>�Jd����͓e}c��0_;�+�o%5�.������'j��! �s��J�>�7Y�0�
ֵ��F���'i�ɵ|/xO����o�O��#���|E/���7H�p⾱�w3�=xt��j
,��>,/� �w�Z���(P��@�th���~�%��ץ��^�hU��7U�6��{�������6F��H�u�x�=cM���d�����g�U�m{���6@��L�<t��}µ^ɕ��nW��&��j-�	�	�GG#�!ȑ�N��(�K��p]��u1h��!<��z`3�P�׶�b,�f����ʦU	ˎ�l�2	�*ɗ�����&�QL��m���n&���+L�+�cK�$c�Z�&��v`�8yLu�iC%�h��M�ӕ���Ǵ��RC�Z ��Y#�Vi�}�`�U ��O�i�{FE���Tu&c�\�4Zǚ~����O3e�%�D�ç�N�� ��.�IH:+pG������W!�*	Лf�=H����兛«��"�*�ݔ��*P~�;̸%;�y��R�S�Ί�G���7R��|�&��S�ϳ&���[V�ޞ�߉�X}d&�NT�	e9�իhdsDt
�062�@�qU��� 3��S�+-�`7�<�9f�pj!;��v{��#ohJ��d��5�F!���-��B�̳����|,2��7�C��0����mR�BQ�3�]]g?R-|��`�	��,�x5�LY��|B�	Ec�e$�������t�C��	v�ܱ(i@:\���Tc:/�|���d�LW� ���2ǂS�|c�=�����t�و�g"캽gv��$��/LHm�S����Ft� �~�O{-����/��{Î��F4�y�b��|ETF��S�Q�,䠉l���Ȑ@M��R~��	��Aqx�J�o]�Ir;��(���C=��x��[	{��+�:�b�6�S��� �����˃��i���ݽy5������5�_��5u��R�n�Ϝ��c�U�B��]+{,��!EhF�����Q^���Z��6m6ʡ�I�����Co ����z�����-y+��G�2��q�5�#�D�=�_�}�_�{?�l�(L9��1���_��e7��l���;Ä��F7�=�[�� ���GW�7���������qO��d ����e���!;0�.�5C����Y`�J~ԩo�:������3�&�(i�5�^Ƕ�.d�G��g���@�p�2���~�UQ&`�@��q6�׀�`���(���fT�p-]�$��TF;?;�|·gMjq*�Rl,k���uI��B\/g��¿�؈�A������3vE��e�e��L�tF�Ѣ��ud���R��h��HZ@��w�;8Z^`��b�b�ŝR��A�I��I	&=��X�F������p��殦)�0O:0��˝N�No�1����89i����,�^x5������l�S�U�V�B�y�O`7�h�I�y�E�����x
Ag<!�Y/0�6��-�����ݝ$�"��K�3�:���/s؜�>�+���j^�6�2��$��{� m�Z���3rY��9o����k6��ȔLN&~u���R����?��tv�/�:����|�r�X���~\`�0�a����|ٯB�`�~,a�1��Ĉk��u9B ��u"��y�"}?�|��%�s���3��j0K���*�<����0oN�>�_�����]9��!����*�͈�{aDbR��a(�!p&�p��p�5�: D��9{N�o���"��]m9<+k�����k�C�|vr<?�?)=�=I�Z�5!�A%KAvOv��Z$^^�{j��8"�Ld��ܭ5\`Ti1׾6M� �8����0�v���9�4�����t�	=:�40��ˣ����=o��a���UL� ��W��s}���^83`�ok�7c�o��m�bn��� rY��ON�0PlL�t�p��V�dn�D�߈ÿ�GPsѻ�c�=� �m��h�怋/����Cj���;��Vӈ{	�2��JQ�]q�Q���@��jf���'�U�te�8�1�|��<j����L�H��R�T�dM�f6+��n�D���y�<��Z����3M�z)�Q�αxwख���KA�m��C�����q��Y1����z�v|�0���;��_Ws��RKr���i�����1��ݪ%���Q:�%{m�
���j�Ee�P�+�\��q�8�T1`~�M�L�@�Ҁ@�6f2X_�VRXՇ#F���V!�K����3:G��O�2�BS��Ӟ��O����Y�i����~y1��*����bJ�%����_��������Ì�>-�Q[�T��~�P� ּ�f�ԣS�"�gAڂ����yU6p�v���|:\��z3tȶPF;��PP'���K��o�6���P��~�'wrcE��z�Ho�����+�u�*~�:�jW�,0}j�B���k�dAAC�͜�p=u����_E��׮ͼZ������g+��1�b�&Wlv���K8ԡM\-��&�1���rרs�=�ɍ��`�A��f)�����V��#ڄ����A[�!(�kC+�;-����U8�O�T�v=��k¯�:G���kc�KbA �fZ��&��;(VK���&�%ӂ�[t����'�I�1�i�Z��bA~�~I�'V��'���� h�QG���]�j�L|�����m;?��ϡψ�(��],+�������']T5UyK�ܼ��G��]��rC�Ks�C����U��4�:�-;��N��+��1`��z����� ��hP���5����j���{B���qI��Xy�I�K�$�Bl�d>��!�Z���`�3{���q��/���p;LP�zG�i�p�R�K�z����"&�/-S�bt\K|������p���T���O�W�Oc'j_&��0�?��- ��:�)�dA4s���e%�hc[�T��\VƦP�=���tN�������XL?«*�1&�=�
9HkO��q�c�}���J�#���	�������<C]����vv�^���w�Cy|wb�sk�Foй��x����F�K�A\W���n�� ���`�� ��8�������eĄ�fa��>
I��4Z*�VM�	�غ���Q1aY�t�]{��+��㛭l�`ck%^���[�e����i��w��uT�Ͱ�����]2��tL
f����	0}��t/�2;��y8i"o��9&G�y�-$��t�q�vjXdר�{��Bє�� ���0�g#~��-E�q��1�� ����C~��[�����h�r$?��m����N����z�8xv�y��T%u�'�\)Y\�������`�	�<jɈn���og\�=?ujmϥ��Zc]���v��pѴ��<u�z}7.M,V���݆��=���;�^�r������".���%�u]���3�dx� �6�]�P�5�*�����Adt�#��<zfbR׋48tHC�s�S�T��)z�l��.��!d���d�<��{~��
�QF�V�|1���^+664A���6+�%� �#|ݩGݢ�,ٮ����3��2�|���[~�5���ŭ�}�C�إUѮA��F���-�y��˨�(�B�]p�������Uwę؎u ��ۍŭ�LC�\�M����e�e���]_
����/���z;������3l��HX����c�wݰq_>�����ٕ�a���`Ά;o?_�3,�N�a�~"~-["�g����-X���2�R=Ny��5�݅������m>({�����bɁ���y�nR��doKM���?n�:UV��h�N#:T���M�e���nB�8:���`Τ�k|L|R②��~p�`c�ʦs�wj.uX.��9���)�C|\S��27�"`���v��[�R���p!��ҬM��Si�V�'0��T~�C�۩��â\(�W%��io��
��a�{.�{mS1�r�ɰ���� �QD�Z���#-`�SL�.:u?͓O�k�4Y�o�_��筶Ó�x��$��!�x�%�%k+@H�l05{�B1����d��y�5�8�,��03�^���3�oL�����C	��8g�W�f���C��_���z	�-�I)K*m�E�4�rŲ�5�] BEU�I��[�kh���kL�~T��ׇ�A���A_�^=��ߕ"+>�M�� [������Ă�ng�ay��VX�iLC���8ۻ��wd�n� �յ�A_�6�;8�f���������2W'�?Ph0�1���t���Č�1�`]�|�z�X���A���ŚOo��p-n���L�uf�o�Q�^l ����_#p�w"ӛS�2L	|�)���n�9<g�X���0�������$8Z/�x�,�����~ Ձa�	��0A'�M$I�FB�7=ݓ��>\t�6����E��V�O�Q��z���7<J��U�}m2W!�Z��b_?�O�^V$�9;)����X�E�nP��ӣ�ϖ(�E��K�AV'���h�g�MB��ps(Թ��������
��bO�ӼԼl��7���)E]�!���
�Wx��k�?U� D�m�i�ibآ�b��$=��U���Oh]��37��>�EC���|�U�U��A�Lt�[o�QAJ�o�:3�Q��s-�\Xag�e�vV�Ћ�t����=F��J�/��ŕl ����͒5��ib�Ǩ�J_���t��]-�v�I�h�2����1�J$�\!�ڬ>����?�N\��q�)��ڙ��"�xw��}�Iv�*J���k{�`jb�4�|-��0�_5P�b�aA�]3<#E���uz~$Tf
)�9�U�s�uλp�i��=�[^l&���y6qp=֣:r��
�R�x�0��-�e#����*ͨT�k7/W��)�gh?c�)f2�8:��K)ڝ�>��(����r����8�آ���dxH瑩�4��k�e�\��W0v`��i,�*-�e��5�e���F�[�@����3X1��h*F�I�����mXڽM��d��O��U`��������F���UU��v4�Q��ZX��1񘮧�"F�����Uk�3 W˸�i�I��z4H^�C�c4'z�sXB����d���W x\�yj"���=P|��d���:@��U���%z����EC `�f�pFG�ь����A]?xn~��k��O	�h���~lh`��{8'���O!���Ĉ�sv�V� 7yD�[��\��1�1��t�w���������=����D\乑���f�S~$���ȶq��~G�3f%}Boq�*7�`�>�ņ��'��1��PD]>tʯd�Q��J�[J\�n:�ڴ���cY����a�H_���lQ��J�.�3����G�T���`ը�������%J?P{q����Q'���z�d =�^���,��A�{�Ef��u��y&&W��	�%�J��A�d�yO��>G�(Fj���8w}(w���[{d 8B&"<�^���U���f�uqh(0z�ǟ�4��#��G�kF5'�#q|va
T�0��Dct)x�8�pG�htI�4W����-,�2p�9+�Pk�b�����,�PÅ�d����$��$�?���N��^�	k=�\�;g��49ޫj�❍$+��b`K9JY��d�k����<F:bKqK�ǡ�>�/Қ��m\M����R�����M5��p�����^ɘ�9�P�����f#'��0���;��Ԗ�E�I�	m��x�r�_u��>��}y�dA�=+*^S���B���K1b"�����Ln�x|O\�^����S��m���ZХky�t	 �#b>?!�ju��xz@z�B��]��l������)��*��V�0׬ֻ��/>���#F��Ū�\'��rѰ�T�<V�P�:>M�ޘs�U�W� �"�^�4�f���2B�K� ��hV�}W�4�Y �S~���Gˡew������A@��1��ҟ�Z�#�BM���g��?���<��9��N ߬7�Б���XR�k&��;S�)��p,�F฻��n���Y�L�ȓ�	�+b�Q���r:{Ǧ!�±��,9y&s�?ܕ�tW�HL,�;W�qZ�j�D��	��	�C�4�h�J�0��c�c�7��HSӫ�y���<�õ�DA�±�=�@�D�(��
���m`�n�0�n�F;�j�+�z�ٻX�W�q[�9��z����a�^���pT2z���$[
f��A2W�VP(Q�z�N�����e�0�DUb���1�w��|;���3�k(�X��$�<���ڽ+�mU#M���An(�e���o.Sj��>i���V㫕��㪨\��=Q�}8h2{��[����Q�@Sq�@"�N�Q�aPt��:]��~zD=�9�, C��\��SU��5öy�*���y
������ΧSL�ʸ��#�5#�>�R0k��������jt,}�`^����Uk���\�tI�����.G�($��`9�^HI�%��H�Z��z��{��pk��4��iu�����j��	�0�Jm�]>�i��G���1�����D�xeMkIS�n��Q��� {>H�����錿�70y��:�d{g�9����t˺qi��tN�&�i������؉�J���	��ȋ�UV�'j�Ǭ�+F�>4���J�t!n;nR.8�9(I%�h�LeT�!�F1����E���Ǆ�G��t�Б�X��E��rl.��:�T����h������+V+���`�k�p��h� ����"?���眬�)���e;|��h � ӹ�_��]��S�(_%ݚ	0�G��N��m�L״���oc�$SU_�� l9�TPЎ��� ,��N�2�ad~Q��;�� ���v˾�`�{df����"L[j�f~��������1����MM�=Q�b0�������`��|I����x[����&��S��u�q8i����z+��)%�i
�1����C�3���^���I�t���X�5eWN	+0;�@�}'��$��Jeyr���C���P�Ī�i�1��jI	;���$�T<�r�M7��#�
,1�!d�j�~�`���B��VZ��P��#��v|����4�Q��.�҂ժW��M�X1�2r�[öp��%*�J����{1F���努����/��S?����B	* C���ùH��-����o\���Ӄ�#��ʡ]U�1�#�~Jp9~�C�$p.f�̸�_�^3E2=��,��)��,���۬H������fN�=�S
��i���G-�;�)�w���@f-�dKI�=5�u��_�測�
���BcQ]�a40�QT�"��g{��#P�4z��bݑ
@�T�s"?D��lP&nEue,`ѹF֗����%�؆p�q��߾<B!"U{��&�S�Q�G�(�͟zO�kFY��Zd�ZP�ē�t^�R>��ݟ�<�B�8E�'��Ł [�/�g���R/����f����#�4�B�������ɥ��
UI2깰*�m��;�&+V�$�V7oQ��m���>t?5<yn*Hqr����f�]�e�N۾��m���n��#x;����$U����k��͏@<�یeV#�Z1��cpZ��W<�P�ϕ�M8���G�7����Ke"[��h���*���@	t+�S�4�7xcҌ[Zp�/�1˸/��ұI�"��4�U���1>:5,�Lz��H]ؔ��{xj',|�6/�K�p|��aIQ�]��g2�]�g6��wH��x���>Iթ�v��_6�!�1@;�9� ��h(K�(�Ӕ�/>`���m�'GG��-l��xGc��(׋�o�����;O��s8dk���xX׸;/�| ��k��Ћ����H5m�p���O�v�yҫM굄3,�,�a6_ůG�������<;Y�tNNT���O�����!R����t}z��������I�����썣�lϝ�	�B�os�vV�f͠���A��J��WX��W(K7+���L{�|(p��d�9W?ͫ&j���q�p0RM� �f�b=�/�dw�s�8���o���X�S�9�Tn;*��J�p�I��#c���N�����{�����(:[!H�2���/�n��Q������{�53Ax�>!�E����A
|�LT\wlܘô�����9�!�x��o�D�w��\{�9��$Z2@��2rB։;(T��M7���D,1�A+�Ϻ�Qs��g<��Y%�`��uG�s�=��e��!J{���i�|�VR�Zu32�"��c���MNJ�����P�7F:Fؚ
��|2���Y�Mך֩���,xU��uw�{�c(7N�J
t@�	'q�\��!(>Md���<�'��<�^�4k��k��L��Y	�'^��K3���6j�F� ���.b��\�nP�'p�R�9���~S�`��t ���EOw�dX�4L��Fz🍊}��DɀL%�H��т	&��F�jR��i���,��յ��c�c\>�g��"_#$l�k��
�s�Ia��Ⴕæ�����}��^�>{Z}웝%ͣͯ��_�76J3���|��m�c�c'�ue����p< ��7I�����:&v�S3�@v�����L�]I�XhozD
��f�7D����"+$��;�3�?����-)O�����IF蹐^(+=	����/��Wg�!��G+����Z���b�D�f��o{'ӵ)��<2̀C���0��勤�d�ύ��jek���3$ ��[2`�MB�9��.~V�4�,�'*����
�Dj5�����f���ly;M��֧RRw'm�:Εy�1n5k.�y�ɜ��\q����h�����ÇZp��E��ǆ�;D2���q9�FS�e;��'�X��g�YÛ,R�c֯q�kv���҉����=1ƪ�5���8�3U��@�p@i1���J�	hV~b��zA�h4���]`nP� `���/
��"��ɪ��O�lU�(7攘�wоV5A�_9��^�L�����Z:�fF2�Dʮ-�����я�-E:�����D��u�U5i1z�RUB�]�������6�ѣ�ҳ�*`k7���7?��d�kռ��L9�R+�ٙn�ev�f���|�/RIO��ԙ&ջi���}�xC*�����f������3�s5�X�(��O�P�F�v�.==�\6a��)P>��L�.�8�YҡNם��D����d3n���'