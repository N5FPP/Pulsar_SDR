��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@���$U[H_#�/8�y��,��F��`G�m6f�f�aiI`������tC����dl���=eZ��^�٭����B�FYĸX�G�����݁�]}~�s�cC�_ �c��2)�}ma�dظ��v}�b"@@�c�
l�bx���,���M�4A<�r���w�$�S߇��`w���~p�lV8���
��%�4�0Q�Hj������8�Wnwx�5|%�B4|y��<���C�bA��T�N���Ζ�:U���J�::��;��B��O����k�q��Q'�O"�h$ZrgtI���IB�Q��s��P=�=�F��Q�4d�mM���v�#��D����)0 G<��^� �_�\�y(����¬.��	�y�* ���Ob$�}h��@y��y���ѫ��A�".R�]�hڳ��2��}Έ:�g�wQ� ��)��E�w��V9w{cJ�d��(�	0b�9k�X�� mKٺf�רZ�[4D��<0p?���T�4)G��L[7[�4�l+-
X�tv{Z����N�8O��B�埑{�	"�=%����Q�FF��bi@7��J�5V��n��fo��; ���Cn��m�s`%s�*�+u+��p�m�|:��d�%Oʴg�6�A� i��8��tK�K@k�W��'��X�@�0���K?n{ץ4Ej����=��l�=
q̤��+'<�-AOU^uO�����h��E�!A�M�]������w�l��C�h�a+�����?���{��}e��_����9�O�н1���8����J����j�H�R��T��f��ڛ�.}��դe��;rJz~ل!���̽v�Q(����O�i:
I>{��d��Q��r�D~;�������wB� �����AP��rB`�\$�Bg�E��Xzy#0-IA~2���A�K6Q,��z������JX��	�����%ӟ�ݙL�?��f"S���s��w0���i��@�j X��P{q�$,�q�Qi�l{�̝V{�-&,�'g��V�jht`���XoN���~Z��=+z�F�	"��M��LՁ<@jN���t��s��o��,�w3!5�>�:+���y�F�"�+����}����7Sd�� ������h��U��UIf�Y���x��6�h8Af.���� ��Y�}9��!1gCZD��1�P�u��S5�Y�mN����)_�n8�n��S< 5��Ś��o;�k�f�<^N�
�'����U���m���hI؅]9h8�B[�T��3ǂ�"e_��dj(l<�N�t� NL����'U���o0�%ga>��0�nG�O
67y����ГI<����я5����_ݤ�=liJ��R:�a�/����E�]l��|דю��ܷzH�*0��q�m�+�N6j��bx}a� d�1(�l���	��+6+E��ֽ~�G�K7j�cͰ���Molr/3ZQT��,���t���Ǳe{d'�x�t���=�-�c�H��L�L������~��@A�oYf�*|4u�-�]u��/�2a��S��m�q�M��X��3�2}��$d�m�`�{`�6Cx�N����T�;yx��X�+4�4���;�����HK~�YM��M���@��d}�=B���?H�O�y�T����4������Xs�4I9y�9�f�y1�XR燎}�W%p�U�=j�.�$��W�K�5~�AW+NHhK��~�t����t���'p����>LXv����\}+��3�ޮ��5EU«'z=�Ҟ��#��>H�.!@Q?����FK»h�D�ǐu�5 ��w���C#�+�hB�Wb�j�>�DQj��PF#�5�K�@��n��͏�Θ��m2�tg9�)z^�c�N����s'�Md�e��y�hj=���z���c�T����C���'�j��#3*=⒄��CG:l��z纬�9f�zym��}#�d,'�V�9��G_ �8Z"J�lŔl���TU|k@P����:>i�m�8��&�cG�t.-8�9 j)[��[�|��r>&{Q״�HH�ߘdp��M��߸�M�_��%TL�/�Ƃ�\�M�nK��e´����+��d�gt���H�#���E24E#�!
)�Ҩ�YMi �;�,؇�̻I�9�V��?K(�t����9�tN��"<N����1���~�8 N�E=�������7��
��"/����U "4v��+!��_\��F�2�0����wIL@�(� ��t,�G�����d�Ѹ;UBqV0��#�HD}�o��"��G՗��j�ixd�z,�F-Q׷���I�,��wY�p���Zc�9��E�	Ml�uʙ%]��1g��������Z���>��?7G�W\To��������<����|���r�c���$~)Bh��S�y��X��O�������&���N�0�r����*ys��~�)�I��gZ2v���b-�d�-4o�b�(#l6h��p��\:�B"7��]�]�b�X�xX�������#B�g��/�?��Q�ݞC_�!p���r�r1�8�����ϓT���'v��v�KL�m�b��	��v� B��@�".S2�VB|5�VW���ܗ%�����r�A*8v���O��pk�/�f&G��2�Tk�鉴�?�~`�PHm�1EA����ǎ�=��Θ�O����$�B���
2�Gj0J!*ʧ	�L�� �[�3����a���s�w��Eέʼ�n.��y��j	lr䕫QߌI�l������e�5��.n<h�뫈n���=�khX����˂�P���ߎg�|�Q�ò֭ ��R��)ʕa�GRY�a�o��O6a8}} ��ok�D���( %���M9h���"u�u��A��_�=�ɢK~��b��t��J.;�C�XI��B��˳���Z|�+&�~�Wo@~���32�#N����x4�G!qV�����Q+�R�э:P���G6d�Gˍ{(bL\�r�Ooow<���S`*����ē�W���r��Cy��ԏ8Uޑ�u&�)D��;)�~�cz����r
>�^�v�G�n�ɺDU82��x{���A��k�Ѯ�
��`�Y��L�^��o�(I�2��6���X��n�6����}�y�7Hb�̡:��Ғ���3q:'}�\���hN��)݄��Y���R�Ӝ�*H�!(���Ig�
�'�H��z�Mo�!n��MUM�n��1��t�a�^�#Hn��A��"�d�t��t�$�|�f�[�u�E/^qZ��מ��p����q�8�^`��b�NWc�Cu���⼝�����Y:�S;�5�T?�����%?�����#�]w��pa�����4��L-��B��c��%��!�h�W���GbG&���0���/�s�z쟀��[tt6v-G[;}�{�LA�~k��
�_M�Z�z�w�Ih-c_���֥$��d�
��$0��uU�$���jf��儡m��Ra���
�g|��o��4���@��g���`p�3B]�r���/Z}�9&�ݘ-G�ݠE;���;ͮ�-���&�x�zN��*�sBJ1��&p|z.9�}�T���<%l6�Tg"<��U�� ˳�D<�=��g�.\g��]`�B"D��/�<�p5;|(|8�n��գz��~���bܨk���uD��udy�zԒ��	H�Qk(�NaE1��*L¦��f�.B�yg�!���b662p
�;���Imbz:cK>up/-�����{ ͇����I^_�C�	�Kz
���z����z5���c��q��GE��]�*�8I���"�x��u�^�&�|�Rs�+��l��g���ql����EC�-��?h��t˄CL�[�=Uw~����MTe���6z���,��A��)�ਖ਼vBB�m&�k ��L����3bi(K�$9�S��"�����CȮ0d^���ޒ��|����8�b�>d�3�b�ֲa�o��?@0����;�~A��ͪ��#��k8�2��WKr1�h������F����E����4].��h�b�:� �.#�J5){
�������$��C"F���JC~�]��?A0Ν|��T��25��̝�^�te���0#�U{V� ���r;%D����%��w�����ѹW�u��`-�u���L�Zb�