��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��)sZtYzѦ�#����������^{���f����@,�B���ul@k�"T�z-��0��{�oQU�<cM i��CV��Ǣ���j*��>3���B��1����ݿGi�b�2g��8��H�2m��@�}
�G%�p���.�x�T$X�v
��;�b$C����f$����D�j����+���DM�#��k/��|�S��p�k�ҘMw�����t���3��	�ΆLww���LG�\��*B/qR�n�d�"O��
���<�[�ٮ<��?^�+�#�����\`2Y�Ϗ�cR�W�G���	@oU�z%�� �˗�#�fŪx��>��1=��&��mErc��ϿY>g#d����WQ��Q��h�.�8� {J��=}�17=E-�挴ە&0�3HFq���F�W]E:ń�{�B:�(��=Y��َ�o5qxE�~�4 %te���s�6cܮu_�b+�K�s�_H��м����-�]�Ô9s���f�Y�5@�(�:Fl���t�����"���s,*�D|�ޝ�'/J���v5�������n���4��>� W����� ��驣�֢�7]�DÚ�\�y-DӢr�X��5����}'�E3c�j��6�۫�����0D>��Tf�G3�>�~�0e� ��d'ɔl�GP�j0d�S�T@|�;�'���t�C����K�j������E��n1�$b9��z��!��o��1V��%��xh�Xy�����B"�u����hk-)���7�b�ψ�V�*�㿓M�}0K���.��"����6�4�yjᔌ �a�o��������6�1s���S��.��j9��;�;��|K��Z�n�>D���z,��N�y\ko�h�a%lc��ᚣ�a�rN"�wH<w�ś��ŋ����S�E��!<�v�#�>՞J�r��)�UJ8�������I��s���H~d	$�<�u����y�v�|K��x74cjE���w����v�[��P���i�@H�����{%��l��~_�T~���UL�*vv�Eg�H<�*�X�o[T��[2�ٍnX�D2C��驜b�&�R� �S=�΅ƙp��`��F�Y��j2L���1D_�t!-��lMfl#eO�r��$��t� hK��-+p7�Lj�6�d��I^kJx�m�>�c���r��D
����*���h�R�Ű8��R/�F8t�9}F��:��|I����l� 
H	ƕW�T�_o~F��^�f�3t�_py8���P����T���F���F{�xK
�fb� �T�sy;��9� �C�>ŀp�yw�|�� �q�+Ѻ�Rh�«E��0Ȳ���� �A����܅id���΀k��Qn �}�4�\m��Y���>D�H7R�N�9�=�4D���K��}�4^u��V�s�X�(���$ m.�(�+�4�Wl�χ�:���T�n48� �|̞���m#	s�Ia���#�J��8۔�sf�ݪJ��{s�X�b��R"T޻��91Qp��p˯s�.eR�eT�ףN�h�r��є}����k*;i)2�!�YI���qn21��� ��&�[*)�����F�
p�����K̍�i*<���q�9���=��3�J�����`4~��)�<Wm�����Lj�$O��p	?#UyEN�>݁t󵜜F�_�[D���f��a)��d�VK���(�$�αtn�x����OP"���������<����,�P��!U�nT�Z��2
:N���O�&���P���/��iWbv��+T��B�Vюm�&���g��8x,�T� ɩ�)n�h�Z���K�ŃsEa�q5D�\�+p�m�i����ʖ;R����~u��ӡY�0ۢ��zY����i��)飔��[��g�c�����q���rE�'เ1�W����V�o.8ʮ_�u� �]���!�`H"G�����чq��1���'6��l|t纍��<�
M�[�v�,}�H���1n��U��q���ws캏q��䥢B@X����{ �4ۯ%���H sޘFW'ߎ>z���ͭ�)�������`H�3�Sqx�j�Ќ\p�����0ݪ�EM��e��`�D������Gn��'�f-۷��J�`���$��F��4�bi����]��ўk+7��0����ǡ�L��߱t6�,�90a��0�iw[9�o�B�5��⬲�L�%��c��1M����<��Y/S-��G8�M�ӆ�������i�QX���V�eI��r_��	6b�Ue3�7��:�z�~(�X�x&tN�nK%�FQ�x	ʙI2w& L�֐�޾�+��-��J��E|,\*:����u�����34P�M9�2� ��q;u-!4�M�ʫ��z���Dt��X8�Wa�S���=���(��8�D�d{E°>�7�f������K�(@1����l�{R�כ���rUk紋�=������r��Rf�v1KF$O�=�0]���g�{ղ"�H���"t��Z	���06 ��F�v�G���7w�7���L+�u8	ܤ�|��K�D)i�
�ŋ¸G��� SX�prD�!���r<�y�M섊�(xV�2�l���.?��Ǉ��v�����&�#�6���+w��n���|=/قܾ!���#_kqowƭ5�M���|�k�z��åM����TJb|��=ϭ�/��zW݄|��^Ӻ��ٶf.g����V�X
���SDٔCjE��_�P�m$�5��$�n��C�0V:����wd&s����k�����G&��\�2aMv��������m��6<������kG���m�%�l�`ua�F���*�H����&.��:��üK��B4��.�����z���1s��x�~�/�O��-����q�l����`�*�3��y�с��[�@�_��g�w��ф�e3��Ȑ:T8��q{Kzqu`��.�h�#�m�1�k»�R��� ��>T�+]�=���TI�������i^�O������[K�m����c�Ѯv%��1���8��*W��pᷗ�L򫌑)<6��?mB�ܷ�8VH�� �Q�S�"r*�o=A� c3R,��+�$� ����"^���D���T�-��ɸ���RI�^�!�����p袴����S�s?��Z��f�'[-,�;�o��>�&�%��0j3�3�t��!^A�E��?6=X9�D %q��$�3�P� �hO�V4B�{�Ɠ58���H��V�����f���z���J�A�լ|���kR7ak=2�6jv� ֽ�vQ��ش�|I��w]Dfw7�+��zŇx�Rq���sKSρN���"ʔ��V�p�^$�FJ.0ߧ������|�%B��<�˙l ��-M�cO�s�f�ֿ�7���e�h@�:��8�\4�'{' q�M�9
���+iQ�m�A�^�ky�$�U�8֒�o�3E��0�r����E*{��K��"�s�.��ұbP�
+��K �6�J��u/b�IX.n.(@��O��)�{8�|(�$<XH�S�b��vf7��*�"6՚�c�h>�� �i���su�_�vS�0��k�vu��j(����@"�����v�k�Qn6
���U�����O	nQ�Z�cJ]���b��H��$� ESST���﷖Zpߝ���w��)�