��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VYkM�#j>c߈Nw�&&�x��/�i~z���&�M*�l����e�Z/r��hrh�}��F��\_�BU0KY�:��j��K.�Fgt?�[�N-�a`�U���p.�߿B��!AB�پ&6��9}K0�(��˰��Ѝ�Ԗ-*��|�ߊ�Wf���Б������0(��(��>�M�-0@�|o����;\p��q)�cry�4���tP�*�'���%>�ϸM��ж��}�-Oc�/*�K�N����h��+��<t�Ϧc�
�K�������h����V� ��|�ƣi:�[�U6�kX�x��ֳ��p�p�v��W'G�F8Nk��P,�Y�p�p�S��A�7��D �<�֧`B��=Q�P��9$s�ye���2?���\H����C$#7,��-�
��g�G��.����'>�eVYy��μ�P3�"���97����D������-���/�Z�Vɴa�N������%�$���^m�ngGғ��B)���7��|F�*�}OTd�t"�������U�~Y�L[̂��
bx�������Fea��}��c�'s�o2rAV�b�j0�zN^��.}vz�Z�^��WU�^o�o�9~�h��=�Ŗ���N��.�Ƀi�
6m�"����P��͜�T�dp>ht�#�j�9���:�˔:1*UsƜТ{,�dqh�/c��u��d�^��-��߬S��|c���<}���*3���u��y~&����˷��h���d�F<P��p�y��?g�k���
��}�J���36P��T�XGk���z��҅IT}V'ٱ{��{Q
�`��8���JT�H�۪q
���]n�<2�������6P�J"zb�J�hɪ�4"��y��h��~��E�hdXWx-��8/͙�?^
gm\Z�����<��D��,�;����@e�
��kն} ��C���F3p\�|��}k�]Jku��D�"�Ќ/�8�����D����{�ucf������EIԽOE�d�Xx6�~C����I���T�~N����`�� vCz�-�-� *�0�s��Mf�3��Ѩ*<���4�}�G���j0}h;�+>&�Y�1���2g6g��M�$�0{*��U�ؕ��W����m�I����9��0Q�	p�)�z��{����d�m{\�b�u�d^�?�\=y�N��B�����d،F�m�� H���?�P���Pa�J������cw��ۦ���J3�%k`Ɓ����5�|"�U򠛨srqY�����Sa��C*�XCnN�qލ%�Sa�+�#�!�S9
�(hgo ��f�����d&�J��+��8�OE�Jwn�}�Hb����� �<0�����0����N����U�#�m�d?����[G�d	��g -�h����Ro�Sv�I[���i���0�`秈0��	A��y@�B8!���qI���|ż���M���Ȼ<�[�`k*[Ɍ�D��Y�U)��a�$���	�����,o?�!��s�"W�Sr���4	��SB���9�%�c:��x�[����zqX�?j���Z��u��st_^ ��q�.�> ��dE�*�'|sm��,�r�$k���d��hNW���u��&��/�}�o>�3	@[����R���]fmK��}8��N��ʊܚ����p@>�[FF�:�Rb�Hd�#�=��AQ	%�8���g�	��]��s����GB4�����=�0٘�TC!��t�t.M]���h�Q%dխB���_�Ӛ&
��V8m��5��;l��#� #-\u_+��s�S��k<�*:-(kIH?�X��6^���|�)�x�b'�t�y�lf�Io��9���q�HD-b��Ӛ��F�z�v�eAN�f��8vf��yR� �,�~}b4S4g0^*��,$``j7��g��F�Ԉ�s�e��i�G�h�}$/C��f>EB��s�F���-�a������c�;">�8�o��))�H���i^8޷��{��\�ڴ�'�3��G�������^�z%1&BVvE�n�Bb	���6{.C��T|�i�w�Q�pP��v��M������gyX��F��(A8��Shŭ��^˲F�Qtp��%=��Կ7&(�,�=���5�*�Em	�����h�}u�0�b?��yU�d��^T���g�L�Oíl"t��J둷���\�k�1e�w�;��q�S�=�\f��ʹ�ś�KG��Q�ҫ��t )��8���^&� 0���a�js�z�}J���=�&G���]�&"Zm���?�T]Z��@c���m~���{A ,"6Ӟ��s�'Ԙ���;����q�+|[�4bެ- n�]�'́����s_:?ǋa����k����iB�ou.�o�Q��X+�* �CX�Î����<7x�O�8�ld��X����M�� )w��D���/�7~#�>�|�W���~�n/�Rb?���=M�jt?����7�f�@�e�����䪖籚<Y���-K#��P�e� ,�?�#Xm�=M���U��`�s�}W'D(4b��Y��|��'Ѣ~�	�H���32���3Co"FPSHe�����a�6*b�5�M}Vj��k-�K.#��;�P��L�-�P�C�YN]
lʌ67��6�g�{�[�L�ﺻbG�}����:�c+#
��H�	d�v�$q�!L6��9����yx�Wi�A��՘�����0������L$=N���Z�֣�:�j�K)�� ���p�|��G���]��(@+�۶Oo'����Ƥ���`���u���� �4w�_\+r$T��Qw���=�����˿,��W���f;؋��!��4�bBHu;t��S�	A6;��g�]����NG��܊<�a���:^���%'Ш��^�6ݻ�	�&?�	VК-��/]`J����"il�:8�7�b��rXE@�(�->�m\[����R��i��i��HE�D���s���~M56�6�9+�����U`�*W�AL�O�����T'�D���q�vs{\�b��.�4���E�b����=�mD޴�"���0 q%J���8�<��\<ݧ�ۤ9�d���݉���e3k�����9{:`"I$����Ț&��7`��;���d2i-���L�M	�e�$2�q�os��a@�[b�K����00�3r�$�/�C��=B�K�D��r��h��r'	S5c��mn�d�m�{c�Op�9Xb�1T�*�9QV`�-�ƽ�S�=����eW��!wͰ�A�r$��Ʒ�x���Wuzg�EP��j��:�X���a�m�O�{z�;�����8ۗ�wk<IR���0����(VM%H�m+Sך��O輴�j�sW8�ۡ~J��ܾ)
(�&7 #��~�eI[���ע�K��r���+'0�\|`㷂�@�9���!h ��I��޲,�6W�Փ�����dD�pY�>��B�u�+-�:�����nl��ܜirNT����������R
���3EWh	Xa�޼�<�*�|�u6�sT�\L���@����9�+����U<E�"~�'҆���O����V���l}�P��o��2?�|<10��������j�A�����K���	p��cJa������<����7��;�
H��R��,���s�#�՗n]��5�"	�y�+P�$�$�ɼ�Mz$�m�z?��]��:YMo��5�O�K(�E��n�)��[֣��9�Dw֝�"٥����:>����TU+ �zD�O�V��4�ڍԙT	m`u��h)��J�oBJ}��0��vc�*��d�(M=����;'��LJ�Q���x�����:�rq�5�lL�PN��ܸ�v��ϳ�ƂJ NS��|9m�����QQ�3���/;֤���>����셬�drvg����)��j4f�Ji�F~ʑ�X�����
�#����LV�關�?Vo���+�M<����ȫ�)��&�Ȼ}�����@ŀ<�Yd�c�`p�x��!�%���g��^�|"2}�{(��p_1�T ���v����H�1-l-d���]�w&G�����_jn��l*��t�_�c�h{��}�R�� �4���":�XW��>/�h!B�쐜gG;�"~�v�"p�9���Qn'�3_��Ǉς��H͜�-�c4���R����^o#[�"9r�G�G�3����7G��q�n�ζ����v�|��[n�Ù2�h�J�6Սy��LĬg�oq�� ��\dD������vs1�l���F�0�~��b������zSM�_j,ToPw����6�&<�?�.���,Z�1x"�M�޿��xԣf�3�OM|-'��6���x�@�I���bu�!]���b�f��n��&���������y�3��ϲ'K>��0�"~+��=�M��t-n���1�~OgE�)�L�s��%X�z��n�T�b��qk��{��jҫ�@�H�b��︂��f����Aʬd�r�WaG(�3CMUAv�0����
5~�J�k��܆^y_;BU�/��H��;�ti�rϐ�Q����R.BT��#7�9�[�z�N�VV(y$��X`an8���*f���m偿#?=��aKq�6o����d�-q�ꛙ�M'Q��Jq��{z�`y���HnUaT�=��ZRd��"uAs���ES�W�] UQ�ۇ�+X���S�kN�SS��XM6�Y��$ Oc������"�f��y�߇6+a������qU�=^|"X��,	4 ����-�����/g��-p˔��l� �m!����ת5��� Л�W�h�xyq�31p�ڗ�><�6�ٖ��]���9=JgӚѦ�"Ct�!{���l��Mmֽ?�ְ�5H��Tzn��Ѱ>�5�s-ǝ!Z�M� k�������A`�sk�g����*��C4�Wj�J�۪�`�{�lm�_E�G�31�݌.Z@ �Ƙ�1ưֈ �yM�!i$D���	?�e8��]fȉk�d�cmJ�0{����(��â#r�g�*N$�~��7'��A�w{)�?gaɁh9�.�<�q x
�y��餏����Vw�k#�SO��y�/���Q����c��>#��RoH�7s�/Q�MB�x�B�W2�����,�o����-�!���'jE���2��u��v�1�g	{򎪄��/�/tĈE�apR;7�*���9���|�%���f"	���?�+��C�F�oƗTd(����x#�p��/�N����s�BV�H��\mH�E�N�SS��,�Q�`��ݡ�ñ��p�DU)'��{r��̩���_l�C���E��������"7I�Z�s? 
O�Zb���!iFc@1lWR�<Z�W�b� ����O�&���pa7�]�����"�߬����+�;�V6�v+��a���w��/�O�?�Z {�B:_�7�<�oG����fsSЁ�ro����Z-)

�2�M�|�!_F$��|,� ��Ś��a��D�
��=檣�>2����$�m�#o7~�ݦ�4��ƙӚ�gr�u9|���]�E]-8݈Ǵ� �A��J�R~"U�h�4_X��M�bNJɌ����H̵��f�s���&�0z�ׯ���X� k�ɪQ|wƭg�դ]��#���� �6JM���U[CN����B�@��Y�af�ݍd�0�M\j�^v����n���}�	������5����%�*LtB4�0[i�I�H���Ӳ�\*ќ4֋Y+�I���ap��ɼ'8��S�na�W>�����7QŶ��F��~�FOW��@dv�ϡε��f�����qڬò`i�l6w�8.���ی�5l$���+��F��wӪ�=�J/'ZI�����,���:��H��({EL��f�sI�'����ܩ���u� �~����j�{�u�a��75�f3,�Z��n��st+#�l��H�Ki����}�c7.�rR���ߜab!���T?1��̜���'�� 30`��].�V���$��L�G5�p�� f�����}��1*=Qw�~����b��`L��B���n=D[�4���X�0{�f_��gxƽ_�<�����Q*�8N!����EVU/�4B�%�����I�ח(��T��l�"����
|�x���r�'���ϯn�A� �>3)�`�������cȵ���Y�Ue���$�"�D�k͟\�co��M�1$]�#J;=��������&�z���m�Bߌu��.���|����,�J�V����Q�������s�_h�!����N�A�r$�꣝�xDJ^Ck7��m��5��c�"= z��9~�p�iš���@���;_��6�ü��50Ótv�~�k��� �p�PtC�6�`�K� �Ss�z7Ӆ�$#�+�zLd��j�:YIP��Ex�í�|����X���v�h�"��a��;� V��+2r���%���^��W��,[(��\��"��$����e�Eʵ倖Fe8���� �	4�Z�>+�9- p�J���5��3ѭ��h�jY��9��6!P�����Jзp?��i��%_�er.:��)6�J�)a�������\��#��6��&�@��,S(p4�n1U'�e^&v
��bM�7JV��!�%���Oīs���F����y��zg?��ӯ�ef�y{�VU�7�	�t8w|u<7IR��*n��6��&��O��LM3^����N�%�j��VT]�9*��݇8�V������R��?CP�BXJ~�P�͔�"0=et2N
kMeQG�%L�������I��x9�ٶ�"ʱH,���6fFs��!�5��K��h������	}d���٘�ݖ3�咾:мL�;<�,���������?�8Gi���|�V2�L^pȅ5�n�x�5�k�(s���F��NZ5��M�v�xҢT���ͥ��_��b�PNW��c��s(e)�e�&��P��?�P
������	z$֭ߺŶ���!s�[Ѕ[���0)�g2�>���.ث�����,+��{�a���'7�?�֊zx�}�`���.�<7g�q� �qSs�S�<'��t��Q�^�ޠꦐ�h@�lho��.��>�6��i���L������:�:��gVJ8]f߃���� �S�`S���U���eB��a�O_a�?���k
���b�E؟1�5]"��W9�W�Es��+� I�P{ 2���*�DP��4*K6喨���7���7-)��[	��~_z��)a�C~� r���A ���]J3S��`��T6��V�;���'1��0�8Sf�����R�t�f����C��q�'J��M�:�a�.�o�X�615/8����|@{֩���-)�S��эN[�տ��)r,��E���y�ϝ��|��p���@�HN���A�r�S3��:��g���d`#�)F�i�N�mi�1�!���f�����Jݗc-�p�1��@� ֏��ir�B�*k�k>N�/�����ո���5!�P��{ˡRn�F�=/
`�$h+J=��1B6���
�-Ħ~b8C��ʯx+���F�ֹ;1�|�I���,���`upDY�۵N3�a-1]k'�1���p1����}�{=1��i�զ�=�w���2pMa�e���F������mȎQ�U[lt��PQ���vT�g�K�L.�/��̌Z_��A�
�Co@�[5���C��,�N��e�v:��ުNdD�~\���	�0Ö�	7�Ҏ��;>�'���p�;fQ4ϖ߻7�U� �"�$�����>��L����	~+x�)!�} b��c��CF��AŚ�ps+��8���w]wz�܇����BT�XY�h�� 2��7�8��񋭷�/���?�w�	�%�O�Z�g���9�E0m	�a��I��G��j�!����k<0���_�l��^�].N�~p�N��讌P_��TW����W�qjL�G���m	1��Pe���D�~:���T�7���2/6ި����SB^�̽{�'da�.���ߢ��)���7��C#Ȉ`?�O�o�"�e��8�����s��0�]d�\^6���J�b2R��)X���!Rl���y(���p��d�n�p�!KG
Z����
V�j��̱��Wg���(�F�6��8pݒ�N֭F #OO���W������K�{R�A�{��_���x�"��K�2����F���#�2��� �*@9J��0W/K߈뙘��W��6�*v�Ҍ�uI*͛>�0w&��)�.�`h�	��4g@���+�{�V�dqo���CUm�-i?c<i�m��PO{ ���?q����!E��Ӵ��]W�%IQx���~^�	�lvJ�����`��پ��Rو��'�R���*fZ���1�*sDu)yt�|��?T�}o�D��f%��30^wZ Tx���O;
�� n��ң��7?5)|i=XeV���G�E�xd��Z�������L5��"��
�#@H�r}���D@9��i��;ա�B�=��M�p�S���z`�̭��m�_ƣ ����{�S�m��_Q<�\����f�{E5��Rl���6���0ĳ/Y6/B+Ydg�:�X�f��{��\�sQ�l���8��=�9���?:�9�`�	���;� �I��r]�U���Nmj��An�
�_��JSs�$\@���x�� f����13�10�T��Oc L��(87h������!m�m�^��x]�u���`�dN@IR�@�q��q���w2��Hx�$?T�� ��DO,ȖUP5������|'�f�oW�*�\�)6�A.t�ԁ�;���X���;h�(��_
_(�:o��;�7kgZ�ɷs�����Ru:��
��1<��W��.�0�}��;o��U_Iej~{0������z���)}	+��y5���T՚]�p�)68-,��������yc���[p��>�>\����VR�5�O$���4O�7x�>������߭�����I��t��5�d�Su9$���_�1��٤���	[���,3ћ48���������	����S�!Il0�[�z�4��q	�Sq���F�ξk6_p��nҺ�2Gz`����V��,l:���jޒ1�� )�.��p����}�����=����ۉU�; G�n�|vk�qI�x��i��F�:�m���2�B��Z8d+�V�߾2��\�-����	�qx�������F�.^��X������(��q��Ϩ��i6#�� ���J��+�o�iJ����@��$իNL�m(f7��<�/��M6H�v��E�/�-n\��%��9i?7_�dw�ӳ��7F�m��atR�[,�xSG�����6�J�HNb��g���bo�A�~S�LEjCo�d6��t]k��3�W���6���yS�t*�`�(UrD�me�����r����4R��*���/2��GS-�wwJݒCC�e���m+����s^��c&�<Ҹ�Ai���<�1���bs�)-�H���\�p]Ǧ_�_ŀC#N�L���r��[�/Qu�]�����Gx�`��
5��;O���k��g�?v�0S2Y��ڟ����ԙ����I��A����zh��~���L\[<x���+y����8 z's8������ڿ���/�L���M��pv�ϞuҐ���˰k- ��O;U���|�.	�����7p�xB� �.̒4�*"��.�H#�kSщ��ٿ-Z�Tx4����|�q0k,�X���_�UW?\�fL|��sSњ5[����C�@]#�{^�G;md��%��������:%F�e��K���"�.t�߷^}gwUc�e�*B�<@�<�m�H�x���O8{�/�$�9����S�6���G$.&����%g�?�7����EaP�a6��7s�rR�8%��=�r�����l�kS��<��1Ϲ�m�){�- �Fd
�Y&������ӈ����%�q�]R�+��z��G��uQ.�b�L�>����F=��Z1����W�Q2.��~X2�`_��P;�8�"��
O��j�|�хF���^<(}��X�R�8�!|��6�6;��  ����E�Hݩ~}����Ӊ��"��7ޘ� �S��^>1��6P�{[�Sf[$쵾l5s�JL�r�!,E����nW]
�Q���X	�b�F�Q���Ӥz�/+t��?*V�b?��
��Q(ᄼ���O��Ī]=ԬɆH��/%&��C������6�{�i3u*L+ ��e&f�/+LI�Acq�vC���{s|���U?�K:UgTv��* iZQ:��d�X��*�hO��7�B���QVݒ�U�j�	����t�|�?���@��ڕ��ɗ��@��GG�K|��t�Y��A>zܘ����[z��&��U�9'6M�:+@jex,b^��.��
�������2x:f#�$b:E�������p4��}��ý�\D�97��@j�tN�~Emz�����ܥ�|��O�)1�\0�kV������Cؔ�_�\IFZ����������p=�x�&A���a�W���<e']7kա���
�}��C�!��ǲ��D�C�ڝ��LD����m��b�Ҁxq��7K���x���9_��!�4�x�atfy��>�p�A���h����+{���r��\��ýf�s�`�7#��	���>6�����#�[W�c��ɟ�E.��앶�0�!.�>��4T��v[$v:/����9�E�mvEl���ǘ@��+u����ѽ7',L���s�m���(��'��P?ιr�g��q�T��7^�,�Y�����c!T�?��e-���Bt��;���V�$��>�JD�Vs�{��0H��3���f5Vn{(WO�L�}�������4 (�/�k{��� ���`�I[��|���z��ɘY���v,['FnF?W�[C��S�ɰ��� ��H"}��l+�d���0�<Xg8��1�<RC%v�����z��9�s@:*�km��w"��⑸y�8��