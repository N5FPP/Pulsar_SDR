��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY�5����p}�"�,]���]'������l����Ym��ݞ�$�(Y��aj'2���2��6��aF��,��:>r����P���Ⱥ�i�q����n5w1��<I�c�d��+�6��>E�ɝ@k5����	�pkfȴ8D�VJ��b���H�=�	E��`��'�e�&[l�ٮ<pX���/����bˢ�e����a|4-/&��.�^���k�a�5��� �b�|��f����B�\��mo�(<C^�e�µ��(��_��#k�z@>�����	V>������"a��iP��an��wm�y!Wm)u���-�$�=[���M�4NG��@�=��x�mN>0��oS�x�S��U=�Y�+�w7���t<�1���KR�� �u�,[�aީ��v��T��V��5pH11K<73�C��MbԊ{45���Bb�A~���I/��F�?pLy������3a��J"n� +��w*D�&*(�pJ�h������8A\��2�9i��d�\]�?�n6�-۟�h=�O��wQ�g��w�2 ����d���J�J2��]����v�!�tm?fu����<�4"=���H�����?�i�FZ��юG�3�B��;Y�G1���D��^w��Ly_����6Y~�z�ȱ��3�7�b�$�B
.��YH����Dbι�#kQ������9�89�k�f��<�ֱj���ŕ�r��k�:��G�)��"~��cFJ�� 'bc�]��hs	K�&�Hu˖yp%I���~V[�����l�u�L��<�3�({��A�����8GM�DG�@]C�z��W?�i%�ȒY����ΐxO��xy�О��2y�/�<;��ў�u�[��}��J8�`�I�����w\b��,��0�%mF���Ug;f�tS�XW�������U!x����ڈiE�=��kLQ=Z|�9u骭!�z��e �#���c1C�k�rhu��2\�'�b�{
�Y� Μ}��*n�7g�Y��p�6��L�.��gK���]+�l~�.Of���s�g�Np#��z�47Ym�h�]��ͬZ����k����;S�;��@�|fMJP��y��+i�r��:�Sl$���wetg�V͐��bDX=���/�7Ax��횸���~�����lk�rx�t%�&\X&(\�3-�f��`�l&�D�̿}p��{�ܲ_���9)�E�D��i�e�����p�pa\�a�-��Z&jXQ(���c��������������x���F��,@�pӮ�)X����~�2���χ WW{��ښk��J#�RW�_�}�*��;���|̅��ߩlϕ�0. ���!M��6��Q��|O�,E�Ä�����Gd��v/�"�(�6<ftV��9]�.���b�g���.4:4��.���]��.�"�0���T�T:R\�����aaӫ�{cw[��=�uə^n����7L�S0i"sc6	?�_ku�ٙ\g����d��d�m����#�6f��5|��[Rr������,؟��O��0��zc�Ŕ-	��J"����
��x���0�N�s�/��).�W n���}�sI�� �x���*�f����z�Nl:��ӖbNI�p��_;g�m>�ݩ�l��]�yJ�����3̔�j�������t��� ��WY���9]>�>�	["\�]hN�������sڭ�D��j�����i�񭆮��AgOe��	u�Mk9Pe�k�֢{�C�'�"�!b�w��b��{J�HAsS�����uDb����>���ó��Rh��ŗ3[{���Lƃ������C�!*E'��?`�@�p���ONR~r�����g[s�9�Ĩ�
�1a����b 5;�]�w�q�L�O���rsSXG"����s�'��t�M���#�ׇۻ�/�A�&ݓ 7��-[>b�esy AY�5g�{���\-tQ}C���EWЖ<ts`��(�=;���|Q�W�5��[�]=9;j�_��q|��nD�I�<|��
��|��UXo��&M�K���*��"�1���M��f��Ynm� EfBetċ;���n2:���Q?�#v���5�'kx����}���43Cg��X)����9��3*eg��U:�g�J4�$����ӧH)Nf_~�)lL�γ�qК����4V6b�]��4:�?������h"�pu2��W�x���[���	��nQ�!1�B���vTD��
�TVܓ����UW���b��a�m)�%y�A���� �նÙ�..��s^�F�\�:�).�4����\�N��ț�wӋ�ޣtbo�,����1��J}��Y��5�W�L���0��I�|odg�;������b��B�4s����Ȝy�2�81�K>0���E�X<�f\�|��:�i��4���ɱ��]�oS�G�N����n]e���
 ��
\��N���b��i3��9��V�/a����2{�����KM83T0���l�:ǲuodt�n�~Fa(&�T3�_x�R�<\_���"�]?���?�_f9E�D�Ќ����77w�|4�r5�RY�:����q��L8�6O��3�-2/끁��4����� ��X�y�H&��͖��!��;��!��ʏǉ�a�1~3$�-�
ĴT	U��Av�J��Y2Hl�����(ss� �Ŗ�t�w���Ɣ�� ���r��^��4�g񌒁h��C
���A��Є�<M�h<����9:��egQ>@I>�_�����\��v����+�8��?��9������E׉�7&BMX=:Zk5-����f��t�_&~�P����{J�q�N��W^��K�2C�&�>�V-Dlujg˥D���'!�y���-vBl�n]�M�$�dsÈ?(�sR���y�R�'���$�S��Lr�⃼D��@��G����~]��0�H-�A���m����@O:Њ8��<� 0��!j���Me=�ܥ�H>���z[������t�����}�����;�ƞo�!��Qo�ȧ��ú����ƓiZ�V��ovtJ�����7�M�9�����>�/��Q] c�H˭�eC�0Fh��UD���0+�����j��jJ9'�eV��=T�	��lw�K����'h2ĉ̚�[��g�o\�4ޙ�	$b4��������X�iz �4d,�NJ���w�� [���#l�1��m9��2�
�m��T�h��Q����I �I��'�\��7��]�g��ө�
����q�j;�X� $�;Xnŀ�(װxu�cV�+` �����v�w�1����>C &B\�b�F����Hi��^��mlɋ�1�9�M �ETo�׺��dWC����w���&���H�#��4kr92|�s�FTc����.}9��p�1�PFd�L;B�,���G��辖 Q�E��q������A��"��4;�g�6z=��`#���9���j���G�Q�{ۊ��J�d;BW����){��*�+J�y�Mq7a5o��"V�Ӡz�m��i��^���Z��|iPϦ��՜I��,�害��y*齔��
Ӳ�{�c
X=]ŋ����|b���2/K6G�A�5��>0[.���L���=����$��\����,&ǯ��Xi^�5_�Qt�#;�+/�ً��������`ˢw�q�Z�&6;oV�Y�Ҳ�rz.2F+�2��I
�az&���˜��jXh���1�����oE���7o��R;bx��n�f��8[��i-��W��������CTu�$�<������Z�z�!_�a&~F��K���V҆VKŀ�,�EA���<�#Ns1���c�����aEva�3�V� IG\�����p�S��9e�U�s�ͺ������(s�a��@xUӸ��<6CW�k7�� ���T�H������=Gs@Ѭ�*6����� �'�}T�D-�*��DA���:�e��]FT(�RJ��\��l!�O,F``���:ҩ�j)/��;�s ~�x�uߣ	���M�7��x�{9 ��V&��Z�gs�*�3b���p��ߓ��u��He��Mն[����b���f��j]G���ء�Tn�5�lc���j��SBF�@�z6}�;��m�S�@Z���^��V��h��%�U�d�Ʌ���h���v~.7�Wp2:�W�8����^��&�����|�S-�[8sW���_�y�R��I�Q�=�L��^�0<����yC�T1�"���v��|P[�
E"�>�@G��׌;������g�5�:���U�^%J�"�D{�����d�W�_Y���Cp؄:����k�����_b��_�C�E�~�����JJ*�gOl�Fʍ���<o��8x}���~4�@��4���S;J����"a��;2%imH��o��ٚ�ɂfP0�,��(Xa5L��� ��ArHhFfY)��	T�Սb��}���{n8�\�����1t�~|�������挾�~"�ڵ�7v?v�}N��߸�$Yۘ����ͽU@����m��W+���ay�_v��2����b�qo3��R_���_�|9��I�}����� y������{��o����%�J�S�YȞ�)]����P��)�A{l�8�m����y� �LH���Ի����+�h�r1��WKpk�ğs�+K�_���2�8��	:W�O���F~�`m��QL���Ύ�1y"7~�{����r�]TZe^��)�1�>�_G�&C-`�>�����/���f)�7���wq=��t�b��Up����o��"�*�W0��zh�S1ږ����u ��5�#Y0S�8��ҋ��z�b�5ד"��}�dy�����8Ehv�G�ܿ�ZI�G~�����TX�v�ҟ���ϵJ��O�[LZu�J�W�#8�8ߦdː��\��4`�78rp7�5����ѭ�`�����G��t�L�h�,J���gp\��JЀ�|����=����R��QT�5B4h ���0R'�1l���Ƒ=�zq9)Q�w��Ұ�n�^���jH�Z�WM�'\�I�4�� ����q���xch���!{ŕ7����}s��#��e���6#�s�▢�-
����e�;^��sAYZ GMc�D� �'hJ��4��@i�m{j��O��	=�Q���Ge�cN,L��\��_"�f�q�>�R��R�L����rH�R
(��X�?�̚,�W]�����(Cq�2�(�p޲��rgyj���Zm�<��ضf��ބ�q���*�4�zɴ[8�H�Οrw3Rl���W��`�����D�ց ��%��� 7Շ�md��R��a7н&��ie��c�U���@�~Sڻ��Z]mh���C�]���m鏯��F�TFW��"q+P����@����ɚ�ؕ1��ӷ�1*����l%�R���\F&��v�x���ք󄑶�է������m*�t"�f���Ø>��hH��1� W:�F���S7S�� �PЏ�@oU�U��#�1�r�d8XբXҴûٝ�����ټ2M�O�q+&�����h�P�q���r���:L�߼�W���
���фƏ_��|�M�e��k��XD�A�4��;o�dG�
4~`kU7P6h���Sm3�{�x�#�0�����0��H#2�X���G8���xtp��u3v�F����������*>pצ��4���>���X�m���| 
�5�6�g�B�Ǆ@L،<l��yє0�%eA��,t��)e��]:�{�~�*ت��\ Ӝ�#٦��fE��X���ˡ�$���#�|�'���w��������3���*��g�f�t*ª\���'G#�v��Q�	�"��mG��ޟ/��9��Ӡ> +p�Ѡ�Q�w P��rK�[ EJ�i�X�6���8��� T��׎���	Ɉ�d���j����x��H���U+�(��c~_����ɪZ�u�V	0(��������%��^(�\��1�ݩ�Ʒ��^j������Y���EF����KGݩ�F8E�n�i[��1V�iȐRB{���v��A���}4�,�x�ˏ�Ѧ_�p[a\�x��	�j��6�݉W%��L��H�H;����PD`G��j��Fw4��NF�;g��|)2����y8��H�	��^+; ����?����>��W��J�Ag:���*�cC���ă��j��_ < Ǥ��Z
�3z�9T�&��/q�<f��Vk�ʜ��omC ����չ�� ����.��Y���pT��^KA�	ޠ���0ӕ�!P@�Gg����i�&p�a��	�|m��w&=��4����Ɉ�Mpz�;
�c]���}{��p���ݏQ��"V�^F�M:j���4������7w�h!w�=[`���AYN��X�Y̮ۘ�iա��v��`�O�L/�f�wc`H�a_Ww��������#�cq�D��@��/��5b���?;s��E>N�͡�s���j��C,���zYO��wǠ�)	�K?ތ|R�WD��<��9/�_{��X�)�{]�)!}"�-�������Y{����������x2`?�.�U�����x���hN�ù��X)ǭO��u�X��S脩��r�\��.�e�O ��jܾ������濭�Yh��BY�ڲ�w��#�V�H�H����%�����~��$���,�]�fq ��>A��������.S����<��r�2̣�wD�:�US|')�ӑ6��=`Q�r/�(}>� y�Q� �i �$PV[�,�_���:��N��}��?�*О����h��Y�ua)��a�s�����?k�B���a����I�a^�x!��e"�P���{�%����ΚxXr.Jy��p3�?���?o��-"๑ځg�2�T�̾�
���(�W\+T�ۀ�c�Q��w����Gv���co�媩]5�h���3rp�P��NN���M'�_q]q��:���A�_D����#A��4'��.T8���oA6R��s���elMgcD"��D���Z6���4�{B��wv�!5���z�Ωvʅ
�%TN�eXYI!k�=�c%a~���T���Ȉ��]˝�YLtէ�3��Zo*�{���Z'9�������9\8)܃��F�|���ĂX�IĐ�����iy Sg�UWm�k�Q�&��v̙LV0��`b��ܱ�v�%�����'��WH�)�FA���)���a6��u�8:��S��F���~��C� I}baԟ܋�<c���)��M�����!{g����dI�~$uhΈ$�a��{� [P��&��,rm�"pt���hv�P�3hU:��J�aQ�V�2�ևJ�%��>����ne�K��U?���t�������]-�	z�����P�F��በMc�P�K. ���1s�ǭ��j��9ôxh��Rg��^A`r��������eŇ��!�
4�L�ÿ�*�.��[�u� r��+�;<׉��� ��W����岇�F�zՌ'џ�HNy��u�2�b ��$w��j���O偼e��cGMG��/	�xW(s��Ύ���=���KV�4�d�R��������P��R�M]P�6 e�Wx��$^=����Ǌ�����s.e�zFb��XEr�4^5�����; �W�=w�01D9��&��&�Q���v���#���%�H@:��&��*� ć�˷����l00�T3_¼�As那���UzeG�(�ZUM��Ü|����M��kg.о
p��?�J�54C�4��%clM����qᖦnz�΅�]��~�JJ�����$.�!x��k҈�~�H�
Н�WM�S;��*�e�^3�亶�Itr�(!X�~���)a*�c��tʹ5s|_�����s�F��ϲ��Dw�c�|S���o�(;����1�d��L��Nx�D>,�Vbm�ga���DU$d���-v*�f�հ�q}����2��D�2�d!��(4l�P|�؜�Ø��`�n]�y�"�����c^Q� I������T���a?��1/B��le����i�r�����=���WSm���Z����A�P��z�{��H�^-y�fӫҒ�����ږV��	w��e�w���RG����9��m���6�2/�N�C����
�0�?��op�ůx;Wxo(H:��i�"����@r���f�态!���jԪ=�D���\�2����.%�i0.=TXo��H�L4-�H�u+�b����c�	������$D���]2E��>m�B9�Gy������{�M��h����w�"iҕ�pwߡP#UE�!}���qwh���ū�B�C�J����	Aw�q�+w䧋�����*B��Kbd;H��)U!��`Z��{d��-�����[Ο�+�L���1��VjO���=W����g�+y�Ԅ�F�s}l��g�Y!��N\v
j�����;*8�1��Ob�i�v(N�t�pY)�<sU!����d�ۼ�!C��:��-1���i�ϋV
΀!�3�9���P��mmgoV��[A\���X۴׻3�'F滄~}���Y�@�7��h�^�������
�G?�����u<̇���'�����j/���%��!vZ�F��u���}l��K5}<���k+������B���T�(��A�J�����h����9i&��t<�_LmK������[a��ڦ4ދ�q�2(� Uɱ����LY�,t��J*�V� ��L�S͎h�d	�3G��nѽ�Љ]<� 8�R�s��_(yHۛ��n���ߣ�,��7
hF��XP+�K�ɜ�g'�,�a�P O}�����*D�̐o斄��crtf�l��p4ղ�i�,m�!��{��͘�j�[=N�~�-#�0��Xd&l@��GB��lo+O,KW �d�B��U�;t�5?A\K���Mۯ����kLi�����˯'�'m���>�2T��|������C�y�|��2������y����ʼ�2B�,��Z&�03E�f����u���x���%�UԱ���=�90�0p��������vDuRE`Z�q�F��P�N����H���b�Cs�mIџ�FYgto`�"�K�>��0Hٰ�`$q�"�����;��������2��Q�t���i����E�Rg��1?Bc����9)�v�ά�fN�Pkn���~�z�ѿO���'k��cƍ�T'O2�㽖M�M�
*ƌ%Eu��]���� �V@FG��� �����f���~[�jkj&i?�m�yO�%QIL�z��l��f�Xע���5�_%��E��7��'�	�"6U�xx=�l�1��m)�.����x���R��򙷊SG�P{�]J5���_�ڮ} �,w��/�q3ܞ����˛�B[��5Y�$H�͜.J8�]_#↲�E�?�	7����Q�� �纫q��^*DX�K8��0��%tD�oM��hO��Kw֓��vGT�M�Y@_�0�`k���Q|��Iy�H�n����BJ�*���-=r��^!;lN��#��h���,�X�[=�E'��gZ�zo�_�����X�t����'{��=���tH椭7%��� ���0��M6�������}��G"b����mVPW��K�^�K�ۀ�_�p9���WkI��JD{6w�H�N�8XM\��dɭS1�8\�P:�˖(��0J7{�2=�f��o13؉G�����I:udY�'���5!������URR���?�ׯ"(��c��O�-����������M1jc�D朡��ނ7Ɖ�2i�7�`�~���J6<J�QK�劽���H����;�))�,ʣ˼��Ɲ�}b��&�ȅ�fG�~��a~�e%�)�����:�p����?M�ͽ��K(=���F>W?&/�@py��1f�A
jy�1���i;�7���'N���y�^Ϲ��h�.i`����B<r��$���� �$��o�}�Bf]���z\lTz�\c1a(I�
��N�&/�A��5L�ɞ^X��	X,j�I��ո�v�n�dZ�y��c*-*�\���M��xj��ϖ,�
+|��S/E\�w�. r���g*��*�Vv�9|��N���Z�ٽD���u�bkqVN0@&ȀO����U:��q�\�h�C	 "���NH��AQ�	��,��2��Vbt�a�[}n������NE�݇9�Um�82�֚������7�\j�L�����@	
?VGwR��4dn�>�ڡw�`t�n:��BZj�{�X��[qK���n|�Mb��D��,�:����v��yp��q����1�9aP")��ݜ
�Ue0P��
eY�*�6p�&z���a����h�>����j�'�Φ��E3�D�k�ي�#�2�.������*�M�t�Q�o�`�3湼5da�>=�	��퀂�TݶG�޹��JO�fw�[�
pbDb�h�HǛ�QC����]dGR>9�}�N�:�'d���Z�d�{i����ǱAv�.�.������S�6� �����IA>)��G� &���9��ā���=7U_gW'PIq��Eҿ?^���G<�%&�ƕ�ڣf��Y��l��P�D&c ~?����#��Y�)���p�q�|��>A�$a�0��N�{ ��w�C�'F�v;0L�@�gx�)%<�V���Ru:�\��V�o��`D-ɠ4�PoYCߧ��$�S2�PA��IPd�J_~���� ��A��&:!��{�ʉ
=�L?oBP��E��1���R0�4�B��qY�����xzn��7�`ћ�fo�:s����s+f��I��я��3yt4�%���bP�޿?�9�(D�ʒ�0�D+����|ʧaͱ�]�Xve��9�K�R�kQ����Y���|��:��{�5�n4�`=����n�9��ǚ�F��^�6�րK[�.����8p�r���n>���-	�t� �Zg��~�-3�@W�/�ޑ>�������o�MP�s�Q�3q�C�%�JB&���G�����>"��!����6Fꐣ\b�lu@�Ɩ`�SL�&K y3��Zlw�0�Oo�Qܕ��Z���Q��i�uORߑ*�'��Z�B���mM0% �)刡��;��c����x�JJ��A0bڅ;�ę]��cOA�ͅ�]L�S�`��2��g3��0�6�eU��ܳO�0�3�j�t0r\��x"Zz��`����8w\���$��a0�k�e�{��98|צ�C��%Ȧ�)KT�Z�d�	;���3���$� 7m�Q���y�Vb��iM�B`���i���H��p�.zB�S� 	�O�<�Iw�*8u%9s�r��"�?��+`��P�QG�'e� �6�;b�䚴���sR]͜����I�KjR��
��0��P�uѳ)��H����XT���D>�v�xjٍI<�I/r�nɖz�e�{�P��s��T8�Z,���F+UA�w[����Q.e�����jV��i����	�x����Jj@���i*��Md�:|�S�5IT��!dG����E��I4�^����q''1�E���|R�O�C�_Y����*�U�pK �����W����N�[�$B�u�m�)i;��MM�4jA+�+��TMenN�� W�J�È�f��6#�����L�+�&n+
r�H=e�|s��Vԡ|��s�u&OӽB���`*f+����!�	����(��֒�[��=V��nt��}��ڻF�0���O�J�� �B���#g$�)�'M��s��T��"
�&ɢ��@�����R��OǓ ��A�!P;��>7��̀E|��؎�LA�x����eƲ�<k�r̫��JF0��!�Z�w�6�^��yh悰"�tU����wRGm��[w�i��N�6p�#s;r�8��^z�m
P�9<7g��]����P̤Prk�R�H0G�������&}< ����Ѧo2��_'{�f\E�	?>[���F}�JC�H���h�?�89~��Z𝶘��U*���	q^��*�Ry�.��͋l��#���q[�tV���L��R���U"��-�l2ܲ��%�aG��_�An�azB$Wn�i���+�ԍ�U�"NC�:���z�0�8��|�U��{�]tS��%K:����Rһ�y�<`B�O߼����3Ǆ"7 8{��v���$�p�jO�u��@��#|��"i��o���*E3dD�l�8`s����@��[�F-0VZ��J)�54�I���U��h[��P���k�#Y��� ����Y���� �{]y,�A(��lu^(|8m��6.h���r~E���a�����~�3;��;�����J�C*����2���Y�i?��Yˏ��ӹH���p���jx��c�}�oK�q�.�^���Y��eJ��}49*M�~�k�!kC�RL�x�U�_��N{���5�}0�P�Ⱦ.�i�����cZhٺ�8�{p����ir{�^�)\��3��@�������srOeW��C�X�!�i\���/P/�\�6{$;�,fŀ�u�Y��0¿B0���B���[<��U�W�s����[X>�n�A;�z[9g�T�G�5�)b����W�E�;���ύQ<������9 ��+�Ui#�ʾ[yI�j�f�ef|B/B4�Vи7_����3���$���t�Q:�9+
��%��ܴ��j�<2�(+ځ����q~p�j�#|4�.n