��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ���L�����I&V~u~[rR�C�XT���o����۟�V/]�@�!ӁUټ��)����؊������I�Xa-�w�H}�T0�me��|_��������M��)��H�BK���G֓�r`6��Lg�6�ދ��׌�ŵ�G�0�2�!�J��c]Mw(�C�����Af=�Эh�c��I+ݎ���O�� ��^1��0s���=9�߸K�V}9��^��*!�S�����p�QtVx]�����S`�)|e�_R ���bd���_63Y��UgN��l��"l�����I�Gɏ0�4��<vT�5���m�༇�µ�U��H��z�4�n]����-R������ބ��I>��L�� 4):E���V!����Q##^W`(�
�P�CI[q���Y�ӕ��Cp�5뿳�p�3� �agD oa��EčgF:K�=/��R��MV�ٳ P�"�:����Zk�Y �{��W��ϗ��ݟ)m�F0�XFk5 ����V�ӹ���:>�H�A_!��K�� pxH���КϿ''���H���%��?H�} VL�Wj��	[��WUt��6(2�"��M�2��d�)��*>\o�䝮6g̍�u&���;AV�{joНgl�z�-{@��oߕ�����W�S���i�f��5+��l�u�Q�vdy�-u��D�d�~�W��QX,_�_�IZ��E�]���v,Ik�5R̅<	�{�B�v�ū݄8��Nf�x�L��_��amY�A�A"���g�.��0U�8W�Y5sgVu�e��s,�	Ә�׹�+�YŅԘW2��
��n�J����}�Y>�<q,6 >hO���.����Vk%�:��j.�f�����,�u���u�̨�J?��}m�=@�N�9���;��eXK�;�s�x��ڒ�h�r�
��������ڑ��M�W.�s=U��Z���v]U\��=���t�+�(��տ;��o�>^>P���U�$��t�9� �&��.M�2^��i��jA�~Y��2Lkpo���]�?�a�]��ڣdlH�2����
M�Ȑ��(ǒ��*([�?"/	c��Ę;?E�VӋ&�׳R�T������n�R�z��l��5��Kߞ I�{��{v�o�ct�Ǽ�ɩLg�����vO�� G��#�Z���E��2=�C3��*�'����+���}�1���=ZũS)����lN;I�xת%�f~�lZ����ꧣ�|�t.�i�цY��TX�p@|=0�4�����8`ҍMh���<�]�բ�g�-�9%�]�m�V���$�����w @��Pp4o������nۃ�z��G�amqL��}F	��6���Dm�HQ~�7��霫�/�s�]-��o��*�\<Z= K�*�:�j�_�>��6c����.ͯ�D���cP�ѣ:H�})�'����+�bK�t��9���F�� �P�b'o�lx[=�����R�Ѥ�)�_~2q�Ǹ�z�b��R`0��;�㻖ؾ��̻D���i�?M(����}io����M�e%�m�q��un���포�\
oqu�Uv) �
�Z.n�~&!%��V�C�LH�`���5h@_�bWPY�4��x�!���\{5������W�U�����r�>��zA�j�3������ۍZ6�C����G�'=��(�rG��iEė�^ �RK�@JkbE���D��@�<O^����p��s��b�{{��]�v��L��t����4}R�Gi�udsc<{������0i��̫�'F�E�o"m��@R!c�z@эo�cQZ20��Nc>�P�n>n�M��jۙ���}�L��a|9��b�)�۴z#��HTrn[��BC�F�v0E�lFok�\zO� 8"T`V^C
���H�*}���A�g�CnX�9r���E�wb���؜��v���1��7#'{���b�.p�Z������a曥��� �KI�~.�~?��h��ʠk2K��(��jT����~Pc"�)h���(���?a��l���i�? �i�(��7�j���4q5�s�d|��K�3�z3 =V�d�Q@�.����m?�r���6'�`vJaK%~\��/}�-�F,�ŧL>ao�5i�-(1O:�Si���7�B��3,��T�b�ODiJ7h>����.��k:ʔg3Tv������Q�h���L1��D��}#i~��C�@8J�F�s��vf٢������no����XXux���#���v<�SL���CXS�`:�^WR�+5�a�y�\��u��p���U�c���o[�e׿�*_�]���'���uq��^��w,�P�Bu&�뛤��|�]n�ɝhi�����g��0�Ө���e��5�^U���Q�o�_uL"�X�	��K5���L��*��]8�;�J���\ˡ�eT�{8ϙ��bYd\8��b�w!���o�v�P&�����5�3�Z�  �H��x���Ҋ��������
s֦̟�(���|�3cp��i����1��L�L�ݚ�u:?��Kn><��?݉4��kS�̧�iY�<8� ��Q��ʋ.�4�1���ǌ���M>��2�Hֵ2�3�1�<��$�&���|�N��7݄"�Q��!����{�@�t��"�c)}
Om!i6H������U� ϯj�"/�UL��a|(CӴ9rZ�b���J�	�������9O�A�1-��Wc�����D���>����I��-rm�\���������r��p��&���uRT�'�,Vv*P,! ����F�@���9��o�ih�&�0˕���(��VS�	m�'�O�����wf�笂U����������2��A���O�*�H�)�{�����'(y+
���T �t��.F��3ٔ�vʁhA�F��# �b�,��+,��~���h	����hj��ZSi��,,����=c�I4����9�Lp~�'�f�>qG2s��"1��Z�vkh�C�������ᶓ[A�ҥ5���g>���Қ�F騐mG�u�p������35����dMW�a@J��Ea��x��L4�n���C� ���|2j�z�� �q��Yg3�<��N��.Ȝ*h;P�6��#v�~�!nNe���P���4.G�E�$V��_˖�{�_�A$Y1����ū���	�����d�D��)
2�Y��#غ�֤
��l=����u�I�� �����AZ��)����S�}u�үW��f��E�s:�yїs���{SZy��?�F��ę�/ui��ڶ�$R;�nHx�4���k�	(y߮=�r�D.n�Jn����m��K�6$���