��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��e�ik3�������w$����g|��J^]��sٍ�<9��uB<b~���R.�3�������w\�8�vJ��[
��~|�ɵ�v���ژ^"�/� �^�!e�4�@���e�U�j��Q��5S��	"�v�o[�.$��_�鿹��ӆ=��p�2 ���U}[N23� hȔl�O�2@���5K�tWZKW�&�p�t.�6|�<.���k�NhC�^08�+|5il|}A�ʡ�:p�uWAb����(۶�u�R'.TXF����N���Zzr��B�Cu0��I+���s�������j���莇����Ѵ��4�mfO���D�=`���:`6�5d��ϜO�	���\�S٦���j��7A��k%�����{ �+�X2}��8e�j��ef��^�ǼI�I��7��+��{ӫ�s�:�M���㊇���'��|>آ����jLg�a��E'hX_Ծ�r��[y�>��C���xæ�&v�4f�x[2��4��)���*��er*-c�o-�V����"B����k�����y��K�P糁��6-"�[\`"�G�4��4�n��p�K;��J
�{��oH�z���D�u�U3�������]_���o�E�tw�)W�OO8���~��?'���Vڭ���|@u�س'�`o[dW�� =m�+�]\�:�A�{��1�~�T�k1
ʰ����=,�zi-������z]XҶ�0�3����|liF�Fn�lH����
͘D1�R)�t��²(�J�@�0��&2a;�3K���r��rè|�������9!ɠm�U�y��|@A�6&P��ק��9��j�*�>˞`f�uZ�z��b�/�G�ɢEc�!�_S�f�˷�l'��<����%���j9b�~�!�ݢz�����D���w�@]�v��U�	�Ӷr��1���&�NǕ��si�.�3'�(��k����~�y�+լ�Mx^��[����.uT�O�X44��w|$�G��B�����[������#��&�\�GnA�y#�iqDW2�c�
p�iR�2��8]!��R����E��ǥ�?paeu��:0_e����\�X@����g,l3��j�f�(�XTg
o(�E"a	�<#:Lĝ�I���w8��`l&<�V�qHx����H7a�<)S����u��N
���c�3��ME+�}�@�q��GE,��S�[O�!�^ EG�[C.]3�{0J�J<�'��9M�io��Mц0��9�,~�%:�3��C�����g���7���h1����߃��640�0�5kšY�W�����>��a��p"`b�J���7����?dԚ�CF��@��6��a�����5����m�-h�$�/b�1�ӔV+7���x�5M��Ҫ}Jn���q��x�|ZZ�u���}��Z�^���s��]��9���4������c�hᬎ�{�Ͽ|�-�	���
�lf�χ��6q=<#o@kƉ��o��aoy�����J��ʾi�':��ǃ@]-~g�j�I�V�L�ːpђ�yϒ���(�N{MH^���\M���T�R��$���o�Ȣ�}OeZ�a�b�_�s��� n����[_��
X
�,���F��L<GE捳�+>w�X��)N�(�HGҁ��f����f�5����1�1$E�>��|N
�D̰F22��1��(�&}��3�6����n�7�߶�T;sB=Cs@ɱL_��0�v0���TyL�q��W� ����E����)xx�&}�����)[a�uzVw���r�"�V�O̾�ˋ�`�������uj3��"��.�ɰ_G2�0�(����1|�\a"������+�dkj�1V-���[�OF�4^R��g��/��J�Qb�;�$R�|x�!FlzW���w�c)�q�PTȳ�.�'�^��ǒ�..}�f�"[8�-�wk'���N���^��W��� ��`�t�6�3����J�A��¤ ����Sa��ٱ7��һ)�m�>�+���j���M��cJ)�� �� h}�9��}$���1��ϮU�tB9�3qc�4)�����`m�?{'�;��w(pB�t#B&���)�D	�q5��ϟ�%S���m����U:m%�t�o��]� ��Ҏ�����s�Ѓ̄�\B���x�o�"Yp(��n�(��!����&Ƈ���t�x��&��Mt샋C5?S�L
���4z��3�+}�1D�+s�Z���b��UPDgHe��t)ϵ�k�*��s�W�/]�`������5,^�f!����s^]�D"`A!3�T��՚�߉�_8Ks���U��c���-�MD�i`�h��U��/�(q�� ��9!������*�蚝x���*�GH�,�7=P��O����&�����__������
h�t�!��☴=�P�Dd����<���2:�|�
5�:e�z�C�/W��ZS���J�����II���ӤQ���vȅ:̵�1�g����i�ڗWܗ�����Āb��f��ߤrn������İ�}�K]�=:T�5�T��XZ�H�_����3h���nF�Q�R�
��{��A��������>��ʳbQE��kb'��Li-��Ԍ���:#1��ף,��z��T���:p8���Hh�������� �F�1�c�|��5����[~ȩ�"�J����vc����.���Fe�4�p�+�r� ��/?6�?G�b8z!5��T�>ˆn�_{ka	Yf��&�0
����D\�Qn�Ⱥ��@�2�@9t��Fڛ�1K�S.$X�-�YV�-��+�B^6˘/j0񕭾���o3��ӱ�nc�)���9}'݉�pӆ�v��	����0�$EZ�Ѡ��4�A�� ���U��-���J�����
e����C�E^�E��p���4�$����}6�-���;!��0Fæ��hY���猆�
�>��Q[ӝ����ȁ��U����2�S7�xuQ��H��VƩ|�(_�C����X�dY������9������Y�I7��܆����/Q�&�ϭ��V�F&��7�l碑lm�1��tN�%[:��"����1I� �0��, �Q���y<�0O?6쁤*�ʹ!mS���E�ob8�m�]����p�9���,L7�o9c�
���Ho�WF�z;DL��D��r�x�Hx���U��B��ٌa� h,�4�o"�ƒ�F&#^�	[KXN����T�=IL��8�Pas��ξ���Z�T5b�M���~��"�(���\%�'�Zd�;�B��/�A���]2=I�����XATz�Y+��e�O�Ϙ����6LhM�9����N���pڸ���j�P�U�Mz3�n`"n��"�����K����6
w���O�HqU�,x�T<b����	��mm��f�)йY
S�+��^��m8n���`m��7d}�RĤd�t��ne��b�m8?�!�ގ4dl��Oc�4�+R������C*�#.�5����vH�˻��]%��ZA����Kt���Dt��Os/��AȂlԝ4Iߑ��`N�8Ukp�סLi��[�Q�WN�)�1������3�D\^6$�1;�|0�NR��}{�i���IΡ�]2ʶ�X��_ĄG)6W��wg�tq{��r實����-��'.))�G#�3wɢ���8D�>��$��]�H�?f���d��s>P���m�q�`Pγ��C�)��kVϚfs�KY�s"b[|��>��>lj/%�,�~"7F�v3���u+�i����4��_�:��mq\:9�'<A��քDw���5��Uс���s�Fĵ!���^�ǫ4��ڤ���q��AN�y��2�A�e��D��lt��^�6؟@ &��?W���6���ߕ�r�G��|ēB~﯀���s�J˂Nt�X7�����?�U��9�����g�__Y��9p���稂:VD;ꋦ�~أ��(_��P�
-���������\=�R�5�k�א�K���|�j0�$$�l�6�N��"��i7j�E�j}��h�-�1 �f��ybn�Nb�
��$;���Y�ό��.�$J������jr� �c�L����F+}|�U��bz��.�lϖ�H���\����%�#|� \ǂ��9�jTc��(��^����7Ԏ�=��-6tR���UZ���"���g�a)I����fӆ��k7l��
$�˳���=G�f�Q3*F<�|��I��T���#L�Zs6!dMɀ��4{<	�SmK@���Pʾ����2���V#C$��݅�,2������66LBoЄ�!�4Z�酠���\�.�I�����6E�4F+�T�����=d�|�=Ө����n��}.�����Ym]�(;O\S�ףp�%�xh��,o�:�04Ў�+��X��ɡ�g�%�e�~#��Z�[m�)c��ҕ�.��
>xhk�H���c�
X�.����J���Z�͚_/KPk:��B	��x����q�z�&�Xi�V6x��
��1�=~(��FWJ,]�\O�n&�5�|]{vQ���T�p)2a4��.���s�ٕ
�Ki4�l§����r�O,���9h�͈'v���e_�����DN����+l��c����ޔ��Y��{�5*�<�����uV~��۠��LOh���t��kX7��d�j��$h8A#T@��l��z�ER��D#Pd?<�@�X��X��:��yԻm��KV��6wA�.1��թ� ���k|J��s���dü�;&��C�4��Y��FJ�����nj��"��� :�����"\C��:xT�3? y�g��o������JMZ�㹈%����Ļ�]è���kd2��o�-i7HZ�VL��j|�`�;ˆ��o�;=0L�g����B!R�Љ�{�+|��h����#�X�I��͋�O���X�rD��7��<�-�R8-��v��S�h�7�ƪ6�>8���\u�ڗ5�ĵ���(}p�g������$��	b��Ŧ��i)N����<Rw������@~���/��~m׎,"��wxq�3z��Z�Yr)$P��R���z�_]��kR��a�������N�� �� �[w�[�a]2A��l�8HL.c'��3��ZU�	M�Ѭ4���%���4zI�@}f��N�*���n'G�
Bsj[�{��lçzcB�C�9k�yv|a����ã��uq�c��#(�0�A◥���f�?�+�R���G�yg2�.�r0$;f��}am�����Xk�ɼ�X����d�>�}�g��4�oU��]è��~��4�jM�6�0�<�n��z� R�}-V�5��.��l���c�����J) �iJ���-U�X�&��MU��q�9�#��*���[g�;�$��
	�*Ǐ�������eyJ�Q�5������|x"=�dU�t������Q]>{d�5m�ߦ9��,z̆�V��2VKl�7{2�٥��1����`��o��cm�ʓ^x�U��+V��G�Wz�`rK�� ?��I�,�Xˌm��4�MU/?+=BG �r�vN5�����wQ���o�7��\�	h��A4轳:oQ :;�U4�������FHېI�1�398�o!�h��a��Z���wV*�9�8��<Ψ��܆���j�&��ߘ?�/������U�ri���A|�����1;��P�v���E�U(Y�D<'�t�Ia���B��$��v����0R8�X�/���9b��B�2n
Q߱�:vI.��샩����˰i���u�M��wO��1Ч���m��~t^�+7L������zp��J�q���]yu�Δ��gC\)>T	`l�����,�:�VRŪڜF#����D�Ie�s��h���V>ѷ�8�-.�&"��8�{ߣ��^EF�1��#�3zғ��[At�8��-/�/x�O9��[`�g*��+l��S����3v�]c��?���D��X�ݞ��5M���k`����Z��)��{ү�U<�5�"��NL�g/�#�G��r=��Xҏ����6G�'�}�N��To<�^�n/X�>?��m�T�����`�M����vĆK���5�5����z*do�v�����3��1`mHcX��	�w��XKMTMl��6�N�YD�2��{��E�|ി��z2�!hX�fG�\
s< �Y��tܯJ���#�63,��0���z� �d����S�j������i���b��L��Xf�����5����1�"j�̄X�

c�U���7>�x�|��Qtu߉Ƈ��],7������P�Y�-A�`O����|��yN�k�t��x��8�9[Wq���Lϥ5bb*QuT�n�`mU�>k�N�H*I��n�O86A�M);[t�g���7ڂف+,?d����F���NC��$ea�J*�j���a�L��.Y�}v�j�[QJQ���+�鞵ONA{�aWe=N�}sR���&�řb��>��nV�j��+�}�Ȃ�D���XE�w�:�a����bY=ka�3V�t��C��A?�j�!*'u�Ta�[9�뙥[4�w��J�W
�"��l.#�Y�]�_<�� @ u͜ c ��F�wq��l*��W��62���c��(P�^0�z�<�����:��y�Ktu����M�{=4
��`A�ތ�R8�hƪ#h�����0��d�ϓ��`������~n���&"�1�aa:��1|\���k��s���%�Q�H��
=�hl��-�v<X����=��ʩ2��?e����;K�^�]�~^��b^-�q�.&6
C��k��������Ht`}�4��g��`7
a�<�� �4��L���}�,��Zn�!�ѿ��J�1�L��4x��bS�L��0H�ni��;A�$�f�]9_�i�,vbq� �M|��U�� ϡ�Mx6�'em3��5�;�J{�Z,ZC�A[u1+��i����@ �` =��T!s��U��M�w����H��f��-IH��yjd'�w��P�sxإ1[�4�H$��φ�ŧt6�)1���0�7;�`t��6Ţ�a�u�?C|
��Ϯ!��wN����&oL�_?�tbK�	�|15b��3gKm|5��o���=ޛU�"P���#��^��
|v1�r���ڿ)p[�Ո�SE@#X�W����ƣ������^eᘛ%j���+y���}-�8����={&3;��A2���u��s�?G�$o6&Vk��<�!������y�/�`��b�c�qω��C�n��<H�<�"4�e�{���]���r�[)�ҹ���6�/&�~����N����Jځ��@|���y��dZ�?��
Ͱl<��FD���Y�:_*!��^�����Y����v���[ϛL��
w���%7�w������_�~�������U0����0N(���k�HHs<b�ۘ)=�1Ѐ�q0�GDU�.M�-s��<���Nw�
oW���V1�|�/�'��b���c����AS|�QGa��~$;�lt����Y�μ�j)�qV:���$�w���`NQ�w��:M�jB�������Kz%��l�gUPHq�����P�)�� ��5�����<E��Y�9�#�wO`EQfHh�2��Z3o�j$[�T.涯� ���͒��ej�1U�K�_�ƙ<�K~��j殳I��ȭp��*>�^��n��+�ג1M#n�?�(���9�oB}y�B��i��Òd��Ie3�gHi7�ȁ�L�'z8\�ICÝ�˓�z[�nj���B,NL�$���_�����`���w	�b���8����},�a�N@ ��f���[�0�_d�S%�8*ݥ�xV([��@Gˊ��|��N���V^�AE�vm\����U�@5�ߣxN�ϧ��[�a���
�㎯?e�`�Fi�J�k������M��l�aP�D�@����[t��q�s�wA�1#�i�"ea��{�c��^���"X X�ۇIR�� ���Uۥs���U6%�e�N����n�-�oo���&�V�E�7��`�����[��B�1��^=!L���_�j�?ݿ�	��������F^B��K��{_�φӻ�o���� ��ݢeSB	�ZrL� �SA�Op˖�A�|��3(��8�֭"�L�ߕ��E�t�9��$MP}�P�aP-�|�?��fREkU��k�C���__�����<�h �J�_#���� �e O����p�Q�9�}dAt�!�<�
G���� �Ñ&�֣?�Go�zG���~bB��.�+�� d̐{W����u�9��f�r�W<U��N��1�d�E{�o�1f���Nw��λQ�֮��ꑼ�8��{9bQ=��Q��t�������IF��	��wcI�uke�$B�m7���kR{28����O2UY� ��-�iQ��H[����}�c��:�C�@�nl�+p ���f �D�@�=�,(NUPa�"ܰJHu~��t�X.^ �E?(.E\�3�.9F�fM�>��m���߮�Qm/UoY�~��Vv�:$cQx%�N�����E�}�Z}���^h�`&0I������k	^߃�0d�|Bj��`� �{������ӣ���f��I:�w�l��A�����Ụ����r7��V��&�	:s5y떭�&�=����������#6�*Ӊ�6��b˄��ВL5iB}-w/���V���}=0�!/j�;߱O�Ń~���$���ۯ�{Y�����H$|/����<rR������d�����PX�1�<R�����%F8ɘ�Q��6�m�0��P:3oW��ZU�Q��>��E'@�.)u�H�`�l��l�!���05~tu��,�®|�y��E&�Y�;��ѷ�}z_~a<Q���Z--=�Aw�P�:���@銡`�Sx����P��^+����'[����~1�`����|�d������d��� JR�����p+����W!{����	wb)Ų�;��/oD:��'�{pE?S-	{�<:����ޢ����=J����5SW�	��:���FW���Q�L��-����aD�,dj�����v�^3:�F�# I �8G�����"=rh���!^�.d!��!y;�,������x���>�z��_�X��)Fʽt�/Y/�D�U����F���J���K+�������E�#���ji[�����f%ƫ=I� E6�@>�jd(�S�s%^�V�-�}$-����n��7A���E~HbQnO6=o��T�d�q-ϵ�"*�%.��3l�qV����c�q����F}��}�*�!�5S�V�����J�۵�f�n?TlS��|j�9��A��lh�ݖ�<�w�2{��lߎ"ҡ5	y�
���*Ө�V�jWI�H�!��^��c,Vֶ5�3��6���g�����D9?=���ժ��p�K�˚�'���rQ��M�j��&|��bG�@���I���Lծ�Q�������Oo�W��S�-s����D{�}��C�#�O,���O�b>�H����~����cy%eW`�,�M֘�ء�W!�\��h̎�p,���5�	4�p%�q�Y����Y���?�J;��s�2X�/ �$��o'�QA�򌡋U3�LE�;�t(F��{mߛ�?�>i�殎Zͧ¤�JJW����נ(�e4��T
�\^z"���l$&�P�������x8~� u�[���f�EBi�ǐ$��F��j�)#�7��N3�*N�����I/ovW��:1N��W�����X��녴�e_���5�y��'�gR�c��w�y�6ш_?�oǮ�	�\'�:z�zX��Ġ�)
|Z�q�[��e�(��l�I��Vd5���KG�!ԕ�`�r���O1�\W5%���ض�xQ���hN�o�4I�02,W��ZI��?��1�e� ��4����تҸdTQ�k���#�x�.�۲�-Tr��՚7�+���Շ3�o4j��`�f���#�$��9n+�o��Y��X�'.�^��9�9�y����"OA�L�x
B�}?:��N�����{.����<�}�Y�z�}�f�T�<�cd��|�燐C�ڑ=�+��o�%߀&�;�隘��u�cI� $�h~O��T�~���h<���6��mY�5��~��-\��IN����C�E�'�p��� <Lx2�ٷ�j�2#/���ydFj�"��;�9��c�=ަ�W�Q!��M�-W�e�K�v��M���*��	H˔�M4�P��^>!�G����Ir�0�I���,$���&�9�ru�o\�	�YP�w��A����h�n��T��Q:����5���T)���)�|NC�~ʜa�f�>����C���fԇ�uI�
�Ϟ�Y����s�G�N)�Ѷ��w&���Ά��k�~,cX��]�� �f0�x �����jX�/�2V�kώ���V�JOK��R>��J~j�u�w���Gi-������Bq\V�9������("+�I�� =`gej�
@| �8�^i{S�O�̓:��\a��dga:d-��v�9�5qFC[�SdZe���!H���xc�D6��tH%��Z��T[��7��FU7v�zn��k���)�Qz�ܟ�M�n�4
��yw*b76�|o=T�b�x�dY����M��֤
��Le��Hͧ�{#����_𷆈�����s����,��Pm���5�1j�;	�kP��4Wj��,;F��Qq�^7��_~o=���B%p�y��m�}i`X���(m��8|� C[Ì�5��(Sf7�ݛGX�}-�"u-����!�F�6�	��o��!.���kHd�'�O�~Ɗ�tPd�3��|�9"�׃��џ�:e�dFe��XY�VS�����Y��l�K8�=
��f�4'�}�=G�{F�^��F;�yk���lRa�9����o䳍8=����1��E�e(ĺg�)��dX��u�����\d��#�&�;.�a(�׬NU�� I�R�:w8�^A
\B��V��7'�Z�;b��1��o��7|]O͌<]�x=�6�I,��Xԣ2��4��c7�A�5P\�~nl
��Ʊ�%�Z��^���u�N�A�^͈|'c��5�j7(��ﲱ�P�s>J♋����Xz,B�g(�\���^G8��T����ЕH,��Z��t���N ��);��P��E�T)Tk���p3��������_)��5��6�Cc�����"ȳ��;j�<k"e�pb?���=ls'{�O7��[��2d�2���<�uu�G��ć.KC���|d`{�N���^�ϵI�i�6Ǹ���k)�Sw�ul8C��h�P�,���#@��JM�=�|a×1�'~��\����က�k�p�a�c޵}b3���Q7l*iV�wo��5�[@A�ɵ�gГIq���sUo<�w��#��Īx�����h���'��l�-�Ն�\�rd͍���,�(:g�3�G"BK�B��J*XU�XU�3<������K�^``b�o/����"����HjWn�����k�Ҝſ����b�R�/����h����O�ء�u~ԟy�3*u��ɓ�$/�����W���;�D��J���!��~��ޑ�4s�I�
�������졪6YR�:b����vI_=8�xSCl|�EtoLZ���|�Lv91+�����e�3��`2t��[���9��
Ӛ��K"_$�	�&Q��������T��qg���=F��d�q�u⣿�� �Ę�u@Ԯ�]%�"k{�i���]@x�#�����'�)T��������!{z��@���<��ե�J	�}zwg�	W�e�A#l���@���cҲ��a0f(�.2��=�yOo�W���;��`m,����`�x0�H
��t12��A��M�zm!tP k>`�qwhc�@xHr��K���� ��}Rp�YטI%�g��2�4>�F�����g��/t+o	����I�[%���t��ck_���W8��ү~�^�-ݸC-��/�>��|��FO-X���`oY��� �!�t�m׏A���h��Y��uެO����w�Zz:@sd����r��vRs�a/��~�8
�>����⫤�������IxV�/q-mݝ�6ŉDm���D˴C鏴+�u�#����7���!�k����\T'S��U'pV/{l�˥�\�(.㊢��d�u�Y�tϸ���[Cg�o�uz�>5��0�
�] d<�9�oF!��ϻ����r�2�?�����v*S�-��W�mH�.fU���d�n���*Z~d&����}"�.���(�� �Hd��M�g� �S��t 7U1U5��B�����^�**Rx'��z˕Pr���^?�z���cl�9����}��������IHh�Ȕ.̞oH:��CdV��o��1�r�z^�QHy�2Q�qb��?<}���V[��Pm���W��C�A^.!9p�3�3����6Ѫ"9����O1j��ǖk�'l;�´]�ev*�\F�������X,Z�P��<y �T��1��;�o�|��?u'�h�F�?�~jm�§0Ꚕk�$q~�IT�O�*�z��-�J*'��������$\��{���um�[F��.5:���`;1U��������̣�w���<�.���\�^�=��	]<�ɝ��%?��+�'���9�2z%BBq.�u��n��W���6��.mί�A�H�����/��\��)�Ԋ)>�Ʌ=Z���6�t]����6���
6��b�891\��j��;���ﳘLlpI�oh�`����Y}C��V#6)�,]�h���i��X�<V��N��S�э��4;-��}<�9�f	����*�;˳@�ESl��>���gc��e��ɸ������3�{�U��̰c

�Ob�6���J����.�$��D�ų�JV��s�S�ҕ��g���J��x��xN^Q���J;��u	XtNH|�����1�<���u�Y$4���Ҕk}��y��<�n+�/5g+�ެ����>oqa�<�)�db��q��-,��$ľ����>M=�#(���ҿ�I�g��̑ʏ�e����'Z��ѴY��u�5�@	�b��� �������PF�
����f|/��̸�)^��H2nx\g�z��<�"����n�� �ZA��u�⓵��;���=���,��˿��+>�0(Ѵ�3���@��+t	{>�!�=N��c�n<@�E��e�TK� �0���`^(�IVD���<��an�D��*�@���j�coP��n�~�*$�9���d���"�P�IF���+/C�\��TJKMd�|����� ���aQ Ow����1�������t���3��;ijJ�uᒌ#���j��񫡩�_	�(9�i�9�sv��$Zz8�˽1>Rq+-I����l0�wSJ!�2W�:����~�c��r1�';�]�{u(�1�e�/���s��t�]�9ǈC��F	q��Md�H�L��n��Iށ1=�ݻ��sӾ�o�ፖk��҉$��ȶ(�0��P����j��|��Į$���{�gj��W� �^;�#F���6�ʘ�øC�cS�����"��7?���<\�u�wtvh}�׫�ϲZ��SL�5��(PR�����{���K��C!xҰ����f�E�,��٪�d�>WR�qئ�W�x i�5��B�����ew,T�ٍ��5שC[��]��^[ M|��t��N\������T�;�&d�T���:��<C�6	Or��q�.5��5~����K�֬�w����U�f�C4)^-1�6�MO����tڰֶ�����H����i��$���zzKR4n������r�U}9B���0���4@��N���^���|:?��xJ)�	W�ͰRL��G5�J�˾9�[�5��I�ε %�m�_�M�a��mͿZ`���	�I��V�<��@$X�_�ɵe�u!
뱏��G^�A* W��iT����pN�"��v.�t�#�_���ಉX�Or�
�S$���Ō�ʾ���si#\1q�"�-U]�w��O����:�}��.�;J�8f�>p:!�?*���6zDYĸ�-o���X�{r����bz. ^���H}�R<� �+���E���7�X$���r�'���̸�V;��J���6Y�i޷�9����L��1�����#��j����O�l8��H�����η��Ț`�!�	���+�d��GRИ�jf>�\'��5�01�B�H�s��+�������\��:';c j3ӥ��e��G���jV���a6��b}�	��S�]��
��(�� "�ęr� :��,���'� [��-v�A�CH`@!t���l���
Ɖ<_���<��)�󳄚��X�A ���)61=`gAz�̵J%���D���a_w��=n2#��W�62�&�^J0H�m�VV-�'��ͽ䳨��_tP�0�Q��:	<�!Ċ��+B8؝�(b=F,��{G��n�^zG��u��3��k'�kc0²|����x/��,릳���1C��B�B�s?�M��y�}F*x���[Hvo�8\�]��v�� 9�=��?>�p�1B6��9��"b���t=O�WK�)oI����AV�E�B]Va��̑l
|,��</�&Â��zW6����9�R@ؑah�^33Pg�#�����_�6���ϭm����	?�ի��w��u�8�5���e�X��r�8Z��^ۮ�r���󭌶�|���y�����z )��ExC�d��E<L�b+X΍0����S�>κ�B��M��^������*2l��.����I��`�ܖ���Ծ�Db�w�6�k�VH2 j��tB����qaw��� ��f��B/�����ؤ��V�_�a9L��΃�*BX9y�!��߶���|�o>�"9k�mY��՘+(���P�^�n��|�i���$jː�d�IE[���=p]'%�w�]�	ӹ����+�>$�wY�f3x|�h�z3@�)�Iω�.�@�&����[#p7X�pj��$sv�̶;�e,X���k~̪�g������Tsǥs*���;	 �[UDi�CS6�E�@
����!o���f���6���q��Np�(F��v�կ��Ha6r�RJ,��c&�鲜�_���	�2<Dj������-�x��ێ��^�ó�]�Ō�w�_�*� ��8�ߐ$t�y�4M�R�2Wt�NR�ؗ�;�D�c&�,T����w����� ����!e��
�����`J�)$P#>�`{,6���̮琌p2%�h�FbL�*�m^�u?h�Tr��0f�+�-8Q���?�b��Z}��#�?�A�@&%�H;WdbIw���j���������H7j�0�ơ�6_,�:[!S��?h�Hc��6/�q�R���3S:4��L��3B\�������T�>�*	���>t�s�w�V�XÖaH'ׄӆ��D���h�.vZ1�^!�����"/&�7�6R��C��>n�jzeAB0��{*F��|��	Y?�\� cVŝYӹ�o�L���"��oAko�/W�X���\\�B_�X�j��N6dᓇkU�&-���v�1�ǥ�f�-�X�AF����)�I��8/���Y79�F� NX����~p0�n��>�ߙṼ;���cߞ� �>z;L>N�'�cu�_"��k,�D�a��S"���z�z�L�;S��ڨn��mxr�)�ꉐ�PS�}~��k?/ğ�8�I�7���nm���}��?(���0)�s��,&`�[���������G �����0܈�an�J�C�Os��LY�10�(� �M�/+S1`��Ja^F��j`\�8�[@�=��h: M�����H��4ir�Ȕ���I����V���M�]���S�%Pԑ����<Q�şj�^���3�~H+��&d�^��/�j�!i���^`��dQ���V2�b&�7~�A�2`߲0��?����gUr��OC�e��qR�.�P�׿si��ߤԡS�N�*������RixK`y�S84vse���Y��;���&PK�x'f��q����~�Tl�÷{��JW�\.C���A0J�r,q�v���(%�	Ս+��R�0�C��ؓ��[ <��bst+WO���;����r%��BU6e��ƹ�^ed07��#C�k�H�S��{�E�Y��:��<W�o�s������D��>��sU��!(H��$x%wsd��Ej7��#��"�ޅ�U�9i�[��A��C�<K�/d��v-ԟl;�F�꥾}�3:���_h�wF����q3��������j��h���n�2q"cz�B�-奻��I\��1����fE��E�t�G��7 %MwҨX~B�VA��?��0,	e��m֞ 7��{��V�;2��}��!G�ҏ��4���`V���AO�h��Yj9�V��w�iud����\w�el�\N�/<Ǎ^Jj={��r�&VP7/�~n2�8�ଛ�uG��v
0�Q$R�[��5�Z�|og& l;J"�oC뮖�G"ZH[��	�"��0� ZaL:3p�-(�B�j,PՌ�1�e�S����Q%���\B5}w�Q�C���,;g����x3�tL��PYw9؁0�KT�~8/�.z)���`+wP��3�u�X�z��ʾ��%�K��J�8U�4�@.��� @�c�'`\ϼ}��X<<yt�~�S�U>*{��!�GS�~�x��� �E�|H����p�Ԗ$�D|wס]xl���BN�"��+���TK�D�Yey�^X�����y� NU�  %R�p��*��Q��
��L�떷F�6ϗ���+�7�B³�3�6|�}�|��`*�*(��v:�>�mN��g�jK\/o�y58�O	�9A�m���?Q��boFno��'���Nr8pk �O�:_���������l�bJ�����d�mi��,�w����w��f�=��'mH���X`1�A��E�m�{�eA毦�Zg�ySc��^���rxW�
�N�Q��bqv6݋��:E�.��Lя`Ȝ����4�s(��~�S���WE����d�vn�Z-y�H?�ӧ<ػ+�u�@I��h'~�����;d���j�n����!f�S�!�_���``�"[0�~�F/��;�l��Z���ھL�o-1e4л�U���
q���t�I�C�E?�N���F?A��j�(���@1`�}_%ڀ_���8������U��#��	�����ƃ���u��Y�ׅ���ՕF�.Fh�X�S�.ǌG�Mض]G_�Wy��{�9����PaQ�Lڿ�l׆;Zp�b֨w{�������J�[m񟰳/�ȵ���z��(A,9YW������\P��D$������	Q��v������Q#f	��EZqpW��{�ےj���9�����B8VZ	w�������93� [� h��Tv�� �-V��yUB ^�� ��j�����$��P�E�vPU��!m��^�+!��R��h(��L)*�ASЭ�?h��(]�;<�NB�b�X�m��1�؏aژ.sm���Y����#�q��.���u�:�m��2	��Yk��e�q��:3PA܋{�oﴌ��K�]ik�ɷ2�(�Vn$A��mU�}�*v��0s|���d܌�����DG�殟G���R9]�{!j��6�g"�8!�Ok3׿��k
��0���h�T2��Ѹ�=KY9fn	�5m>��^s��L����-�wwܴ�Ϊ�����N`P��������{�{D�q���b��Ma�v�+.3/�ۇ���lu�I��i��l#�j��`�Sh��tԲ��ឝ"��B���=c\a@�S���t�;w[�ܪn�x�;7%���~����v�$(먏p4y�o�i�0=��&�=�c�ގ�9��Dc�NW��X!1L�����& ~�w�cneyG������D�C�]О�J�t>�3�"�z��|�U�q��������5�:¿�]v���K���!+���7�x�x���?2R�6��3���MN�{��[j�����&u}&��1�Ҟ;m��J����'p����<�y"!*350�u�L����S��a+%kF=TO#��f��Um�52}����Un��8vAѐ=��qq�~ث���{0�	�;�փ\"oW�v��8b��vr9�H�~�Efz`����8{E"�C �<c`�N>Qf�(}(�s���F�5녻#�Fϴ���b�:��Z_-��=�#)�+��NYp��:�:qR�-S9y� W��A�N����E݈)�q��'ȥ�@�#  �
?_��0��qv jQB��VD�Ly(�y��xA*��FMՅWr���n����/'��?2�QW؛q�XW��HC�V��TU��.�ʤ����q� &(7�ќ�`�q cy��@�h��N�:n�Fk��*����Y����}fes�s³{��:�Gf6��l5K%�m��f蘦i3���}<��L�]rE/S���д�݋QJ0||I�I�/��0��) N����Z�4ߪ�I�H��l"�`��B\�ľ}��(Su\Q���ղV�+���e�]��9ÈɅ���Y�E�:��Y���|~fb&t��S,�W�J�nY�	7[�]o��B��!"|K;K��{p�'�����h��l���}f���:��'|���&�1��K���=�-i�xr`�ķ#/�����c"]�1����>G����K�_|�����1N_���43�S�QV
m�S��*y�^�e<�Y�zg�u��#)Ѭ���3���{��hx���:m�fl%���`�Wv��M,x��I)aU�Ŭ�����PSΜ�?�T��)�b5�Uf"Bal�.��sNڐ2VrC�/�צѦ\�j!CH_�R��w�#�PC�}���KyZ����#t3j$O���"��Vyzn�8�N��=�Ny���;���B"��E[�P����� 0�����f3!tT�F���"u֠-�	���
�m͞_�v:t��΃�SL�͢6�^6�Qr�a����͈��h�钟�w�t��{<*�f����/���)��OH���Xrq��G���O8@�� a'�kղ|�u��WI���l2��������9����>��Wd��{�!�����"��0���Ŧ\�)JX�i�p�ԅ��� ��V�0�����AB��2����ő�a���b�Yϙ j�z�DR2�,�b��v��-�\nEd�A��.2+��j��譍s" �Ip�8 J��J��\�	t�GV�P�梓+�������Qd��0��lУ�[?�R�ng���RK����f�W#;�XU��F����[H�?g����^���$����u,j��� Q���U�DZ�x�3�k{�Dt��oXG������x>"�����w��]Ѡ������ s��{Z0G���ٛU���%�q��Z��=jZ�P�`�׽~N��;e����*np"����vPJ�h���|���Y�Q���'bs��v��J&���K�0�Љ�ӣo��?0�����v� s|K����Rf�� ����f������hTӌwS �H��k?��&��v��O�Z��A��"���6�F
$�-u�{��/.j�;��G4�3G!~k"��0(1�"�t���ljhWiCrnւ7a��*p�0��i����p���~�=�"��ͱ2��{*���w�V�&���TGuq�`r�L���(`��qi�٫+>$�E�
��;�>�����dʪ��@;h��*rUf��7J!�ڈ�}P��z�Q���ω�F�k�@�'���/���C�|�
mJ;��E�wFhl���.���k�B�{y}s�0�����Tk\ҋ�s俪�U8��J�7���6��]-��,54�o;�o��U~@��8П���/�5�q�x���	�Q����(��x���ߩ6kn5{�K�1'�4��;�u��_�]�O~������Ep*��v������hW=��Oq�)����0^�:Q�5�����&�T�3�9�_�.��j�Y�,Á]�d�[���/z}������_��Z	�ʀ���?O0���@/��f�j���h�p���B���?D�9W��2/��������SCJf�4q�瑏�fCn�0d �&.�4���HP핎vW|���If�|';<�&�(yn�������>��U��	��ilJp�Я@E[�
cL�yg�_���P�[��s18:{%>Yf��� ��_���AET�\&�Q������9�@�G ^��}�a�&a��.t�)zL����X����8�(��5��:��t`o׶K�k�����Н}��n��Gi��դ�4_� P�����R�]�� �(�B�n�L�0�E�c-�?֎��5lu��\��*�z��$��f�k�**�P���_��\+}��磺@�ɏ��p��f�(u����K��:�T��&�[��?�J̪ګI�>z>&vn��� Gƌ��{4�	�a (�@�H\�`�|�a7 )�Y��mM90+�-����3���+*������k5<�vF����q�o>�`4�� X+P���S�i�}���i�u�4U��������}jCJd�|+j�}X�e�x��dL._�+�d��>$��p���z KFQ9�n��x+�ձ��������U� Λ-�^qUe��z�����to4:�^�)\O�G�����>F�2���jJ)Q����ߔg9���@L��7�L*O/��*72��(��B��VV�Q@� D�����K��ӕ�ǈ�Ȑ������SPY�MaH��P��DW���N)�����h4}a�֢))���P�gʰ�]�-���N�p�W��[1_�	�PA?�ze�%��+Z���_�Ԥ&!ݗ���[x��\;9[�$(օB��o��I<v�v�ћb:�$-��W��DBf�₞���9�����A����6��MݒŦD7�G϶��IvC����|-�un�?G�E���nf8̲����k����3�+�-l�&�K�s �.���O���<2�J��-'�avL3��^sU(qV�5m�K�Ƕ��G��^��K�!	��[P���K�D�q���~�Z���}y�����@>��_��00��W�|B�'��ak�l��C��^��X\x��\�ޠ�pPz1�.�ӈ'#�Ǻ��-Lm��$�u��t�g��2���	z׿&G;7�Uz�s�4ϻH��IJ��H�����P-���D{`[�BS����[d1Ud��]���;[��L��U���yc�O+�8^��1sB8
��{�:��Fm������e��c/���;�ڳ[���<u�\'Tu��,�zp/�#�j��·?6A��S1���eP������	Hj�4�m�7�_Bߩ����Ť@�K��B�1�z�D#��'�"����)9�� A��)^CT\�2�r������@t�O#����x��Em��(��ɪ	�����W��`oح�WBu̪(S Ϣ�|Pij4��+ͩ=�Ԕ�����A�+e}�ȥ��6�H?�5�PC� �W�B\p�g����±���cߩ�]�7� ��������l�T�hƧ.��T�:��ʈ,������dp���wYQ�&�S������5�"��6��68���^�f��e���Ɍ���03\�k���(�To��$%f�oq�踌d�	����a6���G
��P�MҿJ&����9��,�	|-Q��wo�J��J����y�=2 �]�3�3�3��e�,B!g���I��ϝ%�{�mJ�|$���r��n����M�ؙL7��w�品[*����{pL_tf�U,�k��Y�/RH�� Pz�'���~@�f"O�kso�<U��;A������B/���ҤnI�������#s�$�o��K��-e�p�v��T�/����x���w�D�\ۘ��	�u��HR+������uDH$��t���A{[r2&��uT�z�Zs�ݡ��t���	�?�0�z���n��K]X�P��Gx�;[N�!�'��T����\��\�ϊޒ��qT����̉��Y/ ��b�;�n.B4-q8��9P̩"ƴ��6K���Qgޏm
�B�X;@_u�1��>�,w�=)iۛ��Ib}����� S4AS�����پ���V�ܜ�ۀ��v����d 浹���^2�2��W�យ���uf�����p~Ot��-��z�k\��!�:��$$����X=_��otG���R �����@���SE8;���52��3!V=~6cz��+{��n�q^���	��)������+j'�e���s?)����h�E�j���X�|���[:\�]������J�ƀ�FB��c{�H���㗱��0"\��hӆOQ��M;��_����݅?��\���/�gE���u,��R�}�j�Q�R��0�*�����n���)c��z C�q_O�M�f�h�I�d�FB�o��(�+�Mh�I�g
�7�^2}�3���V���J�4u�ꚓ"�{��u��f��5��T�КO cdæSK�0SNE�(P] F}�jK�E,�*#��F�h�B�\���/� �V7�(���}����*^���,�9��R'������A��ʚιn��X���"C ŐUhY'wZ�>ԃҶ2�S �	`����<"��1���!���?jO7f�q"LЌƒn��������vx���m�{�����&�![����G���`�/QWG+�8�FD^�6@���x��-�<��'-� �3��A�ұz����Xy;����h:��O����Ǟ�L*�������̢D�g�G	|?��)�r��C���cK*����:i���M����%yC@d���7��9'<,{M���4���הy/���ru��״Y��"yJ�w�M�+<-��Ns4�!�})���C���"T�~T��fG����a9���ul����Z���z�:as���H6҄ȩn�o����s������a�rț�P���Qo�O4�)6B��bY������o���+eU$:3N���]��I�Y&�Nfa���.ii궠��O�����~{dЌ��oUdwp_���٭Ц�C��#R�'�J�̼za�����ϫ>E35u�KL�j�ېн�Y�l��
���Hӣ���G�,�P�ן�hv�%%�8�VQ�28z�����Ӛ�I��,zm����F�W�n���+�|C&�<X�	��立c��sy��:hO]������d�:�2�E�ˉ������ʫɃM��ps8u)nԲ�S=�nE��t<�'��n�v ����6>Sq��[訮/�ͱ�5�2�p"�{y��Q�O����ܭ�h��*@$vs�/�t�{�������W�	��Xƽ�t.)�V�~�ڌB�H��߻&��o�qKl`/ZF�ar�ҋ*�#��yb����O��&7�'$2<Qΰa�����}�����Z�̬�В4Pn����s��Q'�_��s5&��!��d�|L�����Pr$����i���c��]�,��-M�_�xX�H���`�3����Ғ�Ѫ:��%U�@p�]MP٪�>�(�ɢ�.jf�aY���@jOM7ʦ�>��u ��C��+b�N�6<�)����F�����jb�K[b����~n��师/*��0C�Z�F�7�QN���
>s�߹�G�}�]�n���H��$��$�gf�e��nq�Ù��a�4%9���������+RS����
���UI�̴h����o��5m��e�qEVB7�9��i.O�E�=������;bSÓ�y*��$�S�R�Dv	����|�Y$O�Za�0���x����w3(���N�;GH�%U�S�y��h=�{����}�C̉�W{0�3¯�/��������W��j����ʴ�ݼ����y�	�@k/� �8Rse3�j��1��q
�Yu����&�{���h	n_�I�G  �m���.�[�
):�9��I҃M%�]p	��&Q�`������.{=�2��V���5�L���_��.��V"�r�(\~(��xjO5&n 3y�`�) �љ�}ǅa�р��҄��$��XI�C��^�;M��/�N4<-��@,��C�$��W�|�ʔ��,Ad+;R�~D�u!���%q"Ф�=d�Зx ��z��i�ޙ�Ϗ��E;�F�^�&�;��%ĩt��W�y�p�LS�-UYd���^��6]�b4l�N.��jn���aD3���ҥ�1�U�x�>����8)��ʲdG}y��o�G��?��0\�8�Ű�)I_a��1��P��������i�W�(����)�]s і��F*=՗�(/��)����8?����!^b~Dr��k�1� �� ��l�G��GN!͖��.�8`��(�B��LL1nM��1~�`w5���ky;4�+�~g�屻Za�v�J����!��Ư��g���֤�C{y�c�������?�ϕ���-����Xv���W>��-V�!2�f�� �K(� ����-���n���5v< ��OX7�@�^<=|S϶�	�7����Kn����7�Cu�a̓eY\d�M�o<�L�]�b��C�U 0#�`S�=��%�����0�s��/�'��,�mP�����?�γL+�Uw�/�z����m���ެz|��R:�`˓�z�W�K��:V9��(����$�VtnxÇ����8��@�l����q!����zt��0���0��;Ek�%��Be;rd�D@^�c�d���a�4��Vulz�!dE�kx[oj����u��X2�N����%J����9'����/]_�r7��s�2,1��KJ�(ι�-�QK�Ҵx��vK��M�4�w&B�]&9d`�*g4�ul�?&���6F�"�ý}+c�%�&_0� q� j�wh����-,�LAB��m���k��]�`��%���y%H �������t���d�n��a�O�B7�1 �\DN�B�֙ܢ�h.)Z)��^/��PAs��6�l1�)���ە�
L��D-:ќ�*Kǵż��ۉ�w�k P�q⣪��C��g�׿� c���P<4��BWz-�*U
Ҙ�CQ������>�`˜�*��@�{t����/�4B����<-���`mCe�?��H��Å#�6��*�"&�D  q=N>#����xQ��%>�bđF�H����	%Sӝ�2�GtV���Y���uU�`���U�.��A$�"�|���{���j�� ns���(P�'��V�\qӋ�0���?w5���|��I��ُD���vV���h�?e�ז�~���k�	&�_ �>ba����5�ݵ(�N��9���� z�P_�B��̆��a,�Xs�6t9$U��a��^ʳb��t=��'H���xWk�&���=����P�
���_��Jiwo�Dʞ.����J���(b�@ْ0�����9f����NA�b~�jR =���,zF�@�i��/��>j�g3�)�L-�]�Pph#9Δs�¹��Ms�؂�ϨEi?���5z()�Ԡ�^���^���&~���'Zݣ]�=����h@Crl�A-��^\*MN��OT����4��V槂���8��$�b���Bj ο�Y�|�K+����{ɋX<9�8�|+Zlo�$�~��T.�D��L��֬6:��ÿ&O���,�m]���?��s1���I#��ŷs������y*i�ǒm���۽d8��mg�^X%��p�tN@��o�{��%�b�[<��ؾ���ڿ fՕ�w��]��9Y�g��>�z�D��(�|E7!���	0;�����&��Pe��*�)O���O�z��;q�;�����g�cs�u� ��QU��"�lA�r�h�a]��f���Q��NB�[����Ue���� �&�<V��fw���4L}�:䂿hm�#���w�
�	@�=T~D����4^A��r}��Ǘ��k�����O;C{t��K����Y�v!rT~o3OfH�Б&/�ϋց[�"[�F�˳!"Í��cvQ�)�����,ݝzoj&����>(|�8URP��H�&�I��������g
�y0��Ғ��lk�+O��a}�K��zn.®3"%λ�	�K��pr>��n���1�����Oغ��:w�Z}/b���
NA*ޯ�/�p�}k��04O#C�p��Q -6�-�~^�\3ECJ��Ě��߾�67���P�ي]Ϭ|�w`��n���.̒C�A�b�������piva�c�u�$V����pe���:M�{ݙ��b���fڊ�@l��,
���&;ISR�����o�%E��{�{Y���?i�?a�:������*?"1�u�����W$z��a� 8&Lvv& 0�0�g"���G�\U/V2����V�F�֖�ؘ�+"�#8ʲ,Z��(9�`�n?�`���jc��t;6�Q�^�45���(g� �հ�_-����ϘWO�s�t��KKz,G�&��IA�'f�!��%�}�,,2)��%e�x�V�g�#-��D�fNo�g�h�MCr��!�[��m/O(�؈�\�w�k'�-�R�B�G��\>��l��Q���z�̀fWO7��E\�,c{2�A��dGe��t��Â��������1N��@��DG�*ȫF��c[wv�n��[D�:!��Ui �~i�/��Pm0���~:��XL]5�G�h�'�H�$k�ß}���ڥ��]1�
���b�.n�� ��"�_�$d!3�)wJ'����1�n�+x��N�Єņ��?���)~mα�䎾�~T��� ��	 )�Sh��6����\� yO���ܓOE�G���@O�v���,P�m/���.b�$t\A�Ʒ��&~7]\+h��p?��)��ݸ稛{�J旡A.�-i.���q
�b�"���F�$� &Yy��#)Q��N�m�>��~3t��J�1+�i	�4��P��~
-dF����y|�A��(jf:����������B<�w�ڮfQ���jN�ƒ������kU
z��kX�_2��*h{0��,��	o��Ң_����K��k�{X�i�j��`а'�}�O��0Z�'Abۥ,-ac�"���Uo:��+{J�

N�
{�?�a���s٩:ؾ�U��7����J$;Ҿ���������2�f�BkP/z����O��c��1����ؾ�E���W�6D���9,����K�ag���Ֆ��)��D$���S���AL��[f
|�J��-yx��s7��d�j�̄�� 

?4x̵d�PD�����7`J�kP��<f��H��/X�=�񖒮�j�i�s���/h�A:������'���UMQd�\�]R���C�Á���őޘ��u+���!A������t��� h�
�)�r~�K�*a������0K�[ ['�Ξ�����t4��D�њ)��}$�Z�H�H��#b��D~��%߷�f��\��%X`A�7}����өu�H8[[/���ש����k�]�0U�B.Wa�c���['u���� >a�[�ƥ�/͟xB?���?�g ݜ<��b���T�ⶶ���{�͝�M?��(�D �VX[ҧ�>�q��3����yV��r��IC��4�a���7Uz��N���p�|3Ҽ�k0:6J�a/[4�/�҂\GG�@�C<�t�
��8"�P6�ʯ����J������jH��dX�mɽ��$`;�聁�J���a���!���M��:-����2�"Z��E*�HOD�V� u	?
�D?4MxB�R���o����������RC�t�	��#�T����?���������߅�<wQ1��T�d��Y��t;C�`�v&ܐ���z�b��ܯp$;R��k{���+��jRG�h<���/��V��%1�Ыe���56��V�|�f��e]� ���QQ� t���X�v�X�1F�iS�t����;�M�L"�Kr�����>*��#����h9�:0�{�,A���҂�m��;d�k�^��,�_��e��?�Ƥ�!ARa��>0�������/��Bs1/�9)6W���˳�t.�Z�v)�jRӊ0�ذz\�M�!,����C@��\&�4�
p�hd�4�����́
�Ѿ�<�6��Y��Ȟ�y�]��FT��6K��V�ߘ��
��`�H��"y�F�mu�36�f�V�>R��O'����z��u�x�?�<�mt=���7١�&��?&�<�����nI%	V�g�s5����U�ԾC�T=�H�JB�Ŋc�X�M�:���z���=h���4��@��/N�&?���7���}�7Ħ�\Ŵ�pjPp�]�
B����2�"���g��\e�E��'m���~6E�w�ֲ3dС�%à�Ƃ9���u�9�dD�	��������;�OO�>�<��_oeU��-Jm������Y�o���aF����Ot��#5\�,lǪ�����x�G3,�����7^�Υ�	�:bg�R��Y8�Z����t(��$=�2����z��O_�vء�۟A���
��ҭFm$�R̫j�sh��D?������e� 
��$pR
�o�Վ�Pm����*��/XV��m�ɏ�+�ג;�\�YZ��ӽÈr_����l+6�V��z���6��DL�=NAa����B�K�R|�,;�ޗǬ#D��/|<^mɒ��� N���s�/,���l�V�4΢���2��J��S]���-������	�Bؼ���Z�M��U�(s"�S�����B�?;����h�,��1A �,��r0inZ�FǶC��c}ٲ'�5����k;pl��*2��^�'��C@/��d�Q|�����A�%8:�i�� ���q#G��ж�vW�ؠ�����o!W .����cO ��lb�[�$�_� F���H%2���LP��A�~�����Z����n�R��"C���CP���iB|�J���1�k�l��B q����vӻ�1�z������
�y�!��E�w�;��a�Z���;�$��_���6��V���S��	��53"������~W#�v|�$V_FM�T>Q�
�gd:��Ɖ���!���c�ز�c��Ɔk�HШf����o�/�;�t��6{!;�_�Q\�-eG~M����v� �}�Cũ{MX물��OQ��|V]�	z	�tm��@�L7'D����7]�圗����Õ@��~�O�S�~h��I�}���8�g�5;��8[��"5Y�1���j�4�.k!��"ޱ�T��<-��p�����SΦ�������E㟲��jP^3'V�n3�����(&��-�`���I��D��T>�!��� �k�s��)L/Q�by���F��ϋ�+Y����[���8��?�/m6V����촦?2���������EXF>pH0�B�0�H�~qj���N�[��#4,�Y7���L= h��_�K�#2e�o?����~ط�2�������#Y34o�\A�>��=�(���G��U�T;�Ҭ>�A�wQ[���K��+��G?(,��������fb\�h�؛o�0��$vM?J®L�,Ue8��w'�n�2�PP��^V��`BǕyDɽ�p��/o���4��`!2Xr�c��8`�sgX��ܔ�P�R�M�󦇒�cX!f�g�
�H:�l6\�LE4�m�������{�����s�}��)�A� Ƿ}!�����$����̥��þ�$���/�S�q��,?W�k��G��ЮY��}C7���W�{{��ﴄs�vz�2�0N�hDƭ����-�2d�F������2�n����� L�#���\���TSuF�N���0�Ճ�)h�J/e�K�K_ܸ�`"����gg1��_4Oy�B�� Bg�(�!�5���������R�G:�"}ϋA��{�fw��r�Gڄ*�E�Wnx(闀�!�>hP�j�B��9r/=��0���9�/�;��h���n}F��A�x��૵��D��L�b�)�E�,p撍�w��e�{r��p�����N�6�g�A5pY�j(f�e1�����:���=��~�}�z�x�- <dGX�{3b�JP�bA�S�d�觧�1[��_¢�]�oz��VkOֺ� ���-�	H��O���Aw(�t��Z[��[Y[C�\j[r���^$7�{��c��;��T>��km,a�<�K�/�]z�R�ke�(57�Uk|U:5��ՉyU[��&-K�d��2W�ǔ>�L���W5҇v���O.�C�L��~vm��쬚O�Z �����y��6q�p�^�[y׮Fi�LΨ���j�A�Z���vmu��і����M�hV��-����/5��ʋ��K�ـv20���6�2�u���i��1_C2d��Iy��$U ��Cy����;�	��6J�A���n� �B����
�˼^.۾T�k+(���Q,5�=�S2��
>�#��[��h?�Ca�u1"4U��*`�����K���E>��@���U3DG����ތ5�99��K9K��x
X	�T|7\��E����+�j�`����V��mSE���%�Ģ�u��^�&=T��\��D_��.�ӈ���|�-�F��w(�j�$p�?c�S�y�j^���8��<�&�VN�?�/� D�$?\`ף�ut�6W
b�+.j�����J
d���;j�����Q�.G��8ŏ?�	D�_��s�|Ls�ia�c��akїH��.f�|���J���n�8�c�S�ﴑ��]���2Iy���� ������0O�{_OФ!t�*�� 	��3A���Z����yR­�<��9�-M�0�l�k�ZJ$�y��V�u�3{��j��8H;�	J,i#=0/lV��<�b6�z{O���~��ҋ2��{C������8S��^�5.�O�Ѝp�I��_�z��=[�?�Y#�eɱH�I0�� �{x�~}�A��S�v�_�Ӟ��<��C�~����(����� �����c�9=�y����v�Y�)���yVea��k��bO܀_�s��3U�o�v�K�]�f�GCZrf�u�+��h>���J�蛒	7��`�i�q'��K#�J!N�Ik;�IF�l�s��~�3b���e|�ZC�(#q�;٤�ɬu��}�Y.�W�-�sf��ѝ�s�|#��J��@����ˤc!W�$!�o�z�����!�4�`P�s�r�7Q�5���o;� ݟ)�4�>���	
4���oO��3X��x� �B|�J�y�!a�D�;yi�F���%R�loOa����hG�\쩸�S��	\��eg�p�s:�lq�/�;�֣�h:G)aK'�>�U�y.om��˷�g�Gʼ���"#��6��)��kI��Q�xﳈ�3�s��fL�R�t�.꒖�k:i�����)�t)��4l�I��_�Y�y�pS#]����l
E�s/qX�/­���y�QM�;o�CMy��yg�qaq{S�m�ݚ?� ˞����q�����Ά	�e]_����z�pt�		�N�б���lX�2���qR�ip��[�����+�V�w�5�� ���7A�s�|*�����]�'�F����B_Y�����b27���4�K�q>o�o�%�E��w������0���|D����a��'A�%�G�$�譺��ά�;U��{>�8z͖8��n3JY�ܩ�;��0N{/�2$;�h���y���e��Р#Y$�(�L+[6�H�A
F�IǛ���,Ͽ���&Mo���QQ�D�Blܧ��p��YU�4�~а��@���sD!/���^����s�^̜>��N��(|z�
�"�=���[�?A�z��np%v�ݬ�lL)eS���B�B��#ʀ�6*}��q�K��8k3�`�U/��f/�e��9	�籢i�w��<cß�q�g~/�s�8���W����V�v߸�=�ׂk>�C[6딬3���,�����-2����0�7��2�Lv�{��O����|�
��9����@�HF#-�v�z#��F*t�˓����Q��s�+�.qȜ�L��;���@7�&�E6���Y;#��hHrFyA�b|D�c1��iot�����3;�\E�e�׵O/�ݗE�:�N�B�q���M�]#�ה#V�|CE���M��;VvL伺����V�NEɧ�!�������pe_A=�ur-+za��`⠏x�c�0$Ƹ�����O�Y-z������W#C�qDywyX(e6���F0rO��zH�#���\\g���q�5��)�ͭ&�eL��4p�`�f�����6_$*G��Ǒ����ۘ�D1�k��ɤ+'Y�Z�������˲��D���Z�j��(�3����n�rgI����تf�T*���E(wm�~
��
(�rL���3�(!vg�%C�еSB-�N�f��8i����ܪ����'���38~m�T�K|�$����|2�
A�!��  L~�Ж�N�s:s'<(��2�jc��6�G��~:b�ʯ�8��2��7X�~��q��?I�,ᓡ�=�6��!S�I_��Pp�(�>Xzv�$d2r���!:����Cvt�Ų��6an ��OF��$.����k䧎�_��q��xm�<���14l�J��bz�f||��W��o�4J����.3Q{'�)0��{�	1���k��2\	+�3;��l��  x�����7�s9�����hi����٘�����ϔ�)���F+�Uk3�/�Y.�W���_)�΃�,���w�;z�6�\���䈅y}kp"��$w���d���`��KR�x9�*�� �����&��A�z����q��jYr�wvݑy
tJV���GT����,�|��8��rFc݅tG	6q�/��t�-]�I�����L�����F�J�h���|8�lL�H[+�&��ZF��I����eӺ0x�#ћ����eM?#$�`I����X4��n�}{~SrL45�"�� �6��ϯ�I��kf�[��\�`�Uw���D�Lr�dE&5���l�|sL��w�; ���$�o�?��Ȅo�e�˗O�|�.��ڸ��3�+�bg�C�1�I�ї��5����RƜ!?FL��8���d>����q� �$;T� Z� ��4a�iP$s,v�S>�Rx��*���a�\�݈�>K�1��c�N�2��E��{ Tku��� ���2#��:����w�;e��+E��e���M��l���#�ua��;͖>�/���nY� �~��_��T�T�#�x�Va�x���D�͈ϡ�lrTA+,��DP����@XTg�b���=���v�g���k��=�7��v�����`/��4�M�c�
`N�m�9Y�d����?u?�|�34���k���%�7K�bs����I� ������qSM�C��3_thIMå�8Gϥ����u ��d�1���ԇ��h�P�+����=�1b���lH�S���A3��f��_�؅���rU�1��N�����R^$��f
d�ZJ*�PC�_������
����Ӣ҅��#���^%�@F�i��@SSa�I����DQ�0��@c�o�F��ni$}�c �?��=��T�k��0�w�&M�$|�Wb�oh#w ���=[gfy�C U�G��V�G�b�kOUT�<i��V�vo�X���ϭ��PQ���-Z�q8��n���%���Q"����0��!��5�G��?Ǖ��v,�}W�"й�C5�:��t٘�0!��|��ZN��B���MP��u������f��y��)Or?�i�SK��T͏�����#�Y�Jn��e���R���^Qc򔬉��w���kZ~�5F��1���x����H[K��o��ׄ�dj�}�.\=���iX�o����	��1���� �y,�R����z�pӑ�+�ߎЋ�FZBE���"t5 ,zhC@G峘�mty!�)���t{	�L�Xvܿ4�~�R"܆ҳ68�-d��B����~�=y�&l�%<-�U�D�I]6������	�&�B�6Td�*,J,o����	�ˏ�Yv��W*,Rp)��y����%i+F����1�Z�����T ^�L6H���3w��w	�l�.:R�㎷�$cϣ!�U��D�K@�ǽ�/Q�j_�Y:mvc�3GKM���K����kb=�	]z$�'���'AUC'�L.�ަ(~�$��]�h>ǧ��'5��F���2|�y�GW�u4:س�4���ģ�hn�M�G%d�]¶��I*	�쎩_x�=��\�����Fci��|��E��,(_\�Zn���ځ$E@�ǝ�4��S=��0I�yLL{��^��O�oj�n	`�n�Z��~�����l^4I�9?$�ti�h��FFO���=��/��KƆ��e���?N�v��Y�%���|����V��"L��aF9����f�B���H�ac��Y��K��,��T��:Ǘ�rx6}E��S��d�.�3�B��|0Q\��rL�����i�Kz�ۏ���:�#W�E��g蔢(�0se�Vp+�T�Կ��̇����0A��"�D�"�5(�k,�&�'���/l>���vp'�+��#���װR멑�%�@X9Y��|�.����t�O"�2a^>����?A�2�P�"�xM��"�W����c�b?����k�z�Y/���W��B����VPelqj������-jhf��(�J|��@Y�����~��xE�^W�,J6`��Ɍ��by$�n�K��KA���U7٤��k�\F�|��w��\^Ϟ��b'=T�������ly�J�6���n��|��6=ҙi�ܻ�������ha��D+v"?��Hi�i�+%���l��P�JO�#3�<h޷�=��}�/tNlFp�=�Z\�?v�s:��_&;U�1���-[������u�-1�[���9�fY��<�*&ly�e�=�fmc~��_ަ��#
~�)�`"���#x��$�U
K �E�Z�@E��ʙ����+���JƋq&P�S!���%;��H��Ӛ�۠Q��ru�w����PBy�`�I�-b;	����\��E^���+i,����4�|M�ȴ�s����P�(P�S�����n,�&|}��E�S���N�5�<X�� ԫC����R�����3���K�1�3ѻP����Ȑ�����<s�2JE&�؉/�֥�t��[�o���MPp�L:��SN�L��#��D�f���1C<TQd���KԈY��e�[j�!1�O3�~�ӥ�??w��5��G�Ҝ̍�ua�Xw�<�o�\�d)�[_��:o�
�_���KTmۗ���
YN+v$�8E7�a�V����{]X�,����n��h_��6"��)�op����O%l(,\Ȩ�:�B�Uy
�<�n���;a����=���5W�%8d�
i2��)�V�����p/p�&�T5��z{R%�Թ�i�`�m3�[��D���\&�C��at;����p�NSK�<TD˾1	�i������%6-�|A~��w5���G%��jԐ�j��݁�ʝ�����tB��`	��Q#V�$��6��ś@G~ʜ6��k<�{��Ԕ��Y]C�t�qQ�<-��m`t�n�&���f��ޒ�z�[�1`�^ikVF"�^��o��[�,�KM4[F���&q�� _pY�3��F�Lh3�nyl�Y�^� �'�9�����Ňr����^��9&�%�GM��l��x�UW'Ϗ����DV���Щ�%o����T	I�^������}07�I9����(+����+;Q#A=K�M4�N�g�sR���<�hڊ�%����B���Z����
�E���G�#����(�]�&�q��`�ėc��!W��6��^N:o=� �,���ж���1�$���R�.d� =ĈO<T+��n�*3���i'��
If�qɒv��a�6�g;c���mqK��4�뢖C�奊_pt �4�A(�%T`G�O�D�sL��M�M�laT�3�\�V��4Mt	5' p宜τ�e�H����-#w~��4��Z�՚!�dK��2t�VD{cP�C��������U�����C����ꌈӛnFdTr��zH�O��ԗ�$w���.oz�n
$�w������H����kl�IL�b8���B�".�P	��Kb&�8~a��9G1K����TR������7J �%EW2ws�$O!J�*p� �x�}LWp'S;�3��Nf��rU=�8c�!],��0ϖn��BT^���><��
���N-�zEz���/�#.f(��0��w?�;Zv��$�ݚ%;�4��t�g�p"���W�:>n�7G)���jI��{U�$��=���7I0d�/󎸧u1MTnF�n{Ǿ��|����Wm�ڇ��J���C�T��-8�$z��@� >��y�eu��V��{���
w�	6L��+d]T>x��Y�T�g�X&�t΂��y٥R/�Eu�D��~���!��k���ڇ*j���]�>�����ֺ��I�0͓�W`��uD��̓�D�*�/�H$�`��D�}��b�N`Jb�������H����)45��Y0�.�[wi��`�_��e}t�[͕mZT�����F��LY�_�<��|�\�� �(h$��asp�\L����X��������X	���4�G���S\�-�(���t�H��&�)"A���Ċ���%48�������O�e��9�� �iGZM=������Ѐ�K�L�=^���1����X��UgG���!nMqYAD@���OףGF��P �A����q�������SR�,k��[���ҩ��Z{���M��gP���������li���֩���R4��o�P���w�(`S^:�JtQ)vCI�K;�����T8q���|���Ux�u� �y���[,�˿'?aQ��P�Ӝc��o�'.G x�����	NA����os*�v��GǗ�wdT����� v!��Z�Ya�B��m�c�Ե���w*���t'�v��8`�jL���:�-(b��R)��j��gC������Ÿw��!/E��\��D�tG��E�7%A�~�w�����q�|���_E}I�`IQ�Ux��\�W�l_�\��`�ʔP����!en�K7��e�
��\���_��j��%�����L���[��&����8�<l�͝��_]Z��w;-�7����s?��8\�N�(
u�]ID*�LCn�<���~�[���+H"8�� ��#u�L�2����uA��U-PT2 ��s�Iǿg.��l�X��9GLqN�v��)�܃f�i���P�oG���:Wԡ۾�ފ��]`n�]�;�A�����6�$b�e�C��c�S$u��=6!|���h*���lN�����&�Z�O�Z�.pDƯj�����BP����V����њ�=ع�z�|i���ޡ�E'��L&�~5/&�;e}:�*(t�!&��M���2{���;W\#��=W�q���u���$W����b��Wy�tǱ�p]t��L2�O9�/B�R�:�{W����qi�BB;��l�%\�����^��~���?���s
��-�s3]�("�u"��t������JH�w��R�~�%W�uwR�g9#{gĺ��hP5?�0W���d�7D�M1kX��8�4l�O �$5V�~�F9� �u���	L?���lu��C�8Ʒ�͑�8,�*ɽ���O��$�]#������0��?���bx�+<��ƒ�5��'x��sA'n���Zhn�J�V��Vw�1E"�,g!��-�,�v+��΃�B�>:0qKƨ�U�o͓�j�w��Я%�;d��B��d�b��Z�9le��[-���z�~ ��h�7���Y~�s�l�J�ĕ�S�I�{{ RlR���)�>$��R����t"	�Bv�[-�>��P�UŖ_L���ZB���l�渆x��;t��}(S��x��\��E��$����R��T������*�$�#��f���M��g#����Q�eqnsH��L߻B�k��k�%h�e'G���jJ7��6�RG��K̈��`|�G�ҿ;��	(T�=?F�'¶V�h�Ӧ��j\������+��	Ϧj�(��H���N�UTT����:h�z�!jN����B���h;$O�"��r�l�k���Uw�y�αxκ�B�LP*F��*y��yg�l�ʯ�й������7���D�e�mv�yM]�����@߾-��)m��8�� YAj�6a9C�_�l�J����o� �O浑�_ڗ��#�T�w/����^G"�eP�RQ��,�_9�7/�>>�0ve=��h@����N��?n�Z֖]�	�S�r(�4o��\��/�4��tז�3O+�S5�T��m4>��9v��w����1�hG��I��ca֞�UĨ���ؑ�W�^Y|2 ���홾��qy����#�iC��� Ⅾ��u%NZ�D��3�l���8]5��?ȣ�~XN0�9	���$��[3_��s�|iOX�VG����ө ;�K�Jkqa�������'�e||�9������XR��#+�w����a�l;�a	H��Aq��BL	,L�"�&[G�P��J[ޑY�:~��#෽�"�>�Wf������HCI���dC=���V|�8�!S�Mb���*��!�{�������c�*��@."<�+Ls-���Y���c����ׄ��D�{ɏ`Ӧ�bv��1��谤 ���ߛutWf�P�{6!s�1�Գ�Wч�>b΂�����%V,�c�3]����x9��������USC[cd���	H�	2��2�ulI�bl%�8ć��wW�t<�_�:���~��֥�8��\��h�?�:XY;[43O,Q� �i`��,9��ᰒz/��3�1 ��I\�J���on=�̝$ƔZ$Ѯ�z	%;S�W"�\��|�_�������T�ѣ���l)[���V�Q���K��,^�֚K̂�&v�z�#j�$��Id��~�x�c���c��1'�dM��p[|Dn�*X��p�z/tM��؍������xJ�tz�Xt�O!4�B3c���>��D�ej�R�["��0x��(��%�yl��=-Y�1������92` �ܑ�u�z$}��<K����ۘ��`�D��D��/�R,����L�!�5ݺ7|5�k�а�'��,��1�����1mo�����Ƣ9�N���;��/����K��i\��'1����l����WWT�����q c,�ވ���Q��pfi�v����X�R*;��li��®l�~Ъ���U$��5���u'��U��a��ά!��}�y���n�������H��U��U>c��"��:T���W=�nG5�)��+�^����Z��k}��4f���8�=�S0V��u�4��`JSuK��D#��?�vB�a?��cô��<�:m�G��S�g�LO�9Qa��_U;fo�-�����~��6����
5[���(�xO�=��ld���B6��z��2 �'m��q�;���20�j�V��d�1`T�p}�Z;!�<���� fo��t?�дH�{�Hhq�����F�X����"ea9�*�6�gʒu�)�ֈ�-�R�����^~�Lc��I���cuI_�/�PyT�1g�N���X��Fu��{��;Z�`�9bX��<�:��߫Dbt���x����i�^�}�8��3� ׹kq�FS���8�"�c������"y�����ٛwW��!�������:�%�LT�q���N>W�ոm�*�Ahݻ�v�]VKG��1DG�p^X�Tu2�Ա����7�>:�>�aG���r���v=��L{z�(ޟ:_AB����R�x���҆Ȍ�[���O!%�]Fڝ|tDS&��)�!T.?��X�y����l����I�x�|z��|UQ�l��!q������Ŗ��6����<�@[\A&��U�tSs��k+[��~1�mK�ڪ�w�X�T�S�f�p�,�{����������s��m�W�+���;�Pv2R���!k�X@&��6��K�E��+
���/��I<c�s����dsށ���0�nfb���yanR�22R��<��\���j�ع�c��96��a�s9c��`�_��*��ͣ�,�\ 6Țf��Kvmŋ���"��Eȟ5�a�>Yd�&TS�T�������g����Ə4�Z���e
�J��E]�s�����Tk���;|Ph:�n0b��2=��w �(��L��`���h��&a��n�����Uub������j�x��@\}���ܖ���ύ�~�����nڥ1��tf9&����!0�%�9T�����qx��Vk�?ژ���d��9�v�v������-7�-b$����� -�����-��>����r���P�tӚ'���(�t�?��V̺�r��/X(�.W7��v��9!,o��R/X%(kZXݹ���
}�ߗ��_7�.�`!'�N��z5f��aT?���S{C@@�['2U"���f��h���}�+f�#�=�d|zƥC��1ؖ	���.u��R���v�DN.7�%��e���įd��?��m�C�>V���ܪ�79P I���!,^i�~�I�_AX�ƺ��q�Hhz�b����3�!8�鶏�	�sd/���%U�E<��_s������ʓ���؇��OX4�p|K)� X����7��a��H�07�!�	\i�Z+�< i��y8Gր% H�_b!�*>(��*���|E����Ї�Hn�]
�JMx8�>�p~��Fv�d�a[.���W���oN�#���`x/��n��6~!v3@%<�BMy�/k����ᠮr4l��f�x��b/�e�e=��O���L��o6� /��]���i��g"F�������z�LeI?��nf�߶!�.ެ].����TX�r�d����w��P㜍_��w���B�z�L�cv/�t���;A�K5��+A�QO�T�Ҥ2�b�	�GD� T�p��������)՛���s8�˃0�-m;M��#�3�@aX��D"V�Η�ET`:�r�E$؎E�┌���Ii�o/��:�5����Ҽ��^��n�~��H��Q �h��ڦ`'Z~׼�Gb(7-\�f��H��a~�Aֳ���1~�ZLH�b��o���
�γo3�(8�����L��d����p�%6���i�(�� :�N���������������
2��#�+ҫ�j�S�/�RB�}��x��'��L�n.7S>��
e�L��A���4��a�DÒ��'�G'�Y��������-%�^ө�U8!��7�g�;R���#�p�*BI�sIӴE���*�ќ��?	�8U,XE�¿Hxݘ7�&�W��dC&�$�Mk;�_�q~Y�._�K�Qj�hƥ:C���u"l��
�cnF��0�/K�@���ۇ�:�F�Hp��9��Y���Qd�
G���JON�)i��D��b�v�Ţ)�q��w$�um~�W�~���鶈����㶦o���5�C�͇�m�e��!���7���|��z�4K��ׯ��!��N8����%C��N�凍��Y�PE��a\	Nk؛���OOp �44��QI*=�mظ��J8f ��fI?�e�TL�����}l���\ے�H\�� ���pHo�X�'� w &r@�5,�Q.7����k���u�
3լ���L'
�?4�&��ݏ�@d����@�Ʃb��L	SsD��J�]��k�u�MF.+��?W ��k��Fһ{��I-��i�E�{��ȥ�q:����-�A�#�"��s����T��_���YJ�Ƴ�V�&�w��cn��S��?_��?@q��n?�k`0�+��St,�������"2dq�w��;v�]����#7�@��l�Ue��J��ٮ�^+I���d"���i/����ʰQa\�#�uB�f��Oj���P�Bl�<������n7�g)e���Ґ�4fO�k/��SRvˏ��u�T簇� }U��ۅ;�񴲦O�o���_g
�Q���#�#�/�	կak��e��k����s�����Nڝ���9]���K�XR�0�`a�8��攃o���B�/��lFc�֖5�q� �SI׏{�*��갷1$�L��7��r���B���v>��8�(�d?=(L�>%UhF�K���$9��̽M�����l���r�+�$��#]�(5�����J��׸�ڷ��?�>?֑�rd����O\X�$F2��p�k6�z>YZ���+�,��S���'`�D��o :<��7v�C���)m����)�����k��py�vF}U��^(�8���;LK���DB&'v��X1܃Ir>��´���	o#ȇ�Caqj�H����OܑJT�k��.z�+H����T�'3g흚s�=J��pG/�W��`=��q�݇ۧOg#�g��fk�P����ȭw��"�]E_?�c?����{�,�t�|���yKX�$�| 
�t+�%�M�>��f���� �_���T��<���*JA�f��¶f7���Î���� ���N��\c*���+b�`�)�L���ew�)hTޢ<5�}8E�Y��{i|E�w���P{6�n	��}��bJ_#��0 ����E�y	|;��&b���� �!���k7�K��/i��R�(Rp8��y�hq%�ȣ~L�oلD�ow&��N��B�_�����Pa���J���ʊu�x�0��t6Xn�� ��� �㧲dy��@�c��[�w�:�
�/�����/�|ZzC��vv#R&q�r�@Ƴ��t�$0#!��nq<��u�:M�ں��X�z˅��u�3��� ��[q�PY��^ׁsl�+g��Y�O�S-R6��6�f�E���:zbZn�A��|<�g�Vb� x����lm���×����F���#�_��X ���>����3��_ꍘ�@�����!����jsz-�����:�)0e������5���a�C��&�k�_��ǲ3�.�A%��@|�����UR��_EJ��``�`�9/ntŦ�ľǕ��Q+֙J<�b�"n�뗻���h���6�����ֽ�%F��]y%�Ԯ�<�w��E&������֎G������ߣJ���|�nR�Ӽ5�K�M
� r넮����П96���``E��L�L)��i:��ҫ���)VL�Ɠns���a�SN?�h�Y��N�����·+�i1�SE�<�*Y3�ϳ���㕟��s(���Y~�܎�,��~��l�hO����=��[Og{{�S|�T^p"����K��\IX"������8�X4���<K�!J_q@D#���Q���>��:-�һ��J����:�4�����}����A���	I0ִW#��ƲUz��܁�ޓ9�m
'�p�f��`Iv.�{1^���m���5�d)M�� �P�~R�	y��1K���.����-��ݛ0�>L��U��h)`��U���7,�M����&�%1Ϟ�,Aq��c�Y뢰=��K�i��=,�7��H����w�A���m�|FS�Ju����|[�s�D1��<�7�K�n�@iP�&JOy��]��8c��, ��)1�*�L��K�H1��hA�6�Y@j����h������vx�P�W���9gwʵ�y��y��	��=[�M�m��w���;��jf_��e���z�`��eٚt8�E�=�<���8�|������S�� W��`�R�ҥ�a���1^W����(�0����6��mY�Z���%srM�� �9���@�ҮhB��,:e���ٱN�܂C��T����y��Y8�aI����� t�JWe��{�3�r��[3�C�Y�g��x�G���� gMd7*"��»|rj��.�\�ϴL[��|5������,\������Jc���ܽ��%ʉ{,?{A$�h�����j����?�x�_J���0�s�$��`�n&u@E㴨G"�}�bQ��l�]!4$J� �8��^�Ws}���}��{z�%��Mc�Ig���k�:���$�z�$\�j���4�~@����	a>��F��4ƪl�k߮�.,�hŜm�re}K�.��B����V�s�wȹ.� ��D6��u��}R~@��G�K�GZ��g�0�Q���X*��$���\�=�WҶd�0V,�4�gL��
�U�y���L;N�HI��X�}�[S�b:g7��g�B�υ/����4 G$_�,<�z1�(��d_����� ���b�
���'�ef	k�/V���̌t`e��k��l��S7^RX��W�F�%�We1��Ȯ���_�����;J�%I�F���ݱ�� V.JYDYC��}Z��۪��i쥑��x�(��E��І�#[c5�G�Ɇ� S�;,�w<q�}f�DРm�}���3����KȻ�M�w�ȴ7l�Õן�Ӟ�s�볍k��?��+vI��6�o"��v�|�풞��H��?
-O�t1-�,����h��"�IR�a�ࢂS[��}���x�`F��UB���@���#Խ�1ui�=A�]��;����e�w'���^7yE�ߗ��4���<��=>�%���|�5���Ǵ�*�2@*¢��p>H^��+�h��3A0k���371m�k& ��$��yW>�`��
�TnD���	�㛺zPwYP�'�HnC�F|?@�ئ]�+|����I�-��B�W���J���TA�+s�=�4�9��<3W�~�6H�/�,�����:������>^C���q��1��	7���׸��fJ�����>����q�����Ү�vv^ ��uB9F_���+>���ZE��T���^%\��(��WLZ�6���!l�SN
ˈy����*���}.<�����mRGy�"���������)U|޷^�ْ�m�l:�L������'��q:bPK���t�
�?E3v'�&���$�L:��ǆ���|�6�
mc����Ǚ�,n���͞-z�:�
�����7Q�=�nc��T6����OO�ԌǨ�8���\�N�M�<�틩g�;��ލ�NA`y�'�B���:����d`�!�[��X�y��1~i�7R�إ(�lj��L1\� 1S+{��֒ʜdJx!p���G� &W��Z�S��0�&�+�q��o2m6H��H��Sk��[�݄��N�5F�i64���<�B�g*^O@K�_$��:�^��;��4�E|HHiq�c����F��h�d�dn��i��2�� rV��9�q��1���w�7�Ք�C�d"&fq*8 �˧��`N�qѧ��"QO�>)hB6��djD%��̓�e'�b��u�p�U�U�4T�7�I���5�z 2�8k����wxᰵ���q
�SU�8�Ws�1����#�x�B3* �@	��� �y�a�=vtX�uJ�	2��?m������	��o|��,z��\q�ɼ`>��c*�0��8�8��r���9�7�h�Ke�o�� - ��p/�p�r�X%�/E-���U޺;����g`�[���NMk�ي���S$�����j� &��(`��W0&([4^�I��~q���'�H؋IT����9��e'�E?΃��}��"���ji|��܌4���nw�������`ofY�ű[�ˈ-�A�B��8=��O�!����KU�6R%����֗�Uc	p��BEl2�9��	����?��w�$'wߔF�_�0K�Jޟ�R����f���86�+��Q���~�N�8|5��νXq�Rz)�-�%i�+�Z�E]��70���N��J����@�u���L�\�XN�럄Nغ�Z��5��K՜N�.p����r�w���ԓ�|�p���H�\��zr<�,!P�:�T��=|U�k�]�v�U���5c��e'FDE
��[C7�ƪ��^�]�#Q�B\@D)�Kz]-P�����	I�?m<����D#�[�F�s�����TjH����.E�����W�۰f�=���µ[�pK������Tx»�p;���A^,w�v �G�����~jE�����E`�Z ͏#�(�(�RܿޮQ�P�:�T������X&{����}��?T	���ຏ��w��t�~?�.`@��3��F���W��͹﯐���ɾs��'�7P�6�Gf�u�˄�e�d��Sq	�װp���I����j�Z��`j2��?�M���d�§���1Kb8|�x�oC���M��)뻡���fdAپ�g۱�+�
���Szg��_=t��% �U�V���bNJ6�E�"%3|XA86�j	9�S�;�R���\I�,@�D���3�NT<���6���9::�2;#K6�l��QL@��M�h7�cm�E�T�s�U� ��8��Y���`���q4q�vz�����kʸ���mp��QI6W[B&	�h��vh����
0�}�e;��FԖ�.$'�7���[�]UΓ�L>h)g�6�Y,D����=�	��'!�Gx_e/��ҳ�}�|x�E�-�U���[����x�-�e�x}1Gg��_�:����XL���M[|�
WPZ�"�nȵ:�<�#���c����^�V��kRJY�6��`"����=�|��{7=���%&[R=�%ٕ��''�4BDb�8�3>�o�N���)���u	��|���:���h���-��lE�9����(>Dj��&J,{k�
��$h�˘�Js�\؜�m޲lAG�Q�H+: K�l��t�z?��^A�'B�A�k��v@�����y؎�1	M%G�d}&e�b`��I�J���W8�n�uz�5n��b*�Cuu�炲U�2�]�h����������"�Ck1�_��T������(�6N�/[w��y�U ү�
"ܞ�C�-��Yλ_p
�U0��EW��T]PQw(6�D��.�!���I������t([����s\�o#�GU�f�f��)hN+K&VPE�h�E�J25�"�q��L���:t�X��Cr/!"p���ҩ���~V��%�f��<ta����q��Bi2������'��)C����f� e�#��)���r�\�w�zu���Q�������Qzɷ{8X9!�B�]ϸ5�e^]h89�R�u��!������~��Hw���(��l�����0g����+OF�>�I�'���P���1�gG�'�J�.xVY	���[EvzjA��q�)��������ri��
1t�?��\�a�zrs�'��}�5)�̉�����I؏�>��ڈ�x� ��>�����(�XdA�I�[��)0Z~l��hUtO�d�g8�Cat�	
���j�
<�cj�EJ$�����ȓaLs�Nh�>l� O�7%^���
��P���k�~���h�b��S��iCR�ڤ��~�}H�SQ������`,�&q�\p9Z�@����X#�C93+n-�
e/��Rs~��c�`�XY�«�햙�8U�����Q�\y�>�Ct�^��?�i�X�Rꍕ7!�^|xA'�Q�NRͅ�7�k���;C�?q��m�eH�n�@�������3J8Q���.0��F� I=�,@3O�qj�r��7̵I3fU�Y�i%�[���k)�A�[14�,�=��.�հ�������(S�Y���W8�m�Msæ�H�d9O
��vb�i:����vh�o�T�]#":�aJ�.��{�4�a7:	��i�OŔ�nT��-`R���R^�<?��L��C��K����?�ø�#1����)�&�K���u�s� l�#K� ���uM9m�琟}�q�S o���M���hA>���.'��ۚ#kh*kiy{�G��J�M��\Ї�������-Q���	��	7�4���#9(1���]Q���D�K:��,��a+�X�-�c���w�&��$���z�۠��+�.�c�n�����	ԯ�Ĝ݂*(�n9C�[�s��l���.�>�WqV��?�Q.�wi�v�G ����(Hɖ<_�;7�%�W}��:�*b���1֒�Q��i,|u} ޖ��0�Y
$p}r�H�?g��uNdI�:	m�"�pϙ�eF�C����*^,����d�¯���/R�6k��}����{X�Q�R��W^�Qvt� |�&���Z
�c�n]��7x�P�
J
�}�����	�(�$���:hS�$K��Wy�N���2#=Poj�.�ݭ��`���{�i�Bq�'MQyS*�� ~Rd'9�=��E
ּeyث���aF+��$
#J�ؤi�DW3�����>�b5�������J&V<��E|_���Ծ.��d�y�������׮���_>-��3��rf�pq�HZ��4��̸�3�A/Q�Y�!j�A�D͐���3d���k�glH`Rp��6Ԗ����	����0��6���e��GY����� �l?X�����R�Ra��ߓ?}H�q^�/��*��/u��/,�O�!��q�^�����zV��ف)�~@t� K׏҆֩r �ɉ�j~m5�1���N<�Tth%�	;	���ԥ-[�	ۛ� �W��9ƨ���?�@_v��K�Y.�G�P�}˥{���/ ��AI���v�*��{K�G�<�����Ia25��%1C2�g̮�}F���)l��7�L6���a�뀍��?o�C��_Ć���D�E�2T;��2d���:�s���N�X�ő1Y�:Y��n�Y�o�9=�z�l������δ��nh��K_F��r5i���<$��At�f���U �&B�UM�rW���7/�����`�@_�;�@�0�4)SЉ�\��qp�0�oZ��ǣ�b��V�
Ӥ�γ������|ߟ�������h��	~�o�w!q�~YNX���m������'ޙ�y��=�{8�/X��:��)M�b¶9����Ѵ��TG��·b�QW�f��(<6�Ş��RD���آdIDVG����/�1�ye�0�5��c`�K�c|�ɢ�U�a�o9�������ϙj+�һ�s���H+��x�b���<p̰N�=���?��ER�������t��i'&u�h^���,}���Ht���!����֋|Y��?S���LM6��}�&�&��n��t�qt]�����`��{NOwP:�M�������|Ϟ��p28�����dOָ���C�v/��d���v������s���;�bJ�A+�����S�H��LH¯'H�y�1����`�E�4����-1�)4�x�S���y�Y�<��[̆8@���|���s�0ӄr�B2�+e7χ�ht�$�f�07�^�e\�"��&	9:S綪w��ܪk��0�i�d_G@$�|���۩��0�u��@�������O ��~�ʐ��]������:I��K=���£��p��(�t�}Z������>�K�����,�Z}B"j���ԓ�J�yŲ8ɩ���h��B���*�U)���+��B/�E��(?�~�]t�]㯔	�l�z0( 4���xG��4#&�CF����³&.;�T`9/����@��9��߷�\�b�T��� d̏ W�Y��l�\�N9�8Rc��d�5�2�����sF�����mg}��u�ּb[�K�Py�~M�WcH��\j����I6����d,�?��\�����~pf���<����Ӟ*P�K+T�h�MU2-S+��I:�s��V���N,���F�œ�jχV��b�b?'U�S��'���+�S�e���լ���U��F|�9�%>���z��M���e�)�4Q��(�P�;�@����;���}`�9��*��u���K���/���/�ږW�ڰ2�N�<9��X>ۛ�w�Lu��a:n�����$���<}�V���\�<"̽l�<�\&t��:���T\�g9(ޝ7	m�CXnߢ�La8�gK����{=m�80"��)g�dQ�����@�M��3a��&�>�b��.��(�{~4�Bⵚ��W��w'M�V�[���-�6�������TO�B��� d�V����A!��C�l��ց�a�ba�ۻ*A�轜0�3�?5���U����g�u��I]}������̃U���[oz�$d��n�xH�ۄF�e3y��[�S������{yo;TkE��k{����ԕ1�Z�����"�Z�H�:Z���m[D*��m(��R;rʹ'zv���V[B����{#��b�-o$�ʉ�Y(��!d��X#
c"��[Wi54h���D��*�)�׉$�,����?�Yw��q�TLQM�K`s)G���+ڭҝ�wY���&��
��i�m(7�Z�L�6�.SVL �����7ݬ��S$	�RէNZ|v�d_���
�_���k��Y��l�#�V^A�4��C��R�Ls4Kw��s0��L	.`�-xBD����y&�y�^�3�7^bG�'oe�\���;��М坅�`�];b~t��
�u�"��,���;g�Q�y����q�qW��1��_��Xj��u��0ǣҰ�y,� *�as�'��|K��H��?e�6d��Cl�� �e�������Y��'ۇ�4�2��D�xّط���?ʺ���RV2߂o)K�c6�]�����F��<��x���}	��=�F��EY����9͎fe�9bѿ�|�٤��~����n�Wج�iE��RF�T[��[S^;,��S������䢡s|��bT<���� �g)�AV�)dW�� L٤q�?x�����mEHEP�I�p �b�>x����81n��Lyv'��ZD���W��4L�-�0���ӣLl���	E�W���(>,3q�t����(�2�QjO�?��1�s2��8�{GzKR1�v̷P/k���"��L�4��,��-�F�ص�ڔRg�/hCݼ�}�1�g��T�Zt�xq�6��)\���A�m�����3n8[�-�n�̢u���~Oӗ��m&+w�D�M.�f��T���u#8���*#
��!,�^S�#���D���Ц��D�E,2�ںV-L�^���.�}��FOնہ`c����;�r��PWD�4)��n��n�ܗ�[��(�k"�Tc���C���ۼ���B�u�ˏ9,ZTgdNlZ��/��kP�
,�A�h������>�Á���s�<�H���=@��0c:iu]I�� �A���6�%��c����^�^[��������m3�/#�ԭ���\�:ZmB1�֠��ɗ��:,vl���qU4�_�;ir��<��d�x$��sШ�fh9�H�x#��[�� ��X]��8���;�&�i� �]�=
��R�OI�=(�2a��@ E'��	���N�,���\��b�HQJ&GW�Sgl����4e� ��y
kճ�	R��)��L���\體kV����ڕ�����C�\�<�����8q ������M���WW�96R��5�)�Z�����{�4�'~���z�)��4���ib Jߏ�pu��	�ARR���bWj�Kn-�$���2�NY#	Q���]�S��us����OևIFב*{�em��:�pϟlAH�����������@)��jR���(�X�uL�w�BР7�������w�I�P�嫶B��J��!�`w{/Uk����T6�&Α��7(i�1�d!����X�rO_nT�BOu���8��o���y�.������B
��ıp�9������^yBhߍ|,Gx�V�ќ�͐��5��F��9������(�Zv΍MB�|H��K�Bg�����T�چ:O���sH"����r�!+I~n�*�X�6��%�(&va�&��D�{�i[�X�qSΣFl2�hq�g 5�Zw눱H�5>l|�9Ő7r/��W�m�n�~���'�u����:�sN�'?�E*���[f+�i7�D��:�_h�:!Hl]�t�$s�j]��%~N{ I�;�R=���MН�k>�`!!$�=bng��PY��1�7?�*�ڏ�a&=��G'�b���#/�n*��K�N :��l0�!��������������l?����l.h�/ʭ�T~X�,&�t<c�Sׄ]n9V�R�D�4��'���{��N�[�T��p�H�b
fȉ�n�)G�@YUؓ\���8��`��pb��]D
��}��ɺ��o��4�|¨ǬV��d�&i�3h���f9����U���{Ԙ|L�T��Qܝ��2:�B��)��;*WS�8ѓ5�u6�uR�=$�:�SAvPŲ���@o<�Uڊc�9�ZK�����!z}p~�a�x�e�NV���t��3ӷ���_�~cg����H����1���t�?�(mL�#�8��rET��F�A��}Ix�п��ڽ�l�#�d����T��xf@g ��޴5����Y�P$/I4�p9��lJ?z�q\WR	�}��d���vL����=���ʟ�Ӵ���"G�UGZ��)����Ȓ���J���)�j	՟\3�\0�c�f�Q0�e���x���慛t�d��\�K%|����}�-]����;���)�W4E��u�'�e�b��$�o�2$���'�;��r�#� ��wP�����Y��.a[��H�~ u^Ý����ޒ�����^�T�fܸ��Oā�K*���j�!�F�V<n��|��O}j����ȼ�.���m,�ڈ��ēܚBחZ��\ZSa3)�ݡ�#��}Ut����PE��:"�j��^^�G�M�P�#n{@��lhU:�7E�1���0��%b᝞��~�/^*3j3��;��v�@<���Н�O���_�m/���HCbN�u�"�<L�&�% �$�_m�d<����e��M8�hD2��� 2��[F�<��������ڛ��D!����fSEѥ{\t�5])}9�����!����ǋ��&O�f�DO͌�)��f8+�[���X][��:-��w� ܠ2@.�lW$M�������U
�u��(zӝ��t�.��7���}Gu~f( z�)�j�񫩔�L0��L��cǋ�t�6й-�z���$�>0���(�̡4G6l$���P�����e�i��M�&�-V[�`ώ!�V���|2�Ұ����#���dz*.:��А}겏�+�.�;�:�d��:`{��u�M�&Ŝ>E\9�)�^ғ�0c6����Hpަ�&2n��g�99w��7�	�����4�.Wq�ps�sޱ9�$�W��qc^Dc V聲3E�g�Y�	vs,$���S�pSl����/�{G��x$]V� t}Df�����F58yz������
!8�	(����/p+z	�E1w��j_A![�ɡ�������c)g�����WL��1�T	bu������8�-d����n��8��?���!Ɔ�Q��g�?�c�:���L��}��ʳ[Պ]������"�r�W�z(*0�	�SF��d�ݞʇ.lܿ���M������L��Z�d�+6�����G�K�q>E�Gm�ѵk5,��zD�C_�짞ٴw׺�)a�֞�D����J��pEɝ����S�j��M�t����wb�ڂ�����;vN`�dCǰ�������Vu��-�nS�P"k�K8��j�CTw��woJ�T��u5�)�4��hu( �TK�4r�p_T%`�Oa�t1���M�RN�7Nu0L�Vo.(l�ٰ o��1%c�U -e�L��>$�W(�����!׊�V2�!X7��u=���Y�O�1������\ݾң~iT��ιK}��2�	7U�
��7�?X!���������\E����Z��Jlm8ދ�m}����2��M��[l��� ��u9�;�\����X/#��`2�am��9)�sQ���8o�8�t#�l��zY�E)�&o6���L����)�)�@B��r�]!?Z�����ݝ���
[��ǔu���i���݁�����j2TҠ�!�E�qz���sp����Y���W�k|�i��2N>4�C��P�vx���\���"��N���#:}&�Z~b�`΃�}���U�	�f<2�G�!�j�.�o&�% ��o?�0���Vir"&qW�������9������ z�U�=�3���MԪ�����z7Ez~.�b�S����b�Ti��O��P��\ 3��$�5Imb'��KX /�Bjc�G\�r~�&k<����x��S�if�!Y�\�m���	k�c.����fcE�V���D�|���� !~�-e!1ƴoA�I�C��T5XC�ǆƄ�
��9Q�ܨ�[����@v@xX6��V���{A`
�*����0��z�v�[M�
{�R�k����;��>��n�.��?��^�b�'39�� �
���U�ֽ1�h�w�q�]��>{\8Mk=w/4�p2)AU��)
m×z9E�@1){�Lp�����$.�Z���R(�!r�����hx�לu��fJ��m�𧊗�d1�	}V+p\g�2/��ދ`����ŝ��Z܀��X�ya�~.<�$`~�L� �Y�Ie����I7�8A�G}=*�ڰJ)�X rseO���c���$E��M~�J��i�y=�{�;�vi0��M��C�$-��1�B����ֳ��F �-��s�p��G�)W��Y_�y���{5�*��Ⱦ��[�h2\�7�Z-�	�[IU݃�v\��PL?����Vi`w��p^�5݉L��Zu��}���~�0�v�!p�Tgj�6�dLQb�S@��Z�"?]_\)\_/�����ȥMwP=��8�U��D1��'�.i>�s;��',�~��1}�Fj�/�)g�4�ʆ���W����Ѯ&)c�ߏI̶�ޯ�M���C)R���o*HYD+x�ɛlL�����M/� Q�U��χ��^<�}��#^s8�W	�*��U8�|�[O�y!�֒�������,�5@���KEk�eZETy�xp�Q�w/�Z�%"�^�)���PoX����DM/�A"鞪���s}���2y^�M�ֽ�%N�p)ܯ?�XZ�������Lg-w�V@���i8$}�]�����}��&a�Q~�p�zv��߇��A�i �%_��XTz9&��M#���ޤP-��ݡ��7b6�(e*�6�A>��@��k���0��>׌s) ��m#�)Ē�B?
��ˮ4?�74\��,�L�%E��=�b����"�]�pT�$�'-zˊd��}��	���P��Z�.�"�hZ��`.� �� 2M/7��|�fJ��`	��F�t��Z̩cYObp��T=��'Z傈� ��2p�-�������ƺ����ZJ��# CCI#}¨4�s��*PL�;��]��]��BN۷άm��5���7o\#���~�C)���}wK���yP�+�
rfo)	-ϷfŰ�5����������M�jOI$!]�H�P�����p����OŰǟ�@h�JH*���Y���{V����>�U	سoUq�J��7�g����fȗ��/7Hp��@�w �{S�DKw��O*D�������G��K���I���u��_�v�h[F?�K;%�U�u�L���6���<'a�sb�ɋ��;G¡������y��7#��g����EK`4�p�!=q��Vk��J�+]'�A����濣Wp/���d�����Gs�����u~��iR8X�"F� DD�}ֵG�v��;e.r�$��W{Eh���S �D@Jn�Z�#��^J���&%ཱིVö���C���!d���Y.��A�����霟�8)�����l�jvZ�2w�
��y��<'�f�iHͱ���9S���[���~4�渋�~��tn�\$�f+A>t^�| x��7��c��)S�y:��Xra�9Mƅ�"O��%M�zN��;'�jӥ,)��Xsʈ�"�d����Z��D�ϡ<��i�(z���+���d��R�bVb��E뤾M�e�B���p�M8Zjh=�i�ѯ���`�:D��6v��+����G'�2��q�ytb\#�9.+\��[@�L��f��N+��`Ԡ�Eیl�.W���U�,�?Z�"�� jMr�;�G��N$��I�:�Y� ��6�V"}�y���͟0'x�;���q�<��ܬ�[`a�K�9����u9���!��6���;HSAD�� 撆���#v.�9w�"YY����_Y�+m�i9�n�L� ��!)D� m���w�s�tgs�Cܜ|)�W�V��>����V[S�/��#��(kp�6��aD����K2���l�<��0�pN�HU�������ejv�(  �s��9ENԩ����B3�V�0ǅ��#��}���([�Ǯ��踞�v%���)4��k�xN ����[ꬻ�\Й���&�CF�,�L���RJ�R�puX3*��3�2�Z*D��r���#���q94��$��m�7��:u)	Onۤ4;j�T��P�&{�wsC|W��d%E�D}��[�2����L䒨����D� /����<�˫f�:��� R����}�Nhb�{��
v*�\P.oZo��g��b+]����^�Ny�a����0��}I�ۙ7ul��W(��jB�Eb���՚̓��A��K���� vpU�]�̹�_�;chs�B�ﮙ�~#p�l�T���0nk6u��h�Cg̳�%wC�U���<ĹM[�NӤf�5�w�Ŷ�O��m��i�$A1\hNO� }�p�>�{�.1g]E+����>������	�3���|��9��=��P/	��A�d��3^3g�CI@�1��dᠽ��W����N�vsT�����9AE�IH��|/^ꮜ6�/���� ��U���� �3�������� _�޾���Ko�2oh�T=j�ܑ��É���l�cg�ϫ��2�
�Eh��:o�5
�k�dtN�J[,x�������,�o ��!I�[/�)P� d7��>N����߅��v�f�����ƙ|
�3F���(�K�Es4��=<ݤcx~Q�,�$�1��˩�v���?Y,w�ɩ����p��`bz���$�ϛRӫ�:=�/\���J�Zaf+9�lqe��I-r�]}�3��&I�d�s��k2h���j�K�o��T;�t>~�3L�\^o\�#��������?yY�M�������BI�Z?��X����}X}��� Z�r?]����r����ҥȩN�j���h1����=R�G�>�]M��Iy��_�7��*`t�e�N5[�pyo_��ʅ��]_�b�䖎�)[]�qs�?���x��܄�K$�M�>��`�يJ _���CF9#��!y|�q�R�S#pP�E!�Ym(Kt���#����e.�p1���ҵ�=���1��/��5��@�{���#4�'�o)5!t��_��H��$��¸.�n1Z��ޢ��=�ۛ�H;�c�s�d	M�v9#j�Զ�!@�_y!�(pH��F2dA�XY|�M[�����'piސH;��1���7g.�ņ�U�S�l!u�� ��}��m1�>�'�LvK��yˌ˦%��ѭO�1RvŶ�1���i���U�]�k���+¤'��a�虦�q�ks�����w�[O_�Ę����3{��e���Bȅ�}\��nԔ��= �S�2�[*[����5t���o�k���=��45Y�m6y~hON�˅��QAZ9���G-j�?�a�I�G���R:�|
�]s��EH�v>����k�kR��讄u�O�.�k��d���f0Gɂ�=Ə��zx�g�_t��#/�I��e(�]�	�8�0�	�Ñ���N�K�V	�v�`�Cb��a�c���kNq�6԰;��� R��0�m=O�������}�<!~I�Ŭ�Uļ2I1��!>�V����
e���Om�C�����N�#oz�D�!�L0���o�A.�q�i�+�8�S֖� ��k�6����H�)�l���8�i���R�g�K�����
�V�
����f�'7�rj���,�s�WlF��4�5J���!#	+��&d��~f�	�(s{�n�����̆�D�t�),�=�<�,j)��Vl=sM	����b_�#��A4�I|c��D�t�:��<���Aa@fV�B��us�]lsB��l�m�Ѿ����%�ƺj݋���x��mV��ʮ&��f����⺋�Hߥ3�~�y��B�����sC�w��c��IC�3S}<�|����B[��V��[��j�~] ��(E��ᱹ�
�s'�B���1�����p�»�Z&�@r9��T���K�9�M]>�r<�!��b�C�0�B��:����&�ٍ��A���y��"s�%1m5�z�t=]F�T#� 5�Z)��
���;f/���ܞI��{����	�6�
���q��:Y�[�"�e�汢�T�bM��e���_�u�sV��k)��jL���ݗ�`��ҷ�0�2P]!>��ŞD@Z�"<�ݴ��Ɇ����"s��`��������с{^{5�^Y�XZ}v$����)OE7��,�'��o��\Y�������`�0�������e�?N�@?� ����^mה�fr�G�9���G[D�N�������g�]V<8���.�%�.�"@d�sef�/�?��e>wߨ^G��P	�7sֻY]ўl���I,�o�-<�Kz��{�\ cͫ1�<Y(�(���c����V�{
KN��Y,*�C*�0ԹT��y��J�B�2�K,T���NnH	�׸ v�������=�m���!�躿G�D�#!�����l��4�d�"l9��&Fq��U$oV���v	EΪ�X�ouqI���kk��P�0�������&��F�%����F���i:�v��fRVs%�4z�~��JX�'��Wrۡ�O#)�q�H�h������۱:q�2� R���D�aJP�Y�o�2��14��PO�)A����.>�.ɵP����vA$�'���ޤA-3��t��؂|�d���S����ڷ��3I� +_��S6�K���@���S����jf�Qn늈�pʪ�td�y0o���b
�����3���bl��?�|CY�E�Lk��0<�$�^�и���>Z1�)-�4#@y�VwT&��������L�.�qC=�A��,�ҝ1Q�Ns�A"�M\��Bf�����JQ����+�q���a�pv
u,�Z�����A\젫��~�$]���Y�x��I�4$���T��qլU�{x��OL�-��׉w�7���c�ݴ��<O��ԃ#�f��ȧ	:���z�7�mFWT���>YZ�	�.�Ǟr�����b�v^,J|�'��_�f��u�F�9'5a�D���<�&-Ð���j��Q=��V�7�I|=�6�@��U����ucc"��GR9�e�n�V���>E�)p<��9��=�u}��q��]�o9ě�=U8y$�]�v�1�EOy� �h~���g�
�� \��]ը�P�#�m���V�"Qe:��1�h�5��P�E�(����{��I@Zq���p�� [\����T���~�>u�,r��7=�OT�d���|���h�m�+r�i^ݜݻ�ul6p���X��,�w�w�8Ct!mA@>Wa���C�~q�����;��1�ΘK�M{������C����	����k.�-&���
��Me� ��Ȃ-5�3%V�8kr'�5z��I&9j���<ٱpw�J!N�{3� 1�C~��	E��%�j�݃K�(1.��ꅻ��SF��9�f��JQ��W"�]l�a�o
��� cŕ�_̷,Z9���$�D^F���O�*FPmũ(��w,�L�|}]|�#&��
���MC,���:@v��u��ke�Ա�n�n�</X�v����
:Gl|GYwa��]��Ah�-b`q!�q���~�/(F]hl����m�k�pLԼ�e*N����T�1��~M��w�r��2�G�e�o#�R:7�MOm>��Ў� ۵i��C�z�����6|_��_.3�@c���R���� �&u�}(b�4������@q�܃K�{��ާ%�cNI^��6XP����|�R+I���AIb��MXb2�
4t���91�g���+l4���d�Rw��;��Q̪� Ik���Sqs]�?h��`���Ut��5�.%�T�a���F��Fuh�� Y��`1��(m����A6G�N6�i���l�o$0�Kp��톞�i�/F��P�`��H�h�[�5�ݑ��le8�Q�󾤴Ӎ~a �NM6�Q�z��6��&Y^R��d�m�d�����J�o���۾�����<�ut�Sn��u��ڨ�����@;I��C�O1��!�ܘ �m2����.yG�|�z���z�ݜ1��f�~��(��N���r�2_D�����fm�qEJv#l]�-T.�Νfc6��ŠRya!�xc,#'7����Ŀ�"Ү�2-��`�q[��Ҏ-.��R���d-��wV���C��.�$u\��P�����.���k�t��(�a0��_��4R�n�i�(T���ql�暂��\�{r�E�&�����>��>_�-`F�7��a��3�W��VQ����x�� \��t7m2f��,~�#�5�0i�;f�Zf�͊Q���U�G��B�u+�z֠����_�u���
�C���D�G�C~>�ל�`գV���!�1��㾦Lni})��uC�q�*��_Sw���M�8���eA$���w���m)\@����4��sO2U��,%t��g.b\!B�,�U���_�3m�ƽ|H�e�\�z�|և��`yB,N�ob�<�3o=�Z[���D�auՀ����ifv�(5��h���ųμIv$��N��aٗ�D�L�2�(p�H���̈hG��g�{�.	B�^�4F2c�k!�����2/2�m�\��_T��R$��_�����ѝ��I�5��L���*v�'b���C�e�S6x'?E#+&��[%\[3��[��|>�M"�|�_�K��S����b1j�����N �5�p���o�̀�Z�[�0�p_���vn}�m��W��l�4e��$�0�d�d���Ik�����b�����%y�͹S� L��nKyP�t��� Ҡ��H����'�b��:�_;�sz�E@�����)��# ��9M ���`��h��"x*����>x l_���^��0�a��@�=g=��xj%F1/�fPƖcXj4+��¦)�>?��0�=l��^nc�z����;�&Â�:�b�Ag).���]�!���@�a��ga� ���y�50�<��:M!�j_�0���6#V'��J��N����xc�ȎI4gHڐ�Ȼ_2��ڍE�_�ͣ��}W�{��_�t�?m�:�ϣE��qm�}] �^؛}X��\���@2���G���	�ϋ툁"�ʴ�T:4�]Pض��3XR^�j��U)��8��� ��*�N�!�dd��ϱ�7�.^�n�;Q���K�aTIY��4d�g�jM>����F١i�lr���A/��t�qi�.�,Q!�A��p�=���1=E��I� ���ƭ�WU��p�#�,���'��m*�Q 
$i��%(�UkI�z/8�[�p�礄*B󂪦l�8�{B,sL73��U\�x���|QL(X�u�l녫�=lmnK`!@K~�E���md�(�w��� }�kuB�$ ]�vѤ����`B�������h��L��������4�"J�����W��T�P����:�y@�-�N�~��(H���/�x��x;v�x��P��C�*l���Ȝ���U��ހ�A�%���f���MU�)�v��qP<�H�(���2_�]j} ����E����L���!
U5� ך��K�W��Zt]����פּH���bΒ����xƊ����v����e1����k�Q*����F����߼�Fݶ�(|2v��v���v�i2��g_h���j:ۥ��B;�鉰�4e�A���5G��S��)H���%QO:�ݮ�+���E�+���~�∫��n@���V����̳�X!GN��� [ѣ����sp�ec�_�*���3�tf��Gc�	\TCM׋�>�E��=#q�bk?W�N|�r��h��ûH[S���`Q�����ȍ��q��r�kK�|{�j%¿_�U��F/mF�C�g��4��J�*���������giS���)B�f7�F삓:S!j��c���J���͡L�8�c�g��������ֺt�$���R/��T0�vzKo�j;��a��:?Qd�������G���[��0w�Ҝyg�4Oz��}N�r���T~�0����������V�iZ�dY�3;�jo?!�8�����#�0ǵ�����(M�"�u�0��}\1�v�gV�3���%��S=�E�ȫ%�y��X�/�_<�l۽�
P���Ng��+1X��Vd��/
K�� c�4��1Ce	5*�l:�m�F��\���]�9O#�k/�>DX�Lo���������u�D�&D"�2c���'U���p�J7�y��,/�5ù�A&q�y��YRH�f���y +�۱��3y9>|LX�@bb#ވ�����t�a}ͱ��uL�z>��#w�.(�5^�$�6̃IR�&�u�6�C1�gCx�Q�]g�lm�݆��]G<ғh����h��}�,5M#�`w_˪����%}��1�n��ߝo�fxD�F.����l5׫����O��9�6$!���P�_�T��yC�G�y+a �!�?�A5v"(`��
H�o�Ǡ���sPh��^	���Ct�a���37��%�L<���K�~���	��Any�ɵe�:,�ș:���h���Y5T)�Q/�+�v�U� ٨s%p��+rV/��5�����C�6�����]H���~�[�%C�X-�Q�h�eG ﯋}��:s�,ul(ŀ"#�D:��6����Ńׅ�\��$!]��b�'�@�iq;�C����$�,9������k��x�Hp`D�ȩ�%�!�vz�9�V�I�r��"}`0H{�&����Ǌ�ޢ�}���6��8��hu�a����c���E�4}v�;��_Qiʢ��>FL��R?D��7O��ia�L5HY�S7�?LLw����zNnyZo�j���5�Y�=T���:���@oEq=��pp8B+��:L�>)�7x�g���g�	S���i*��WZ��0��둦�a���ESO�{;�q�B�	{#ᇾ$�+z���S��Pn.*��!��:�%�_<md$9�#'�!G���?�W#����Rö�������
{��X.ǐf�n�����D�EZuWZ�p�^N�{Ll����@y��l�f�H�т��>��%;����A�JU��v��	IղX
���]n���|��|yf*�ָ�K�H_���e�7ޭ�wҼ�I�2�҅E�!|*�`/L��q-}a��+�K��3:����l���{��ˍ���y%�{��-g��e�`(��Y���	;�Zm�eZW�z@��ӭ.(��g�+�'����7 �_���zMժ�j;p���	��"���?�C�[r��YX�BK &^qI�W]\輬VC�V�������#|Ε�f$.��xne� d��mH�D�a�Ք-�X}�}�2R�~l k�l�㻢�W��k�	A �S��e�ǭ�<R�d�A�_�h*P�+�G^��]|TVҀq����M��*\�t{��OC����W�n�	oh 7E���vi�&����������Ze��m$�9���u���Bf�f�:g'1W��<��4���gD�ȅ>��;�a,?;m�H��@ ���{��5|i�4=�b�J�o��)���R�z�/4����^���BRpT�Y4���6��9	�����NY(N& 7H�f�U
�ǥN��*L��%z�(���'��s^?�ʛ�� ��|���� &�_ti���C���x��p��0S�T%��L��֨��^���K��o���ie�����n~��4	���#�Q=��[v"��0����1�����Q�h2[k���~M�w�l�A��t*uF�gr�ؠ�F��⿬�Ms»��K ��)1>{��Dh��o^m�lЙ�)����M���Q��:���G\�=�h��j����#`]��:M���We��7,�?c�T�ŵ6��ɗd:�{%k'��%/����3I���Ϻ���Eie�f,w�)�ژY�?�������糖�P���2�k9����D�4��R%��o9R�~l�'Y7�h@����{g)��s��P�������zW\l�&+�󴿇A;o��O�L�͓�O�xw���_�U��ADd]�6�-���L������{ˣ�ɐ�R�E�|�:�����
q�K�.�j~1uv�Ú!l������-�J�svs���(���Hˍ����Z��!��ݫ��hN̚��Z_����"F�Lôm����nK���&S�&F�K�gn�Z4ޯD�n�w�ИģoS!�GV$s�z���P���]{r��������>���g��84tD��g��w���v��\Q/��~X��:B�y�Xfύ����}���z?���?�H|C�����<�dTxl�~b��J*���d�i!��91wd>o	u�xu����C�����/����K��/,C�D��[�w��Ϡ�;�?5yٙd��k�ˋ������qiɁ��}�P,B�urdپ��٠.��2��h���4t��Kq�w��F�Q�VI���A.�6��r�Ayl0�&˿�B|���%r���T{�#s+$�ysUz������ ќڳiD��f�����K�{�Ǒ����N��-� v�Q���^�cF����q�w|u��c��$�Zu8���f�*����s)|R��T��̘������0yE4�u��\��`�m��G+̗��&u3c��-���ȴ[�n�o sֺW���
4(�^f� [�.ϙ���a����.y�F~ aZQyG)�<���G���]4f�C�m>@�ڜ��a�f�k3��c"��V�+����E��Ro�������gp�h<W�)mS�W�F}�_��"Ro�_��.~�bV�(�ۖ:#LV��0Tu�i`Acp���oN�aL1�G,���"l������T��H����to*�>���u��|��o�QHB�,歍��0)�&�c*�Z{`��i��Œ�L8�N���j��[e��JO�va��i�qPi�N��R�uS%@}Mm�G��J�abg������NHy-�p��X�[_����a�?qfII�8�����Mr�� ��^���4(l̂�R�����]�VV����!ZB���X>d{������|��]���/��,",sC��Y	�'	�'s�)�v�=��]V��Z���P�IiL�9�Ҥ�� �1f6`����3��ɼ�|�{a,��D<���+yT�G.=�@o7Uk���b���hD���q������1@g���k�lt�gwO��7��&ڤ!WϨ7+�Jz�3H,�6�+�&@�R��+<'ה!EGj��%�l���̒L֯!�G�v<�������)$��	cp�LݧL#`�j�%ݹxf�s�'�+)(ŹqY0��ȿCbأ�H�sI�V����<fǲD����K(p�e��d�aX`}U�vl �*��D����n�O{��i	�^Y��%��G�S'�|w,ʁ�p��}�Ǉ����ީ�Op�A+���(����Dh3Vu{�Ͽgq[���y� ^2�kqHO�al���"�r�FO�"c'��c�)p#�;��)l���!���H�s-n�m�9�x�������x|�2t�}��ʰ4O��Ik�������̭�
s��S����jC�N��)q��Bi+��9������AԞ6Jԅ�ng@L
�(W�'�E�2��du���,'h�jyWG:�HQ�bn���¨?�W��cR��E"�����ѹ��t��a����kx�^V��JZ� چb-*v�d��G���U7Q���WP�q�	��s����^F0l��-�w����' �"0�w�l�M;��5ty�Il����.$�A�u�/�ls�*�@i\<t���,�Y�5}���%�1�Y[,�v�$Vb���c��KCu���d�~�ڻ#u,�K���%�_Z�sdI!��V':�h�k>�f �N���y�9���CA�k��Q��7�<&�����?J���\6'�fA	4��¯z{=��	q������"kռ��}�5IR��BM��	ث@��2A&�Fv��m�s�Y'����;�Ұ>�c�5�cgo�̊�IE�^6��f۶p[0d,��Iq����z���V�TD����)%^��7���hG/[!�F*��G�}�4/.�h:�$�E{��ixi"x���#��ty'/
�?�������@��Kj�˒cl���6Z�&�(�x/C���0��~J�����Ӈ�x���^d�"���L>ӧ�����?9T������/�a��@�YV�{!_�i������z��ƃ�������g���hK���h�6i0��ө8f��y%�[vd>������|������&.�B.�#��y���_����L`�`�,=C�Wf3�8��^ESV|wO�b��<��y���yB�0��_��Yv+��*��g'y�'q��E|T�S�+7�>!'o�<�>V'<�V��еL��$��O`h�Ձ�a*"��D�1�3���%T1.��i��G�YL#8���TSVvȅ�H�=��r���P�	�N)*�v~G2>��������T�u��7�����OGm�ׇ��}��<,|�܃�ɀR��4�J����^/�Я��VU��������Hj>Vq�h���8���;�I��
m�Zq�r*8�V��ћ�ƒ9~/C'K��{�c���� 
F��b{ٙF��ǁ��r;_w��>�m{g��t�@R�#���_��+Nl�$�Y[:4!s��o�;7!�+is���y��x��9�b7�G��|��7g�GL�V�S�39SC��n�L.�/L	�#k⥤b��5V�����_Lm ����:i��v���:�=.�L����=��ޱc�Y��yN����¹���齲`�����g9��mK �h�48:m��7�~��O�:C����^n����ޕj5���FQ���Z�Y6��`˼�Om�5��}gޅ ?��?\��`Ms(	T�{�6Gq��-���j�x��g�9�t�C�x`�����1T��,SO��W�#D�1�߹#��1�Z~�0�G�0�Ut��a��cA1A�����,��5�J�=�6��2q{�B���>��b��L��4{��ܾ��wl�0��i�l\�����p/��%~S>E�����=���+R��z���+�CDƉL�`S熖]���iǹ�Un{�LQ����v�2�:*���Ə�C]#,q2���^��y���n�Gp����Y.�6�K�ߔ-��fO�܍�u^�оF�@���<̥,�Wc�o"/6�J����Y��5�{���O�MD��bF.`��a���w"a���������U���΂���@%JhE5��X⋙�'��3�'}�.O� �+v�wͤ�$y���E�g+Cr���%6����4Y�~lGp/���[B܋� ���0��-gG��9r�Wf���n,���W�a�MK|d�x���D�H#aJy���E��K�W�{.=2��PD���a�,�v�е��x����y�^�*�|���X�[��.�,�K�bҩ��0��♖f�������Wa@  �Z���w�c	d�]�W�$��v8tVI>��?��?b���4(����BS<T������e�1�G�l�D=ߣj{�i����W�C�)vU,,7�/��%	�d��E_=N����� åy��<L6��`ގV�I�e���"e4/�㰎�	���j��S�J�9�/R*���_<�L+F��3��xt�=YڒX�1 |��������f��Ck�@�hJs�C������}.j����A�:�vˠu�7}2���a�F�#�ųC�ʼ�{v%���1���]I�t �}�M�B�O�:I_��0%�}(3T_��搜g<��FC�$���BԪҮ.+���S���]s�pX�UjК�.AL��z�����[ռ:�I�q܍a�����a���3�I�K���\r�T8(��C?[P�Y�F*����,	߶��:� ��l�nd�X��y�	�K��ļ�V�Ѡ�����j� ѣyk{6`A�|c��j���qݥ�u�EϿ�f�e��̓�9�V��3B��B�����P̌�-�3�+ko�J�>�71�$�az�FEn��&�+H����E6�+�%�;&Ǆ�t@ɕ��O5����g��}6�"�WW�'sTl��o|���`���<��*��/Y�۞'����49/���)l�&��i�U������(� G��M`��<�Mu��U� |2!Ox��}N`j�k�MK��C:���lO;��b^d�.����[A�2�[��)}�u��a�:E���]�t߰�F�´$ ::	�(��(��N��BD�.Szl��qN� �u�6��^K2O+�&��\��d�M��א	�p�Q��+AI�\P������@��2{<��_�d��OY���I�ߐ����Zj�T��E
�F����d"��iw5Z^ֶ���>�:ޭ��U-M�$k�S	�B���Ŵ�[��|���9<=@�f����0�6ݗ(�t�	�p����d(����������J�'����G���^�����4B�V��t�!��N����N��G��w,@���7�����O8"K�+�1gҪ��שf�Ӕ�����U�ҽ|��e;L(z<�`�jIP��;XO;~��.�dG*�����#hc%�I���MB�g_��f��6(]��x��Pc�6�s�9tj�S���R�Y=�Ll��T*Bֻ��ɟ���d}5�-Ԣ�s �\'���!�����a�I1��d�I�?��{��1 �qP��o��w"!Vx��3
�Mmj�js�	_�J���[Ok�l7nV����V:��v�a��,�4� �f�o����
��r�`�<}GEy�x���	�w�A�ۏ�7e�z���f��T��uy�M̡��-��*�@�b�jB��
�ɐP�Y� ���u}e�7��$>�V<?���M��ȼ+�~��}-�dL#��WC�e����,�evDG�+t����d���)nK�������w��p.���>s��������ib�@���f��pO�rޒ�A1Q��G�(��-Uꖝ�g����d�r��$���y���^���xon$���U�V�GkD݌�/V<�����2q����eI7c�p7
%�-�#M�3E�N��(Ш���#t0\��؂��]>�2j$���t>�
/�z?:���uF��4Q���{P�p�3Z(ޗ���O��R��̚�/��r�7ɬ�2F�(X�;�Y�
&��J��[M�ʅA��9���*6���1�d�V�s��1���p�9`p�޵��cE�T�{�����!���
�9:�EV�xHNh�Ƈ�	��h�L��q�u�z��G·�]0s���Ocמ�B�տ$v��/'|n1�7��w(S�fk+v� ��Tշ����ޗ�)�(y���O�o��Wl��^'�j��l9`Ԓ�%����fn#Kٔ�{����Z8o�F�L�"�9z=.�[XXO�37�t�}]2��9�Ʈ!���&�wb6����I�f�x��h���d��2�f3���x���0��jw|@%�w�b�|�e(Ú�xє�-v��������ԛ1�̦7�=�jE��W|�bE��>�寝~F�9\�[��G�G./����Inx��7(h+@Bv ]hE�4+EZ.�������R�} v��o,�|��A<H]o���+h���V&�r��;Jߚ ��5q���� �@�H�QI�.�r̳J�n��e��
��
>?���x:=�i�]� }�+�:@@�%�R���S�UoE>��5I�ΫK�C-iݑkJ�7���d�<v��:��t�hY7��M�/<���ˆ�Z�oz���)l�!S8�ЖiO��^lj�k"�O���������=���Ȗ+ӊ�s.ΦTa�'K��`Z�!��(���H}�&���gvŭ�������[F��c��z��j�YvsR��M��ry6(����(I��uj�
y��rV��̋��ab�Ɯ�=E��]C�����Mt��k4dm~��m�D��[�*"��o<\���2�,�A#8�~)hE�5�a��A�ڍC&SL�Jh%+G퓳+_��֮Y��I�!�۶�_G��ѷļ�����p��i1�E�F�玛�n�ZJ����kP�!�23�-���=���o*��/{����I�N���c�C?�ی�,o�I��nC�Ҍ���l��k"�?�����X�ؾE��h�q�2�S��}��U	IρrExuS��r2���;���E���l��N���k�����%tp�@��@�b�,9>�����M�X.��kPO�a
"��(Cp��MN�g�w�_��d���8��E>< t Ǿ����D1�%��?���W��0|:wi6�C�������/x�b���Ô�!�(�k������*�J��ʮ"�`�=�K�����K(���+s`��R��rB轇��,���Է����^���rVN�d�|@��Lx9?�!���X���tȘ��G^r��_��E�����3�>��[͓�/Qږmn���E���cG�������q�L�z#9R7s\��|�k��;���)�U���|��5Hv� {��@S$'���b���ϥ8�~o
�g<49���B�'�q��Y�u藋f�sa�n.��yp����Vc�x.z_~�X�O��Z�
*�������Z�rX����8D(�]�r�J��]�D�v)�OG�1̫I=G��N/���@�x����]�piA~�2����%��~��i@%q~�ܲ����GGK�\?��h���I+��r[���ٟs���)�~o���D�bz��c���'��0�`Xق^,��+f��G��a����BL����Z_ұ�:n�h�gtU)^�u��L1�i�1����w��t�T��������=�Eq�|�箧Y8#ܯGi����Ho��6~W���~[n���"~��IrlEE��O�����ͨ�Rpi)��2�ĻR�g��i��=���� ]���VX��TU�ţ�J#�G~y滀��Wڪ]�Z���Rb�^#O�$��F���"�J$!|q܈W�DE6���-�=�	G�"3DR����b������p7?UnY y�R��@�������v����	���3f��v��Y�~���$!إ�1�%2���EV!�X�/���\O�7Cf<v��\�/�k귯'S����O�H~�K�EL�+3��䍿~�_��ۊ���A#|�9�3�_ A��S\�w��2ʳ���j5$@d*.��!5���y݌�k|����ct�.���=��� ���-f��xBF?0?���7��C2�K�ƒl��q�<�����m�W��{5����<��B����E>�4@�����b����g��M�z�U��r]��R�y]��ՕX����qs�g�۰H�R>���w���TP����R"}%�閭5m�;��뗞��96v+��4�`�p-!p!�+Ӭ<*Pnl�p;���*H�Bպ<*Y�ȌWR9O��̈������S٦5Y�~O[`��dR S�������$G���l衯�`���&�&g0I�n�,po�vz� rYO-/���¹�Ҙv�����Yd��8�3�"�t���ת�Cؙ
�Cq�0��Z��}b�����q���g`������"3:�B:qS�c�o��W<mW���tպ��ώd�[�~���|�:���3�?b���v����!G�4E�Ι]�Հ���?9�%��a
-X٤c҇��@�1�����vD�~ڣ�]ܦ�,C�n�M�����B��}r�t���w]Ӛ�+
��5���3m{�B��dT+dU��^-�1�D� �撍yF����YZI좞�,�2p<�K��_/}�K���5�}��F,�F�]}/�.ںxȊ��e�$�dN���h�5��}D�����.e�k��<�ymU���,?�<�IrC�z\��C�ｳk���ｶ�*��K/d&U��:2w��~I����]�{�����69Nb�&���ؗ��z���j䤙�0��_1b���&� \��}�mɒ��CM����UC�(!S��fJk�y����0�0�v�x^K��UI\�p�/�%�7����Q�4c���+�ŖLD{���ƖZ�������,u3�r����pi�U~����b�DTe5�a�c3(���S�� ���~����{�����C������?�}��L����]��&l@���#��vrXy���rqa���tE�畸&7�n�q�R2�z�([<* �P��pҮ6����)��uR���[���9Q8py��o�B)���P{]l|���v��<8B?ĕ�c1��H^D�)p��>�$T�t��Tq)��������U�59��.!B�ߋ<̽u$A������N�F ����t��d`~��iB�`�c�3	�U��[��)'|Ant�0��y�Z����+OЯ���x�6���{T�"�'
�m���_5�xl��a��=�O�:a �ɵú�hK%����Q����fġ�3փ�͒��'�<�>�d=� ����JF�<���벜q6Ö�[�3;u
��t�%7q��(�0�b?p��S���m�ƨ�s��g�{��5��T���3M�}��Z%�J\�ΰK��|�䩊�F5�) ����0c�Y���l���,����f,(6z_���� �D��4߯Y�82M�}�K�w��U����)r��S�a��Q��4ȅ��?�h�:�B��hn�?��
EW	��n ���������,(��������z���N>*�Ѿ���Q�#��-���aٿ���Ӽr�(��I�MT(�Yh�$��ct��рi��5��!r��r4G���( Ö{���x�����'Rg1�g�v�v�����p�g���3~
�n/?�56���gT�4Z�Y;7��&��?������+v��.l�V~hL%T�Fv鳣�
j�����8#_�$y,ϔx�� w�#��,���d��o�'�3���Z3��=f�{�KZC���i/^�H1x�\;R���eT��H��ģF �� ��qj�}��m��Ba��̢��n���|�qj�~�R��d��fH'���AE��X�bd"�c�h�Y�!��+�As�b��ޫe��QY��B+ �@�u׼�%����n$�ݗ�XD2�̇��,_ڏ-����7��m&��"G���`*N23����2���:��ڞ��<�ZgO.�����ܵU-����1��:��?� ��=���Ê&�F�I�������@������9��'5�ʩۉ�P�2�HM�?UTQFvQ����b�5^�b:�Z̀�=I�V�Q�7���G*�юK���g�
�|��,iI���[��*�U;#X
�Ԛ�z��XJ�'�H�-�od9���q�/q�7���+�Ԟ�zy��eV�i#2Y�� ��	�+h( L}�*JܽhJ�W�>��6w���P�]�̣�Bj�Y�����f=��cM��@�,N���qq�����QvhvT,�p�mO�74��Ը�s����9�/�f@�;��vv�C��6F����vW^�#�`�B��cL�j����a>������j�'��M��:i��	�o8��&�K�~.a7�s��yʩd���cmb3,y>��	�0 K1)h�v���Vՙ��)i^˭�-�`A���9u��ǂ]�$��j*/h�0�A��i]mqۦ{X��8 ~:��>)�Y�ʗ��چ�j����z)L�<�E�p+8S�ؽ��z�Q������z�s�8 �OGݜF&h�f��MC� �gc��l�=u�H�c���l�
�%����Z���=�Pzc+C��}�NX�9�G�0���i�	g�#��2-ں�:D��0�ԏR�ŀN�bg�_��0ܛէ�Єj����k�&�|9}�L#�����a�����0,�������DK�QT�m�>�L�{1c�g��KA^hh���Q�5�F�ݗ�{��Dt^T�����.�1LCv,m�i�$�|1H����#��?��L%�I��M����eJ<Cӳ�Q�ȫ��j�8��5���/*�$�7]�����AWLb�wL�*E�d�Ɩ�8p8���LU�A�{Y,jĵ/2}��|�dl}^��zC��ؙ��(���
ZK�4��[�c���2��R�)� ���ԝܷw�X�[��|;-N���.77; k`��n\��	3b�).��Qa~,�58*�ZC�\����K4��&�A��~�˄�w�"�����`�`�~ӡ�ѧ�j/�Z�b�Vpp�h�X*w,�i�er�^��
�N&�h=N��F�I��!<cet��j���9R ,�k!zd!����#K�Tb�h>�@�2b=�� u�W��{'n�p��S6vxv+�p�4�NDxEﺉ�&c��Zt�ݥ(����/���V�~�E��÷�+k��s�A�X`i�N���g�@n	^-Sܨ��|3��r�Q1.��+��H�00W���y�Ӗ��ʨ��F0#}M�Z��,��G(�?��0�"&'��h㱸i4�^�D��x��**���F�\CP|����Q@[4Cxb<�nɟF����� �?�o��wxU�M�~�p�o�*ץA����v��m\L$����K"���P���4�=Q8����t�	��ltҰ�(3q��QTU���c2w�C��3wĲ̘���v0�c	�[���|B��?��p�+%9z��[��	%��i�<�<.�8!��b49:G�'���.�ʡ7�仿�)��o	�ˮٿ���v90C	�B�,���;ʷ���Pl�s���E����q"��X6������[��:�) 潘p8]�.�.�� ֿ�'%2}�Fk�|�:ڎ�8X�9�0/�ҕ��J\�L�����{�b������\4���I��Q�w��Jl	ry^(~�TaX��$���Z��0:��	k$�x�����?;����J�7�6�z��eO��v�BҀF�t�-T�<��į\IS��>g��I� �\��i~2nx1)����|�YJ�'�햓�l���� �����&�dgn>u>8O~��s�
�{mG@U�O�f��$c5�Z�;���lozw���PB�ʼ����)5���5��N�7j�O�R�h\�U�VM|�:�,X���(mB�v��Uf�����Ǒ"�i3J��AHq�D�h�20Q?=�BLh����F.�0+�<#c��� Ǉ]Ry8��v��SZ���
VEO`�tO(�8��T�e����R$�<X�g�y^t1�:t_�����@jl����^s0�:��^� ���$ֵ��$�������>� �����E�8O�<��ΰ���1����|�����Ղ�r�>n�����^'�BS�����
��ZA�ޡsh��E��/o��KL�r<����*}� ��E&�}m�b/*+��V�˳a���l9�1>�?3쵭 1=��h����hy�ǁA"PTʯJ�`a����*�0ԁ�Q80��t�R�׌ ��;�re)R�ZG�S�U�g!�kw����&���Ot�$���uA�c�*-ne�x�Ek5�_W �)�o3-f�V�f�E�)k�{�M�FU�-�z3�.'Yy~B�p_x@6�z�;"��������;+����Z4D�����/3���s3�ϙ�+�Q��1K�6��� %? �b��{?5�Xܛ)���8~�>m�w���ʣ��G3Φ?`Fd_P�*����ʯoA����LN�@޵x>z�����3�-J��l���R`8��SWTy�����>��� �$�G.j��4��6M#d�[z��vIC��\��*��R���ڦ%#.�+uFv�_�m���n�b��=ר�PF%��/�0pmK���7tNqO��{_l�a����aZӑ������m���K������yF�^d�v��`���3!5s�+�v��)���C���B�|ρK꺵�tFk>���n�T�F�ԩ�:A�l� g�m�"nL.�#�W����A�a<5�b �ږG�թArEO"GR'�.a����4}��|��/�#�4�7�7w~s�F�8��%Z3Y��r7]&E�hS���/�~}�w�9I��ӥ16�.'�{�C�5I�z
LK#�d�R�t�u���^nֲ�p]���k��c�s�h6�����G���"-Ad�C�!�:���ܬ��C�]�\Y9V��9����T8�!�vdx�
�n�6��r,�v��������L�
G�P�ɣp�`�K:]-N�W�Kb�ծws���#Nu*YL�����d��!�$Ā>H�{�7���[�u/�?����A_^���mςQ�\�q=h�ul�1�,b;�ћ*eb؂��j�z�������E�JEf2#AH��) �w��ކ�',2��I\����H"uf�VFCjT�;b��̄���k8�
��}�����b����Ƥ�J_ڊ�X�tuUh��QaE�`��ޒ�/�ƙ�k�N���Uyp�W�)m]/8��A2$J�R툈X_��(}�<I��۽>M�GdD!l���n�*��?d�~�[A���u68,6��!�S�ݥ~�K�j-C%ԁS�F�i�e�6d��"�=����k����v�B�������~�3�VV{�Y&]��FG�����|#�\��ݟ���i��h'L�8P�h�#��`�t)��6}�H<�ad<���+u���D�@LHc���O�� �n����6!�����#�+��d@�6x�7��3� 5�)��*��DF_2$c��K�"]�y�����O�]z��"�[�wљSW�V�DVIt)ES�p��kH��.5 p�(oh8q3�v# ��F�Q��++�,n�� ���u�L4��}mBk2KtX��n�7�����@Փ��#�E뒲�Q��׃.��O]v����f���,$g����R/����ޏ���?d�79}�����zNrޮD�N�}W���f��Wm�w0VQ@_�JL�Þx�(7�wG#�o��.V7#¡��^yBؙ)�E��%�1�䪒�+Vv��Lh�1�?q���������-T��ߘ��>鸊�3��o-,ټ|oEuLg+������1�p��j�k��P��;��2�I��L��(ˑ\s��V Ld#�W��x%�@
�nɈ���(q��נ�*��mNQ�e��?b�R/T~�^(������5�ʕh�zi;7-��9�]՛oD���4~��{T�tt�.���ă5�����zk���=Ít��,���r'��R	c�D�JZm+-�,:~魌}�"K�d�O�K
��)��F�n#��@B���>����q>���sE�\v��I9��D����,�B�*7��:�
�/X����>󼑂
�F�1�AwlG=:ien翆{��Ī���o#�to��U��#�����U��	_���$��uR�ֿ�2@��R��I�ܿG��o�ꉥҡ���Wذ��^Y&V1�l��H\ N�(�����*1���v;*2��	�y|��,h���Q�dY�N�ۧ����D��ȱ]'<��VΔE�� ���30pE��|
٧�[�1��D�K�`A�����[��¥Y5��)��1s�����k#j��T�W9a�M�����d�
O�4��jaU�pǷ�W|g�0�xv~8�7��8�lǳ��cp#�'�	&9�b�`�A$��s73x��@q�;��|��tV��P�� ��Wg�	���,7����֝�<,�������E�<l�{O���9Ԅ���궦&����䷴�r�,+,�wA$��_#�k��+C�9N4 ���߳��Aa��M'�2�8s��S��U^����Xc� ̢"�A��hVr$P�R��N�n�E~��u���j�i��U㰹j�<v<ڔ�2[i{��dX��]`JKh8��\����ij+N�1I����~E��y^��Q,��P�m,)�?K�cbX�K��������F���Gx_1YY�5*v�Ԕ��h�>Π��!�x��R����P�ȧQeH����t�v�^�Iy���$F�����}Z�G�.*��l9}'�A��F��c��(��l�B6�D}���H�C�S��&�K��\L�
���ߎ7�o��jm���ĮB�g8+���E�Y~���~��8�R��@�ny(���8ϡ��Q[���S�r��Mu�;�	�V����c �=���;����rd�б7{&�����)�}�r
�h
��Yc�b��"��h�&ݣAt�����Tߪ4Q����
���{tY׺r�h�ߋO�Cd��G�G��GBŁ,^ze`�q�/��J�+�Uπ@�*��T:TW>^���ȺF<9s?�h�o�]��srg�*��W>I��Y&��P�5���3�3�V�(�'�w�G/suNV������c�Yq�ړI�Oƾ�xr�,�� ��U�r�Ar6?Fr�{(�P9�Q|����}u�1�W\�9٬]�7�Re�w��7|�,�dDJ��d�"m��;��4}�'���AOү�&&���)��;�H�Ͷ8���dx��ax����4&�	��`q\�DJ\["�h�R"瀰���`����;mi��'�U0^���4�" P�H�cr��Ed�ZO 
aw V�G�oI�f�;m8h�9����0��(��uK��6N�|GE.u<�@\p�2|��͇�J�#�|��U=���vK) Bd^�1��)ci��.{#<���JV�Z����9�7�F��RQ�0'H��-��<2_Ӊ�}$O�8~F�X�x�&_><r�ɧ��Ҙ����7,�b~W��A�%�E�T��Nu�2JT� ?0��:��pŵ�z4�0j;ྫྷ\3�ݑ�4��Կ�X��r�Ǌږ�S{�\�ܿ]�%+�(��8��w�V�Yf�`��J�+��u����4���8���'dG�R6xG���'���0��O �Vˢ|����o�a��&�\ys��� 6_��s.�x$@�.@:�?�b�QLd��t��!*�K�M{�"�䝝���2�i�?���O��� �����Mu�P��܊`:ێ�7 
���n��t�Hn�G.5�K������%8mǵ�x�fH���Ǭ?�u�B���3���=SI&�OX��+kₘKC-&_K�G-/��ւ���Zfc>�`�ɜ�NA�O��o>:/"�N��z�k��W?O��:X$��s֢y/Nl��q�;eD���t��#9��j���x�56�<��7^���g`�ŉ��C�d�O�U��u������'��^@���n�e\�n�e2��dka�V�������}T�2@��20('.�ɚI~�������s1MA 6jB/_�V ڗ�r���Aro�#��l��:�C����bpB�#����N^��v~m���ʺ_U�9��0�?�tzH�,jUK��OפJf@��VM	�M����:(��K�ʴ��)�T��=��v?,�蝿�ug؎��1u0Z�I�H�Ux�0�,��] ߸48�o���D���K��� 
��EQp�[�0��'��Ұ7�_K�%��N�Rx݅���!����p�4�UtkCy��Pa�>��Qp�g�{H8����7jED��J��'��{�mZ�5�e��`ϳ��L�@9�'�0���A��0�
w�o�"�� �mw�S�Y��X)=�V	��S��c�[��`��XF���rG���G��q�..}�~��1k;��C�C~7�ݾ�{�[�^���7R�lbUci�;_pWXՃ*�}ik6<� *�!���./��ͅ9�+��7ZfCS���(�X�U��{H�%�/5]'X��~�U!͢�6-3vsld�{�F�&�:�C�2V��l�
8#�D�9���q�SIGC�l�<���+­~�g#�����'Z�0�/����$��p�UȻZc��C�J��W���&��u��!�~R���.�I�~�GG�s�~:WË�ӆ�긕{�OUCs��l�ٵ-��B ̡��`~x10���?��J�2�3's�U/Jn:��5ӥ�~���z�^Ĝ�dk+?��G��h"��M�x��A�:��7�=~$PS���p\D��f�H�>"!�v*�2�?9��ٻh���:�|�x��"��a�X�ҳU�6P�΂����{2���C��ĭK�,���/i�/Q��6���}���p��Q�볹�9�`:�/7�ҟB�&��K�0�Z{i�����1mZpFrò�+jQQodH{�}��Zƒ��J�E���k��8N|m8uh���ׇ����޽�ׇx��TY�_����f�e�mt���⿋�*��Yb�2��.x�w�h�3kӑ�xhuA��`�Q�V3*հ����j�o��'���P'���Ba$�2ġ�%B,��ے�hPJ!A�Չ�9,�)�N�ٵ��`E�cWL��?%�{Ӏ/�%��[��{r��-�mT5?��r��C����C��E�կx~�@�ޘ�Jw�͊bO1�>ϴ���0��N��:"*���DF��\ �ٷ
��L����zq����i�c夸�bW�k�3��6ԉ	fM���Y�vE`O�N��r`����k��V)�c�m��}�x�9
�K����A+�9#�����N�Wށ�1E[�����5�m �"l۬�4i ���!e�p/��"��ƥ����Q��7�Rb�u�>�6t��t�3� YA��?���[n �={Ť��\J�\8�OquH�?v��z�?pXC|��f��*�+|B҃�|Z�J��\����v }��.���(���%�U��:�y9���3��ʢ�܃�U煖{���e+!����'��i/)��X��f��C+Z`�8���ǧ6�!&:�8���[���[O��e�o���h�iʳOP �a
[s��P[н�7���r:�.�WZ=a|���B��ˊ�W�5��o� '��v7p��4��P�(�V�B����'�t��K�[4,�<]3$�JZ���i�)F��g��f�e�S�u��y�6��H��+�o��	*�f��ZhϤ��
ѳjJH`�x�����e���M+^=r���bq����z����Βa����?�[�hg�n���ζ{����VH$w�z9�,M��/=I<��c$���~O���p��D��'�p��U��_|y� ܆z]g҉Y�s�q�?��ʗ��1���8u�z�6j�=P�2حW�(�&i��NB#v#G�]�-oA2�&dS�s����t�!�����f�~�7&�m��T����W_T�_�L�xZ�����?[z���n,c���`�k��9=B+D+W���HjJ1/L�qf|@c�es���qM�m퍬�ʡ� ���ZGzAA��� �4(D'��Up���l���Tx��C."��;�����S�)J���6�rn��ɻ����������i���턡��_>����W5WE:�V%F	�.e�ݴK
G5��2��``[�gǞ'�${I?�/�Α�*�)�#�/�f�M�\9"A��@,l[�����p�c��%��l�k�|	�W�
�.ncN���E�ˇ��L�a���N�lAnө5{�;e��%�����%��'^�)²~�!��)nK��81�xԱ�y��ˈ.�#iaH�h3"�@����e��gϬ�1�q���0 ���!�����u�<����.�(h=�4%>��{�@EL����^ 0�Nl7�y�#��oUI���2C�UN�����d�h�\��ޫ��ʂ���s'W���%p��v\Q��)
m �e�uϥVWor{?j ��[GCCm18sn��)+e���&�@z&��T�ҔhC�s�E9�s2n�)c.�k�V�EoQ���BxO�KfY��:�.q��R]O�T2�������pC� ����
�|�T�G� �	�s�>%�Ǭ.�$'BuN��.*gI�d�r>����fBH�*)�7�f�V��j�o�>�.
tF�*�����SS(�o��*B\��&���%� m��CE+g�=�$,��%�C�,N0��ı#��y��4yʧs���0�qw�!�+Xr����٩7�g��vb}��;���P0�����Ŵ>n,����0�pP����o}%��djϧx`6���)�h���V�k���%���HA +%_�s0y���zV�t�5R�O%��k�@�}­�wP��4r7�C��L�L��
Ջ���a�kܦN�9�+�u�b�����]�q6E�+�y7������Gm
��Ù	��|�^��N1!2xE���p�0��i�F�����S�X���y+롵ƽo�.���!Ƙ��tg.I?�����
T��ŵ쭉����i}�ho�d����%��P��^;~��q5��	1�&d1��(5�]���V$Fv��*�⬜��sݎ2e�q��bWa��d
%_���0O���"|1������h��,�d�6m�R�����\C#�u����Ǧ��J\�g���5��U���?��9��\��i����J�_��?�జ�7��e��ٽP"�i���h�g���7�L%� L����c����b�A�T�f���m�*6�D�0$��0$��)�]���B!b��K	@5y�4��4z��M���;�d�c�WS���3��V�G�_?�e�b����+�r`����~D�< ǜ5�?!��K�H
,��CQU]�j���Ia�y[�0a�����!X�9��(�C6�5��[��񟯴Ɗp*w~'�.W&^���"�qo�l���	�ϦGW��!��b�F���i�5]�y,L��v��{K
����B�t�(izA��ufb־=�C�BFG����ļn� �I".�a�J˅�O�m��i��F��s�SDЦ�LW�{����
~Of,�W�M��A���犦�U�zƶN˲�2������j-�^8��ˑ{rX�;ڜ~tk�	��R���%bE��=��b�4!�����O��&L;���;�.ZK�$�_CϾ�
�u6紙֑�aj"�(��|1��˜�T��#����k�}F�fx���B��
R��c�3+��v�ӌ� �xŋ�1��������%>����7��`A��������:�Q%5�xd�!Բ~�˕�%h��T��M�����ػ~6pHA�:�E?p���{N=%Jp����%�kW@����7qAD�v���~w�O/E�XQ�z0�v	x~
90���<�X��Q=Ҟo_�~w�.��ǟ��Ź�L���<f��)f���d�X�}닙�T���_��F�~��5��97���?��ZM0uq(­5�Ϳ��H���=_̱��"/1٠elQ�}ܥFO��XdZ��K]����#��`��.)���d+)�g܃_��Y�����#{T3}u,�YQ�[#5��ŕ�*��+\d
Z[���e��(,���ܞ�����:��[���2 �a��H�
�t�]����[}�Э�o����v���)��.��l�H|H8�u���=�(�h�%cn�I���RPRb���Bm��6yC��L���I)�/0|���f�2D	��T-Ϛ�(�m���8A�;�ȣ�w�r��k���qN�������nrg��b�s��T	u���� �-��>���d���[�8��RG��'��j5%�u
w�ґ]��&4-���~}�#Џ��D�O҈ުe��,�"�ɱ�@>Q�-RB�m���ǰ�/rb*��zf�z�����,~�h���G2���O�		�Q�e��טD�%!�x^�3Q��9Y��?4Y(f�q��8{%�=�`Mj/c��J����1�[��������B~8]X������Zj2Ѫ�=��ӓ���	�eٌ���A�鮠Ȝ�E����l	!�X�_GT�/��5ybοk�A�+�?����jׅq#������A��S�$�E��ћ{�4ԯ_�Y�'θjo�|gED�w�j��[��QI1�0�E�8
3P����d�M��
K��t���A&Ԓ��I]o�_B#^\R-���\��N���)�q~[�t��e����?.��?��Z������n\r)V�Jl�I�Z����j�_��ۭ,���ts�0�ks�l������T� �0D�T�+���K�D;G�Sl�ʡ߈��;��΢R�\��-Z���f�0�=ُ��׊},d���zȒ�jn�a�P� C����0�Lu��i��-|Xz�:�#S�1W�`WۧW�?�b���	E������K'��ズ�|�����d*NO�Ż�^Ef�1~H:ӆ��p>�	� :.r~+$li��&��i����^��
���T���q:����5���L���f��ƽUT�����a��:F��Ɵkq�����B��Xޙ�k�T�*�%|���蓾�r�u����ۀ,!۞�����ӷ�U>�NZτ-��#Z!�Z<&��R+ �w�݀*�h��4��Bv�`0�0��������6n��r��W�o<Yh���RW��?-�4v+l_G��=���O��/	���wV�Mf�М�y��Ʒ��Ӭ(ߦ
VS�i���N��Ǔ�u�m=�(��Èa�Ҕ�Fʧ���nv�	�]�R�<!`B�𼓊6{�ᙛ���!��c��;���pQK�O��0ҏaQ�d�U�$�x��Ɲ�Y���E�m��[��RS��e�j|�<���;}�Da1�M��]��i5�i���p��;���ǡ+g�ڤ��Q��,;[�|�k'c�����~���Y�JS|�kT��6΀�!��[/9��a�p�y����GPA'�3LP��![&,��N���[)_M��<�q�x�KQw�1�$2�BMV'��_g�/W�h�\GS����N�#0w(f�\��W�#����0Ҽ_�S-\�/"��)�r�s�-iT��4��H;���ޞ��Ҹ�H#v�N�jA����e���Ŝ�֗�\[����U��3�ml��}�$+����.��Ĝ�H�:���i;��������%X��B��'_�l��O���j�9q9�R��-�ٚAz�_��v�@*�E�]���������LH���u8����S���6�ny�^w�YeS��Y��`6�ᬝ���ɺ?e�QǏ}5��D�"+c(��=`9(΀�I�ާ��:�1p=|
z�(� #^�͎�YE`�j!t��5Hg!?RW�vV�q]	�~
��K� 	�Q�X!A���ab͚��o1��F�_�q%�t�<R>_�4��kw����cWa%���5��\Q��� �6����\��b#E���w�<>�כQ�>��S�7���$Ƥ���|��ښ�6�J�(��DF�
��ͧ�)�Q�%�t��Y�%�5���Dȋ����$���ݭV]����]r��Wે�4��W��3Ti@�b"�4 ��х޼	.������/�lI�Ȼ-{����)ݴB��h��h���ݛnm�*:+��$Iy"N��J��ڧ��>
�&J�V*hW�'�Yi1���xvE�3��dj,~���=1�V�����q
Ǆ�����i#�q#=����c�!��nO��U�
��E��"a���2�F�.�j02�]���hy�̛A}���Hͦ��I6�=���%5���P�xS�@-����G�;�r�=�!m3|W�,��D��g��#��i�]gD'[� �yu�����j��K|4�J*�3�����ZR��������+��l��}!����f������:V
���փ ����� ���S�s�?���H�Lo�2imM�Y����9�{N筠���9W���z���ɶ�wX����&�+��	�ȟ�÷��V8ҍ���F"���S�|w�HkK�e�n���ᓠ.t+qKCA��*����ۖ�i~�䥷��<ĸ�ܸcJ��7s��%�<%��xEr�#�����U� �U��Ӆ����Z8Yp�5p#.}~�ڊ&%�(e����h����߱��)Ŀ8�К���.	f����+˧W�+� W��z�$S��|R6�i.�W+��a�';/G�-���9G� 7�|Fo ��=�<y��Έ�
8\��ǡ����65��m����p��Y��?A���+3/�C(��%:Z�;�l�I|�ql�����LR�#�aZ��K���}n+Q�2�/KC��Z���G�f�t�8l��NS�K��vE��m��>�A��6��_�[�4��D�j����a�H}e�M��"{o�?Ԟ�
���'�͒N��熇���z���"�rW'^��w6�E�:&]�i�>�&xS1QV&
�p��5$hŎ<.�#jn��Dc���6�.$�(y���g�X�)KQ���{��5?���6>V�ݟ�z4m�o��0�i$^�f��uزlQ$
x4��q*���
�v�/�Jh��ۖ�tz �|Hw���DP�^8a@��'zs%���&1�ҷ���ͧ�W:�+�����*��k�+���֩�wu�p�I��F���K�9B����ֳx9H����� G�47H;�U8�g�W��	2=�*m��C<]�o���SH�n݈��܍2?{��&���C3�s~��2c�5=٦��3� ,���c�z�5L��1~��by�����L �Cۚw��$�����􆦋�o!�%��͋����/��� ��^p�7�Z9&����Ǹz)=�t=�D)�|b�%%�ʽ#DG -7i�/!�(-��F�&%lt���A$i���&�<�RO׀z���Ľ��"-������ݨ�Ε�bŌ�?��%%���\m�4�G��0��r��zw�6���/��ap�t�����D�D^�>�\���|S�������m^\8�����6c������O淓��ׯ�0�_`��y%�Y��ŀ�m���(99�`��꧚��>i�����1��(��[s�?b�z,�
��
�2|M|e����cƫ!�nK�^Pݤô���|�D��?�U������pE
�T�D��A?��b�g6��
���ȕ��kLD/�n�%������ߘ?96X"��jA��u�C	JV
ܙه�`jQ��z�Y`�����W���փ���R\� ����`5��	���u�u����qYA��SZ�,�HB�u%�����8m_,��q�@T_v�'�q��6�U��������"��(xx8�5�_C$.�l�Q^kkD�[�x,�h����߉�䔺�u���C�0�d���iA:ҚΜ3V�����M���@����Ⱦ\����Y��V�����=,�����)T���p�8��y�A6y��}�GK�Z��S������+�%��^"8�H�
[�"t�d��·�j�������������]L1m=��% ��&H�����
~k^��G[�����Fy����?u8|Nb�l޴�N�P1)�Q	
�=�"l5�����n�I9Q��ՠ֤�@:.���g%���S/wJoʣ�����?����9�4܁{M�e��J���ا�J��s��"��/�H��$Ԗ���hۘD&XXb�7��%�N��k�{1�R���}%Oۧ �%cy?�@�Xk�>�mޭmQ̆dg.�kj�n�e��ĸ��ѐ��������sø��-��[��3����6��U@/dQ����5 ُ��'j���̌�y/�&��Q�y;Nm�$7�}�#�V�F��x���aף�䖧6ു�9|��f-��Ue(��K2�J��T�(���x'�=�b9����`�O������,Y10=����cD{i,��*�tI��;#\Wd_��K� ��
E����"�A��#�ǥ��ol�� veZ���{�ߴ=�T��(0�O��*8fM�:�1ܵ�]���齟
?��@DXv��@��L�
h��懑|鹋Y���`��k�^�m��;<�M��=_+^/��zeS����E�S�֡	���0ߓ���k�3��	@����z1\%�ۉ�Gw���NbS�)� ������R��kBC/;a�z�l5��TK_[f��ߊ��^�������V��_����n�ܳ�dn���u��Gg�x���s9��F���3��풥���{':���5�C�k��{�H��p��
2���%c�7250WS�$٣���2"���QJEY�I��d�{��3��E5D��[s'�?f��}��Eu���������"�d�~WnM��,C�bE~��	�Na
qE]tD���!�W"P�-D��8H{px�%Pu��Eh6���Ԓ=�!$CI�VrPD����e�����m	;�$�P=u���m�P���jk��m�WY�-C��u:O�|��"0jD�W��0�{?��*��g�! d���ja���<E����u@eQ�z[�]�Z^]P0{�Yx0)���|@��߽ՀKр�E�R��|4�@i��h�Am��̉L��t��f�N#d�jV��6_1��2�~��g.`ȏ��F�D�v��1%Pg��a��[@:�6��p�vSwG�O=Q� 6~8A	��<m=��i�N���fr*���E����s�&�����`�4���z����A�9A���=Ӱ��p����nB����hIB�D�!����rqW�~@��׈��m��)V�Q[2���o-�Q�(�T�Se=�X>��0�j��� E����@d�b[�Q���*�mC]ss �����;�����q�6��u��3p��f5�Q�+m�t��g�\�WX2XLt�ѷKOl#J7��~�8"}������]��z*m
g;��g��Λ�E���8]�SQ���[Γ��#�2�S��k��~[�QƤ�8���RU�����}��<Ld��
��^*BD���O����'9kh�Z9r����v���d��I����C����:&P!��%Rr���7��J�?���0~��5�M�{c���o�n�c�d�i~H�fx��|�p(F���C�'��E,{X�ٞ{��X���4a����I�o�����O��Д�?;��rӊG^�F�E�yoMcv��ҧ�τ1�#��)7QG�x"-��d���m'�IlD�$���5|�݀j��� ȓ�W��vjfG�8eI^pgE'����؟Ŀ,ZxK:
��Glfm�d��7������u�[?(D�L������I_V,	��~�ǚr,�Y���L�'�<�Q�A��3Wy�8sO�c/qm�k�Ԥv�QH�� )�Jhz�����)���@?����7�����l�ۍ�����қ�TԢ�b�G�=�\�P�m��q �	��vS��b����Z�1�g���� ��0����~Vnk#����-	���d��N��m?;�o�����i3��^3c]g+Q3X�7(��)�Ү�Qĭ�3�1"A^;��,j����C"p��b��7/��{�F�:���ۜĚ�PÊ��W�p)yA*V�����I_��:C0�|��yE�S�/`�)O�T�q�:C!�&�hܲ���Ǘ9�塡1=����5=�����4��\;F�E�U";~r�?.��b�<�����s�р�(�UI;M�qmg��el4��3h��3ѫ�w[ջ�j)#P-2	�G���\��>8H�28S�q3g���s�. �Pءe��n�M�d�f*G��ߌ�$}h��.�e�������5�S�<z��	�qБ���ϣ���]���H�5�f>I��KcZH��R��47:�Ő��p�e���f��ԝ\��J6�s�����ҳ����8�Fx	�3|��5T�j��F6(3�g.�7M!�1i9� xӥ�z��[M���鶫��{�i5I��P�L��@t�.�b�ӱyձ��ږL���%J�l�j�l�/��h7鬳�tN����GqO�s(�=@@�A��2Lj�㓓H~�c�� %�m�m��N5NH̯��Q ���6�?"��g�T�f>8-H�U� <phs
z��Oz2��`�޸�#�	���I�/D9�<�%��r��M��"?zֲ�DZ皁�j�%�E��s\Z�g�15���|��hqu�u�Z�K{gN.x`'}q�W<��j�C��G���G-����Zq��.�ҍ�E�Ʌ�Α���3vp)b	z����:j��C	�SrFg9-�J�h���VB�.4�0��<��K�K����TN�����Js��a��A�gW}yW1/]f�����9�ѥp&���`U2K�)�E?1"�n����������*��x� ��%Z��z1�	�h8X�d�P���k8���!�J��RO�W�Tvʟ��b�X�0� f&�baYi��W%@Ĵ���Wr�}U|dͷ0��n�>���Z/�<Op��G]�V֝���Ht��U��"��aln�Y�<L~*�H/'�#U�r�<���t��T/��D�T(i�܉�7�Z�����MU���`[��;J$5s�,�4Y]�FϜ�����d��7(B�;�eEu��Ͽ�9��O�a����fb{���|��ʿ��1��X�$�bnM!�ɜ��ί�;A$���� p��������'��X�hh�^���®rKu9,��t�0��U� Ǳ�b����T�y�ǳ%�,��b�!�Q��\M.��u�ZԎM��Ɨ��B�Z�{5�������s�r�R���)�HD��}�AjP=��B��������Gy{/���oǹ [pt=��[�4x-ܞZX˷�ےW�*dv�2KYq�E�j2'���i{��tby@oD Z���n��&�"�'���R�^��'�K(���WJ�έY�\�?�7bR9h�)�&��J���q�	�q�y;O�b����Oܥ5Λ[WDY<(SvD�����=��޶�u�@BM���/��it��g�*mJk.�����j����2��n���U�D�O$�3~O'ZЄB�Eov~h�b�A��ϣ��Aߎ�����\��Yl�t����yΡ��fK�s�/
8td���H
8�~��$��3����3t1H�>�4�O"r,���4�*�{�/�D�s��2��xx��TG�i��� �^�P�������@�I���Z�fg���9���i���z.��]�I"Yk�rmK�k��%�4q]�� 8\�:�Q�g�E#ahO�Z�x�2A7y��5��P���1�;Nx�BV�?����h%"��ѩ��B�ҁz|Y+S��6��>���n�k/�Y�mrt�]:5V����VT�8L�u�g�Ⱥ<R�)M�mǈ?V5p���~�ٹ�o/���z�
M���kv�g���+�  ��:Jnӝq'��C�Ρ��ᶡ�o�w���I�°��X�Wy��c��Z�m�i9��qЫ<��7�3QF}1;�K��^n��^�v��{#���,zQ�a�!�C�b[��0��ՙ�e�<1�(56_���!�Ar��fأ}󿡠����e:��
1�\���F��`�"ǬaB�����Aq���'1	�P�� �4-#WU�x0z��l�GZB&|����E��%;��"(N�^O*��R�JZ��OB"ъ�� ��ehh�Ԋ�N �=�ȕ�9r�d��=f���)w)xd1ڮ�y��n���4��k]��1ο�Vgo�8�%}�Wm���(��F�����4[6�Ī�{s�2���w�����(A�A�sgXWH8`���hq��$^�.����`Ȓ�xK����y��{��X�oh��(��ۢXˣ�
\�#��Ӧ�h���'���g����q���+c��Pr�{�D�T��MUXą >(�B@���
�|s*���K���%怔AL��ރ�,�m�,ׁb��4���fU6O�.�GF'O�Y��}9`;Q�W�K�^�I?�1�a���o�A����x�YR�ǃ7�Y����ц6�?}�7�����m(�2�<��<�!}S�$�Y�� �p-���.T�<����WO?z!`On����$[M�����	��Q"1y���i�!0.��!�<�^��ô4�wc��.4?��c��1�y���A�҆�F\�$w��́�\��r֢CF��@I^��T���-���z �`�`���m�pn�^���f�7�{GC�ޠ_�΋jj�E6��f4�5�
����-��|c0��.� �x�L�E���̀�m�����l8خs��{�e�!��#�����L��IB-銓��q�g��G�O�N�'9ǿrW�f�פi��F%��9�M�s��9V��Q�:p,x���ˍTr6����^rz��|P�@q�*9�in�A���e7��e
%�`q�=�a��y�@�$\�Ij��h@
f!�������A
k��D�de�5�.��ǋ�*{�F�]36j7�S��1��+�����[TǂBF^�C��&qGэh"�Y�xQ		��x��MA��k��.&x��U�\L���}�����W4��\�"�ȅհ�}�Es,@gM5B�G��1y�R��ƭ>.O���pT� Fas�WH���k��ZƦ"�h�+�_�YU�br �0�
�;�����I<��|�Q�R��u�q��aQ-��&otW��l��KC�����|��Χ?�9���wЦ�v��x�~.�@�{��h�˻��qt�5`l�k��]b�*�=�G��uy���穗2A_��xxH�O��߿�P'��#=>��@\�9rF�~y:c����@����WE����&og�y�p�� IK�b^&��+#
����.���G�r6�jr��f hG8(I2�s1�ʭ����>�&Sw,�w�xUj�3��Nےh󈈤�-G��漏�@�[Խ�2<��� ��K��膪��4�?ha�!�W�q�GL�� `�|�KR�KQO4�|��`ۉ��\3�m���1��xﰧ�!�	�!��UQ�wַ��R���O��*���z�����k�`z��W@�_��T ����yM�8�<��y8�S؀��2�o*��"�-�V�䢔�i�~�(�Y�8�&�5��WƐ�!ct�N˾�0mzC��!A���᫏*V����ܯ�=���{���x����'z�os	"��+OH�d�9��d��eM��b�Q�%U�|<�=�Br?'���'�.!��Tf��m,�����4\t!{	MedA`�a�� Q�w톆F��*�r��F�oԹ��:��|*0
g�K��â�F�̯���m'9�bU~�_�i{��l�p?���n��Ǭ���������">W]��k�����:��_(ޒx��`���B�.�Yy�X�4;���SG�&"*�V��^��x`ƒ��䎟��T) �+/a}��O�۫�����bx�,� �lN��s���r%S��
VN�o{���(�R��en=�?�P���z��þQ��}��b_�3���P1\�}�]���X�]��J���4���),�E�C[���}��̈́�&���H�O'��m5"��DMhI�;��
gp�$;P9[��ܷ3��,!�B`��ZA��\		�T�,���-I�OI�l�0�W�q�pRf���%��;[E�҅w S������Fmu%�������y (��<�O��_�Q�]��5l�F�0�k'��+VR��B���b�ۆLC�j:ar�;Pv9E߷Ti���n�����t
Gwem�^�*y�;o�p����X㦜+L�8���Y��._����_���c賷�۪J���K��˨ERǀ��ߗ�~ط�#��p�-Q���m�͌V]a�mSh��V\��<�';�=�<�J1j:��h�'Ӡ7pg���y2Ym+��5�m��;����*U�BU��OLE���!���/ ��T+P`޾Yf�J&�,̈��.a��q����2����D"�x�J<
����Քܸ��:�"��|!)��+�7?�@ҏ*�'�e���&jv]Z�Ӵ��zu_��{��:&������cf⠨N.3��>g-|n����u	�	$jx�pC��J�{Z�p��ũ�Y){��W��q��7-�hj@�j�À'�5A=�b쐞]�wF����,"׷}k9^�k%*��*�v�y�1� 2dh㿗��`�4���3k���y�i�����3)1��C�(,�M(�'�S_����Hق���!�Iz'�T�����1�ok��(QDlU�^�[:|D�&�>IZF�7_�{~ߩ,�u�w�{���9RN�7���<R��G{�C��,>/��cdi'>��ݢ�V{?YM��g����Dď�kJ���Z��V�$E�M�f�L%�����5z;��+�Se�S(�;C!�
��X�� �.�\�űu2�m�[j��r��5��� S3��FD{+R�[]z�2��z����W.g�dФ~��?O�+3�`�*��N�ҦS�޵�@a���{ذ$�%��4��L���6���v*x�8}������	5t;Z�t:��r1�}l~��	㘦��ް�+l����ϼ��Y�zm�q
�Y�Z�RUv�2��ĕuQ���6�#��?� #.S�J�@�(��j�_�g��3bo���P5��P��>e�JQJJ7�~=&y���v���鐦-�~���odޔ�;%�ߓ��<M�����7�a9��E��B�	1�4Q��
#��3��hS��YZN>��>�e����,���Z����/��EAp���ćy挊�s�8m�-���]2櫝�;�aվim] oG�<Ig��T������A0�c��3�Ҩ|�0H1���-d��UlF"��^�*)]1�^5�H�z��WYS|��^Y-��Vz���P�H��^�Z����G��B,Ö���(���.��z�N���[-�8�*�Z���!��������q#X@��7�!������Fv��(Y���߈)��Y��,7Ɓ71F��uZ��Ow����}Z��&>&�INz����ؖD����#r��b|P�
�1��C�5�I�a�N�QU�su�+��=��0��@p�d%҆"��ˀ*���֒2BT�`:&t�#G��*9Ҟ���~��z�~$� �x�S�,*34�q^����̹#�_��Hhr�a�VLO�V�q����b��I�b�o�L����.��'�1~���}�Da�Я4f�nf^lsP;$�S*�w���注���r>��R_��S͵��d �7+�p�8{�B�C����<y�ȅ�c¤����@�_5}o�FCG�Z���?�.��������	J��EY�[X���~��p3�6�˜+A��͎k���\���g5G��1���b޲���M��V<�
��� k����JM֓ǿL0�R��{Ť��s<}�E*�Jp�F�7���L�7K��?Q���!����HZ^������9%ǽ�U�Ɨ�׸�c�=[o���5�A9�;�w��ly�m�W'����F��PK�����#�".?s��Y�=:%kX|�f�C�K�p��O��:�&Wc�ɎHײ�@�`Mq6??��"�A��KY��� �~�,�ߧ{64����ޏ�H�F�}���6[Q[V��u��9�LS?`�6Z�#gڃWjs�G1la쮫�M1g3vq��Y�6.{E$4��BO�4�(�/-�{��en�އ[�.T�ZL��|�c��;�8y�.�R�bB�L��P>-#��nl���8���a�����-9.�ǷU����o݉�p.]a��{d�<�ni�D�j\r�/�\8FN�	����bY��RE�8`��T�s�����������S����Mi�O�-�Cxy}p��`�~����Q��A�h�hsg#�+\*0X\�.6�«Qm���X>� ?V�޿�g�L<�a�`w���Cd�t������$���L\8lѠaɞM���M[���t�a�ߏo�m�����k%��3A�,><G���E5k�>Ü/Wt�K�� �J\q�$d`;������ʾ�����֦�&R���]��+�����yv-Z ���E{�O���l-�a-OX��և���]�e���
?E�.����)ۉP���Ƅ��H= 3S�"�5ci</�rJ���U^Hw[�}A�s�&l�_�]�jU���;&��Fnq@֋%�S��_�ǟvc����9ҟ�� 	�����2��z�$���)�!ҟ��5�x�Z-�23uT疭Qti%R�Z�f���O87����N�w�1���p�� ���}!mv�-+��>�1�^�$�xF���e���}�3s/�Ha��b�7��z�
|�` �Tl4ip�M�Q��0�D�b�`��4�s:�*w��bBn`�ȑg 
48ՑP�FI
_Rl�o�U��uY%���^���f�+��*��,��Wx��ߟQ���/�c0�@<�T�@�NpN�_�>]�T� ���.Q�<{e�SuE���Fk�>�����nM�ĵ#��c*�C���3|�It>iAЦچ�Ky!�Ŕe	5����
d��o��o<-?-�eˊ�P�9$�s-70��X���ΐ�݉���)���+�gC���C:ݡ	6v?T]�ﾽ�mrӀp�^u� ��)�L]�2"��Y.�����~�L�&T7�v� �m��(��;f[�;���	��?��0��Q�b<)�D��q��͚\�|�p�6K��g��&����ޮU�G.r����aB<�%�F�ؤ��S�%�c�3�@���.�h���J;�w03"��
��_������Mc*�9ۮ��x�S��9�_aCa��i���}����(�m�I~4�L��ł�ݵP���2�5;vt�lܚ���PeR�	G;h����d3������'��I�8=�G8ݐ�1F��	Z�C3qw��[l��ɉӽ��XW͡obCi[C��r-*�&�#�)o*�zf
3d}��d�w�t�'.e�Mj����3Ϟ�Ķu����(�*|Z�����0�����Y���������rE���f/�4�K���?�H�<�IO�E6lG|~���p��Ҽ�
U�T�g�ȯ����SX�;�w��Pզu����$e���0뢏~M���~�-�w��뛓�j��Ѥz��u���9`�H5J_�2�n\h�iL��A���LI��N�7gD�ݱ�\��<��Y_^�q��aHq��|��r��v�;���&�S����������%ҷ|����f�'MY�׸��/^'��up
�#*�jq�K�H�1Y��M`h��5�����Jv�'X��+��l��6]�g�Wbn����p�k��ƥ��u����ױ�m<�6���6�'�q[Z��Bj5v�z�j�`���X�S�U��q��b#[��a�b��|f�þ��3im�.�%��\�Z�@ȷ��	˙t�IJ!6�����z<����0��KMWd�z\�DO�ئ�Ӌ�eo�c-��L��P ܑ�����wdUr[���a �=��ѡ*�"6	hw×�O����7B�	��C�xc���ƾ|�4�� `ȵ���L�Ns��i/���ݗ�bVU�5�n��&l���D>��� �O�K��vp{9�9P��� ��i}�XM�e����V��ƭ�H��MYT��JՋ���V���S�A���ބa¢�pAԴ�X�Ĝ3��iDk��L2tШ�"��U�S�<��'�`���?��*LX�]i�9��/}�E�یx;��f�����!��M�ю��4ź|m8�;*����Ob{l���\�j��R�Б��iف5'9�W 2:�h���i�n�F86��XD^yJ!��r��2_�d��N��RvO8�PO�s�Ԑ �@����[�<������>��)z�w�x2O0�w��d��(�'�ȥ�wz_A�bJ�����s���s3�C0����,T*�X�&�N/��>?;i����2)L�4F��nDC(��Ιm�xօ
X*��Y���ˑL@'��c���,�($�Q�˔ c�)*y�ӞM�X��uo�@)#�?�jٯ(4Ru{«��2<#�6M��c��+͖�i=�-���!�'��.����ʂ bi��s%�^R�o����Iu��i��{�6���s��CDh4��_�~�C�1i�U!{�FN�mޥ0G���#~���4�۸���OR�#���ɑnQx��[1x�u�� Ulb�N�����=i+j\ECDN���\�f�x�௙�O[Aŀ�x:��#z?����|����E�w�s-����	���=�P(2�[d��Q��b����,���l���W�.$�[C��#�=	q��M�:D^z��m�����W�)*3j���g��[��h�]� �����u1xzq�_I��zK��j���/�S���@�/��d���^�߅�I'C�O>Q��,���_�c�ciB�&���?��IǼ����:�y�# ,���ॴ� J�����'k���G�&�,Arf[U"8J�ƁCV�_Vp)̳�5j	^�KR �C^HJjh�o�vg[JI�l�W�Ȑ�qu�LT�d+�l��nnΦ3+�E���lX<���'�l�6�wB���@,���5�(���L�\���]8O�k1jf�}Ǣ-�>2�)��u`��:��
�����{��GE���:6��Rȣ�}�6�ǋ$޻�����L���bz_pu`�_o�q�p�ӛj��,��*� ��WJR;`�m`�XDl:�	��6Rh���1��#7��u:GW6�gv6�It��"�Х�OYM���%�>Q�ǖA��F&����^<e!.��t�MK�cs,��7Ǚ�!ٺ��ٌ�bED�Pi�t�|��8�9�h�}��哢�@�Ɲjr�����2"4�9�4.0T�5���h��$�-(x���� #��?3�-���A�}�0�S�u2ˎ��^�!�����ň�nڪ�&)A>Q���!o�3 �Q+���?�V�/0em��b��^��B�9�<��U�=hź�z��.V�R/��6�g#ٗ��O���w��o<��>�f5����˿W�=٠�BQ{�ڞ����$�ɅJ:e�)��nxY���Yo�|��q DRt����Pcb	�m�/°z�{�W_�<�m��o(1��{L�~�p���eݟ�h�Qau_���1�3e������8�:�t�������gux�<���I�C1��V�=D�Յ��+$�Gfm����h�K�+��zg����oR��|������7\@g���
���z�5�A ��C����p�Bf�t�ݐ��Р;����]�kb叾/��9��ۡ��f�,ʠ@1�0�di��6��?~��Ǩ]���+[ݾ%�'�����%o:�r�����	���2�J`�q��]RYM�Hi\uJS2K3����v���LlTB:r鈁ɍ�=��yƹ�*������I�%A�(�"Hb����r,��.JW��\����8���5U��YVe-�t�.�ՙ����8����=�&�����]��cs�[,���U
f�a��"X�ց��F1!����|;���`�tn�8�L��4�"0c������U{�^��u<� Iа'�I��s��n
�OV�B{%�p�B����2���֣��c��ɽ�[����=����W�r�W�Z}=�6(�@����I|�-�������ȼ�D�|���r,U��'Ba� �濝�� 񚶟��k�5l��x�6���L��VMN�ZŔ�d�I�n2������[�|��x����
Xy{�b����K	S���O�=�I��]��bwp^Վ)��T�$�橚m�mbT])�_�!��ٶOxb)��|g9��YO��u2��_�˥L�h�O�q����jv	�Nb�y���
�-�Cj*���w��\��g��v8դ�� 9���^�D��i0_dw畉�iWO7�Pc&�"�����~�Ύ�,� ��>��e���2����N�g�[��<�		ɒ�4n��������� ����O�vhp���!�R��8hz|w��`t8=�z�s�F_�-m���`�)[�xz1�Յ^�~������{M���=L
�KlZ����~U��N� ��
-�e]Dj��T�T'��Q gR"<TU�S,(��
*�b����i�{���"�՛-�/�m��]���bH^����d��G��3?7��}�w�A�UT��5^l^5�9	���F�P���H��dZҪ%D�.x�������1�IEz���/�\�v��v(�'Ķ�~�A�!�LKd��Z\"����%�DM���'� �A������y�B�������t<eY\���܀Z`��>��o�{]�'���Q��/?����<�.�8����3F�]ݐ87>��>YJ �E�s���$�[z�&�ҟ��qv�s�h��:� ΋o��er����_1S_�1��Ώ���'^�@%�(YHR}5"U���m��?���JQ+��	�41��n�"�j���(��-ѡ�����tСr( �F����^%��yn��{~�d5����֍0v�C.��8�� ��L�`��b`����~��w��(�@3��(��$v-[IB��ߣf�,z�?B��f�\�F�e��pDY�\n�WPj��:�3B��ӥN�N�4����J{�e��Tl�������0,��Z&�{o�K��9'��|�|q��=� E_�n���b���V�Z����P��%�%gZ�T��k�/[������Q��H{��Vί
�aP`��s:\/��7
PE{_�PE莋�t���'��5
�2�/ B�i[������D���W�MϜ�Ce�+�(���m{�����֮pz�z�����ʭ�hNe(T���w�I��˞0��>��ŀ�ܭN�Z(��D���F6�{��D����8��`Ngn���hC��G�3kP��T���|@z���ϴcje�K�4_7��Xm���m}�,6��d�6����?���c

�&�^��GÔ�F�o��j����8B�s,�Xc���)3�tעs%Un篃%w6�dȆfaB�ST�-���%���������?6�,�=�Z'����1�X|%�` ~P�"}o���h�z��g�ߣ	_c�H
�em$F������|��*�CI������jc"gv;5bM��Z`�G���b{;&�R����oKs�����L�����{��}=�xM�!��^��L�Ὢs��H�;��G���D]�[���aa������^�X��D���j��ڋ�n,d⯣�ے���m�cD�7`D�v�t��s<���<�+�i)e� 1�HI�c�+�=[S�/l�Kd6��O�#���i�Y�˹t_��8d�t1yZw�HH�M|�1��<��勗}��b�:��%�krwU�R�!»i�]l��`�_�~��{d�3��Y�r�X����%%;��V�?�~�d�`x��5s����!�yX�x)��pX8�Ǟ7IV�l�����W���=���Iz��,�xU�b��1�����?=��?�{>X��o�9�6k<���l�!�~�����ڂ�",SM�;U��p�Yz���W�mW�_�����wc($|˽d+@��	#��08�]��DD+���|��
3i%�c�W�L�'+�T�l5����ub���~��;W�u��ihR�%@��e�c��#���5���:�����D�C��?�+�K�Eh�#�@�%�H�RȚ����K?=�`�ã�����	�7�i�� 1P������k����\�����IV���w�D�~=,b�u��C�I�wbE�q�󽞅u\���Dԝ�?��	�N�����l�&r�K�Hl�E>�"�Z�	��b�r6y �= lK��
��r:��vmn9J~�+R�3_I��k�a�O�zOeX�������� ����6��>���29.:{sR����Wp)��W��h���@=~��Mһ�V���,��`2h�"�����s��q9g�%�|�{��e������e�n�yl9�qV�4�v2��V�� ���L��{,�,U�ˠ�ӣL3�2�[�x|xt��N�1�� z�@�n1ϑB&���Е8����xa�%*#�$(�J-oi�]��n9��ۖ,�r$M�hcG�(�TŲ������Hg�� �nז�mNF�N�k��#��$_�τk�U<���n8��kةd×�p$i��brf��Wr���(�n��N
��{�lY�6T@7��5ukuZ�y�ۍt�+�e1��y�7jIB,"_)��<ՠQ�Ҝ�l$��:1����9�˂؆o�Z��c�.}�`�qyz���@,80G��p��YWC��L�m��(�6L�f��%�;;��]�	g�v:'��g�����̚�F�+�� �K��4�6� X����0|�:`�-_�Y=Ί?�S�Uªȣ�waWQ��D}�c�S��X|6�#5G!&��������-�����E��6�L��~�4<��Ɍ�J��np�q-~j��x���<龍v�ͦ�7~]���VQ�<a�{��V~�K����$î�_�'��+w����t�]l*$b���)��xl����b�ܩ����*h;���*��(1�s�L�L7W^�&�{^$��������O���߃h	�7P'�+$�{��ܱ���)��e!�x;��X]��ǜ�h{wv'o�X-�Z�ro����fM�h�:��Ȝ��%�b�f�|i�<��<�O�b�=��~{���2N�C�G�w����O؀'�c���P??��)�������}�!�A�4qފ�&(�����bf�ח�禘 H���䲥Jj��M`ߩ^�>�_�w�\�^4zy4(���=�@!;�Q�ɫ�aV�u[q]��E~��)�-R����`�ӊ����(�y���r�B�Q��ݧ��-�t�T�3U�(�Vy���ĲkC�b��P��ݲ�"П�G"a!��@�'+3�'d''>����D���3�l����բP� m�UW�q;J��?�⼼�*�<Ng���%�T�������8���9v�)�9�~�#�V>V��9���.KRc3<w;�l��f�����O&�`Z_�*��Psr�V$��.�X����R>�aH�W��6uv�e%�Tlo��]OM��"`P��%JBm�U0�E�đ�@63 �ұ�V:����lU��l��)��h"x(����R�<��2��n��<?�{� wл��f�X(HgY j������� �Y��O��N�b��pǠ0U�1�fg�/`�B��@�":�EشYNYg�A�w��e�6�;s�	�k��M����"s}=`�XQ���ٔ<mj�v���]���g�G�����]�w�P1�j}[���XQ��w[gJQ����#�e�fnp�������s��h��ǌ�@�a�^<�6C�7�ma�zd�N���pn��9���S���W���ue���wK��:�1apz��G�Jc����-: ]/ݧ���>��7���\8',V̔��
���D��D����Xo ��-�����p��r��3e���7i�sm6�31-T����:0�}���*<���jj���4F�w��gw ��-��lH	�����w�K�f���m�^#aK.�-����1pHCz4~2r�Ex��j"_��
 �gOT�^�&�Q�\-6� ��vGUd,BVS��k���Go�)ŗg	jQ�t D�0eY�;ȳ�Gn=���R9Nƴ΀��G
�yz'dF?}��R��A�a�J;��з�������'��ɥi�Y(����4����G i�pP��/�;"6�&U�qx�{X˔���uR�0�m7q#�z��>�ɜD��T&����ɜ���c���7?�����ˣ̡�"�&N���E!tq$ت���.��`����@'`ڻb!K�/o>�Y���]��o�~��R:��`@u�]�e�(��U��JRn?[>��@�yW0�#	� 3�p�C��6G����ٺ���`���s���6�_q�*�BB(�+���c�"���G��3�ޣG?$N���ҥ�����=��~- _/�X�7bU~��y=\EA����^��Tdf��3r�K���|�l�~w�U�<7\���}��o_A7O��r}ޱ�[>���c����-iљ\��M������/g�F����-*�eO��X7!7�II+YfbE�~�$F߹t�̢͔�=�D)��U�k�0�ˍ��~��h� Gv�����g��V	�8�e�}De���n����z�%׆@�ӯ^AZ[���19��.��O�#{K�U��1\w̿��nj>��2I���X��:��!�oʌLZ����a��&�M�'`���;��D�ٽ� �Vw�n,��Ԓz\��;���)�{A����6S��GSJ���[�0qᅖ+|�!�ۿ�%���b���\��!;�'k���972[z��u��a*��bL
�l�W��ΊQ���򣕑�H�n~�>�Ѹ��%�YI$��.������h�<�?�orD|+���CMF�."���۶G����jt\� �Y��X ��?2�9iȕ[�Qy����)�;(�eq��h����ujKí	�.,Po_d�c8x���l�5L���*qN�oR�@����um�`B��$g����@5���w��,�A�S�=:o�@<��5􅯪��`�g�pS'��ܺ��>��?�:�!��#���$�P����(B�Gg^��_�l�j|��,5pjr-�������F(�`:_�<��PZ#~FUL�p���N�Щ�\4��Ae��^_,��2fϑ|�I^@���N?��Kđ�#5���V����.b�S��qa���oe	��;ܧ��+ݥ�1�ǁMrZ�YyIԼ*Y4,�s�M�����W��~'�vt�������`VE#�6VG�t�!�m�|�l�ˁ�Y��J֩�gp=�ߚ�$N���k(�+-�3.�Ɛ�Hb���Rd��1����$�uJ��"�؉��T�j�I��7��J?��OD@������{���T�<�5�64�n-'�PUd|���G,�½�;7{j�J�������Qb<�$�g��	KR���<qǺQ�0*w%�b���5�	W&�!���z T�dtɆc@}��#����umO�#�w^1Ƅ��x3��f	ɑ� ���r�*�G?hE5�Ñ��	���X~m��S��Q���ˢ߃���n��f�"1W��u@Hyw6��.�D�vZ�Ȭy׎'�9>Ϡ�o�s	^V�w?�H8�k�ҫs��IӠFT��j��?Ei�7�J��$�{�퟈����iQ(��V��?(�M(-$�)���{�Ğ�ݧ��	���6~���� ֓>��̺��*E	�M���6x�ڡ���b�-N	�?�z;/^@\��+�������V/��s���:�����P���VUg��A%�JH��\x�
/�F4[�ɾd}���^����^�wh����I'ؒ8���]ңf�1���X����upc �T	�d6�ۂ��~��k�:���$�G�aj�<�&�K�7�����o�s9��y��k��V����8��+ϖ_;ːM��z�W>�(�KI�.����ЊԴi>#S͏��K��F�f�k�C�����l{x�����>��,��vU�x�ʠ$�Q�D�ڱ��`/뷿�3r� ?�
e5�����S�;��x�����Z ����/�v-4��)'ut�S�����1�죋l��Nq��*=�`��!�Kq�����D̚�H&�g�����-�7 M�m齻�9��R�V����u�S����wT.���&wX:���W5�I�
��~�C�[*������!�����"�
�����������������~�:��44���<b�.;�uR��Å�5�l̈́���i6¹�!4� �A�9ߊC/nz-�^��H���=?�nTLf ��G�F�a��b�?�B:z�sy�m���,ʒ5�������<��?��{g�J��`:��:��R�=����q�{�]�����4��kX�W��t�� &X�ie���98���S�ʺb��ȥ8"�sxd�����Ԗ5y(�"�
�-�]34���^/���n���I,��v:
�aӏ�0#`3F(%��ޑ�ҒE:'�@�[�J��PB�B�&�676��u����Hz@�S�1ڋWT�f �t<]��$![�1o;� �G6���S�?l_�����p`sHB����.��������$��W"\+8=�ϟ�t^m�צ	-����	��ؐ-#6W�[ҔAV
�2���%���E�cB{o����v�b���ҍ�lo��]� :v�7i��LZ8L�p�5
�\=��l
|��4��qޣRwT�s�W�S�5'����tC�}��k�e��%�N8��4���H�%�h�IA<RC�� �8�Ai�S�QqTޣg�PPN�k[C�]O��P3��|��m�SEO��u��%��W�yj�PM��7��
)Թ>����k/���α�ĉ��ô6*����x�hO0��1�h���cPc�>�g�OSY������Lvq��R�.p�ӯ�R|N�@P�MV�QT��(��ɍn|Su�U���,H�9���>�(U��r�-x��#��0H��kzoX���	t@������f���Yr:>-s7�&F��%��gda�},�y[}	=�+�3�d��� 9?���ΆM����@�������rд���g�A��ef�b0����'_����TF�u'=�3�fe\��*�|>t.���
��/h����n�����	.���\ecB@��#��
b��]�G�q�Y2�u�m����Ϯ�1�$R�X2����j�T�v�L���mt�	�Y$¤�ۼ�l�%�D��اg11 ��������jThn����7t���qN�c��ך-FKȟuUH7����~\�|4l�nk�櫯�E����p[.P�[���.:-�4HY��:��BW�o��� ��i��L�؀^���	���"������aQ��4���I��d.�z���TVf�Ry�b��̌�I��֖n���&�mY�L���ӑ�6�!��J=W��__uu�qAk�v_�vTװ�H �����#�<r4"��<!N���pH&&�� cI�]l��0�.A�@[�/�$K����$5U6��Gyi������ɤC�I�I�J�� 1�f*cW�̦�/�B���MVgO�Qp��d!UE���%�4��2Gw�y�!��gi���x��~�K���)8
R���;<���ϝ5o�Ń��T�%�5%خkQ\�ڮYSg����Ұ|yÚ�$���nQr	��f�	�4�C�C}A|�"��UN*��6K��:����Ty>�?M#�up�^�,&�;'B7#�qqd�����7�}�62 ����])��w���߲�/O�;��V�m�m}T���,����@QQ�*��a��8B����I)!��K+��������;z8�o�����d�ۑ��~��e����_r�:��޿4�����<�}*�S�2��֧l��°�	>��� ��X��u�{8��]��LLF̝�p^$��o ��Q�<�rm|��BrT���!�y�B������*�%�����k֋�GM@O�� �|1.��Tq�m����&Ms��������:	�k����w�A���h�L�����d`s�JZ>cWH��Z����	��9$ІB鰖;k��	��`a�r�iSf���>�ɨ�Zx��=��BYD�;h%�N�i�߷q�~5�V_*�������B��K͗�[����i�h�l�ߙA9u�G������Df����
��D 14�q�Xa�����<ާrm�(<W��!:�=�0XĈK�L�cR����j�/�\Ι���^�i���P�^���#�I�ǠT~2`)�44�A���ھL����VW�/0�B6���~=�V�