��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VYkM�#j>clM|�a�pJ��p����*��>Q�	q_�A�C��@1�'֨��
[�xH���� �/�BJ?l3�����c��S�U�˃w��F�[���;h��j3�,+fG�oL�a��D,r�d�Be50�8rz�s;������!X�O`{�(�?fMQ�B]�*�%a����/�)+�"���_X�My�7�Z��6)CEW2��8�^`�y�EE}�%�w4���0J�!$sSod(}��շ�?CL����G���'�d�Yớ;ۘuC���M�$+��@7<{�6f�7W�8F12��9y�R�*�� ^���Խl�{s6���J�38��P`[zj�z��i�� n]�:��S��&�}��C�NA�`���=�ڍg�U}g�V�C	�
�V�P�-�����NX)�X�{����u�_��,��|�`�JRNi}�i;��u�uM�lO��R����w9����7OWiː�=L�>�������QyLL{:�	2J:����8�
D����I����#ԁ;B�0}�6��|�S�M��jl�4�u�/���2Z4��Hԯ\3�����Y��%�����3�l//��g��7f�]?�\���6��Q��$�����z�2�.��#����R���\Yx~:��*�²�? H����wp{�XʆsӤ�\F��ֶ%B��7!��j��SЍ!i��t0a�� �@���7��㐂�x��rO�j\��)��L�A�Ȕ[L"X_ 8`��4�c��G���!�w)@��
�ÛầFIx'�({�(4��fٓ니y%�1v�
D���S�P�}L܆�"'��77@��~�S�7��yy[[��)�ڭ�r���Q�����C��0�4R[-"��	E,"xaz�cGyOUXPKGB��-��ƅ}$� �Ӵvdj�1��=~$�i,ȡzo�7�Fo��]�p�V]It>!N����ƜC��'*�o g����	��IJ���sddǡ^��8�Ӭf�)�\a��#�P�K�-�缂�6�N�-W8��"�}�Ǝ
r��^�i�a �M�$�x��~��fcf;�җ�E;��i�;i�K$}�1��J͞ �"�4�?�Ii�ԬsqF���]�^OQ�]ص��'�ݷ��k�no4M�_
�Z�.v)�tٲB8�nf��.�_(ܱ�of�$�+&����S��[Rt���&��%��Zk�/�R��>w��\��""��2U����W�}�O�E9�u؛l�ЖP���3(D�Z���'�������S���si��Љ��ϲ�iq\]�#UP,��6�"�Ȓ�"'tiR!ߺ�����K����_k��*�o�Po�K-��˻�?g��!�G�(x����6|�[fd�o{8'�Ԇ]�!_xǹj�+�<%�t6�b��<$
��֩-!�f*&�Y*�gx�Ś��gp�Z����b�!0��mh�&d�~YyC
>���V��<|��#nx	�B5�m�����1^R9A�~���x���Ý�;G��+����$�n��YJ����zB�*D�)� 7�d���6G��s���pnT��|� K��'��[݂�w�dp(���3 O�j����`�@L��2��8l�Ë�Z��^����qZA�@�	>[����4)�C�g[a���$u��G����?�JI��Jg����.
�:q��snS�jv�X�&r�Ѯ���ĽrG�o�� 7l�&�ds�Il�8y�|���uȻ����"K:Y��G�.cv>��),uJh�����kye��jnB�V��gr�Lދ=�$�M@ �F�u:�{���*7���V!G\�p�0dIK��#,P G&!I�w�jcb�{�m�+n��űA���k"�T����8\���b-��B\t�/�XPt+�n�0.{�$�Q�A��	��LjpW�u��˅)E��7�GS�"ލ��ۅW�P����uf�kb�zq@�0�	=�� !:"q8���*�j��¿�u�q�EW�]�ѷ���D�L��oJ}賨V�0��@������6."��^}��X���ȑTF���7K�v��l×�#���}����>���^�"�Qz�s����H���aq�%Q`.�?#ť���Ow��Δ3r�,p���u+��r܂�b�XT���W����\y�NxԊ� �����\mJ]/�_u5���4��S��yhk �lka�@���xY���TI�ˆ2��,0����x�v�g�E�0�D�����M�`��,_9�Տ��@L�I((�@�z���۝�+5�B��C��)K	��鲏=�� ;�IUͤG�f :�H@~>t����?������F�c�ƽ� S�mV�3�I�kNt�˰���l-��
����:T|���p����vF|�h���1s���?�j�`LԳ;J���`7̍(jsK���v{����j-��e_�If�[(�ٗ2^T�<��O����1�梣¾v�(�:���X�9�!k��H�Ct�Ya���V��| �q�$h��ʶz���KQ�5�2�*Y>]�N��C�۞�:�^������I�iS����l���?R�&Q���*'�	�?!���[6��qJZC��w��MR)�2�k�3��G Z�}(3.�E����z0��GS,�<����>b��ͅ�,䘺J} ��M�:k!N.��QYߴ��CH��V��6��'ͪ�=��XI�b��m��e���\�Ug�*���w��2�-�yL�!�
պ	���[�w��>�S�kKJ�e�������������Zn=QS�� ��F¡�A���p��8�]�	�t]���w�i��QW�-�F@��~gZ�4M��⇱^:�<�rd�2Ŧp�U�#�\�*偹I�}=�y��Qó��h7��ml�WP*7>y�H�ʛ�J�Έƒ�jh*S(�5�0��R��8r�g}��C��v���,����0���}M�-Bo{"�����ݠc�b�M��nY�<q=dd ��69�Q�:�P��C!#H}� ��M��+���t�j��
T>�3Oz�����;�\�Fhǯ�s�rC"e:�Cq�!��<a�3đ�/�'������j�.-s�5�N�D`��n[���P���~M%�!����L|a	~Iܢ;[Yχ�#�W��`l'��X��ݸ��,�2"�W�A0R#��Z�Qr�G��qI�Cp۱< �|�Q�B6�!�SǱ� F�k�8�����&4�J�;�Nׁ���;�lD�Z��woh`	$��x����:P݀y��O;"��V�]w�Y߈�Ϝ�4q����4^%z��h��&.�2 ۝ɻL���, ae��~O���'�b��4%Cd3���H5�?���*�I~K��/��&���G��΄"5L)�0�݀����%f�*Y��÷�K�qKEA��h��6+�N
�1��@<�e�I������ujō�%5�?�Ih7�Y�ڷ���s�+�6S��Ƴ�.�����3~��LǸ��)7�)����c�U߲���H��q�6��y��B��R#�)�č�;YT �/Kt8@+*��<C�����U{2��%GU���{w>���ON9��e���ob��IR��M���èM�ޥ�o�E��c��Ȁ�A���q[��X�y��YZ#��j��ƕ�IP%�tօ`q�6L	�	ER>��%� �Ô}|��VL>�Я�7h�H5��"�w�5[<��w���x�]���e''����M�Q�A@�x��lb��=7�~�Fh>����7���T�G{��E=/�V�u3��+�
Ƿ���9�n�ԣ'��U�,��{eu��Ft|�^�T�q�v\?���X�-�+V#+��lq�%���B1�s�H�z>�.σy�tL�
���z";�C�K�WvB�xͼ�'|������Ǉ��/>G�"�txЭ��Q>�i{(���}1�p�CX9����t��a�d'!���C^�r�����һL�b'��2z&Z�1Yꐶ��9wm�郀;ۀTC�3��K�B��+L��)z4"�J�)8�=x�y'��8��Q���o=�e��� T%����[*o�-��Bo2�f�e"84�����8#�F6�P�v��3��-��h���as�|i8�����v�(�y�3О�#e?A:�W��ls�ɋ��v�*綾q����W�M�r�� u�8�س��BE��$G��?��f�����s�yD6~N�x��R}�&,d��ҧ�h�fIh�{�r!K)j@ߖ�ߏ�'/L�./�8&�ļ�E�D��˪�1*3d���?B�37ġ��a��-��7)��[�'ei������3EL�5a���
�G�Q� �/�j�W�
3��d!-��m���4ycѰ_iY�3�
�F�����~?ik	����^�H��KἬ�f,��TiYu e(0)�rs�X�p�R��}�������hk��.ּ�A���	��|�{J�l��,Z��Ź�{ࡅW%�3�/:`� 1���Ȝ\!T�
��T!8-X���aJLM|ߍ:Dk?�nƐ3��]0�#�ysM� �����й�ݹ�^�s��~�v��7����
�\=U�R�P�i���K:?kX�4���˽�=wo�EfO�N�X^n��G���=��T�"ݨL���+�ݞ˞Xh�ㄧa�jw>)�.P�;u,�ߞ�ʌ�k����;�!�e�*����n.�� to�K�Oџ��)��h*H�)>��[F�4^�>�A��x��x�#H��%�����2߉K�/����N���$&}�0R	��������N�+���m��ӸCFswjHL��Hδ���vN
�^?���}�����~�Aʕ��s�'kx5�C� ���^WFPu�Az�pw��>baǯ<���I�~��ل��z���q94���r�D�d�1^g����u)��D2�Qbʷ�$2�~�t�Z�[�o~j9"�����n�-T���i�P#vo��?�����َ�!{�,{m~?ד�U6�.�L���^�7IsR�����u<g���U�D�mEP�IB2�i�֦ъ�zE*�z`(��e6$M�i�Բ�<�Do��g�PB��z����߉��o��G���,�W�ޞ�~���ͣ7Q�9��ŏ���<C��6��v�R���ͭ<
12��gP9�"����oQ�:��� W��6��.r�%tJ�i?�6�#l���c�!-�y��8���s��p>D}��a�ntN���
3%e)��<���.�Sφ�ˤ�az6�7�y{`�j9tʁ�B�Fᡤ�s��%j�TGq*j�ߢ3*|@�7]�?̬.�%}��Z�wvXB�nU��!�X �2��ip��/$[%c�Nu�BV�׽��Jf�]@7a�ur�!����nh�NOg{���+H(����[����H��@f_��+�8*�\�P���)S�yVu�Pj�:ّzv�q���F�|��t|����3U����0Re�� ���ol�0op� $�7�G{;e_��7�hu"2��^�-�.�7�-�>�4��ii���՟��e�����DVc��o+�
&lè�E���������BN�5��a�}%5X��O��{��~����\a�l�#?��	���ܱ�4@���Ri���7p���b��d�xU����:��E��)k�m�40�CZA�쮄�;U}�Ok����P[���c(;�C�ei��36����lэY
�[|�}�{z� y�x"�eJQ�	�L�w�+�#zÄ]��=�D����Br�tH�o��j?��|�lv�4� �!qK�gxu�����F�b?\z=L`o�_�3[�>�7��@І�}�����B\.�3���{��j����g����<� ��02���W���,�ݖ-������&c�n�xk����W��.�|���s`�!���<���ϚU�s0�e���5ϠQ^D�O�ԍ`Y++�BE� E�d.���ZV���\��
����O���*B7C�!E�(���S��~N�����cD?���\�W�����-�V��Kn�QTe�_�q��\���ꉌ�l
=`>�غ�=!~��ctH�(�1"4T� ��&Xa�Y'>�ktY8��B�N�ޛc����9�9�y+�G��=h�`s�*�i*�S����$H,c�D�	=��
j���^�\��䡩�d���9�e��T�>�u��<��w��3Ʃف�@�U�WÿO�}K��G��sJH�}�*��
E�gVΌ�5�Y�z���\��(:e6k���u�:ݑc��B\��/>>{���7ډ����/�/��'�G�Lʃmۉm�����ǎ�/3�Q��?".�Y��t~%X0ըq�Ͳ�P���v�E�`��U��2@��f%�W�.�=鋑(8��R��� 2��duo�7F�W����!�h5.uo� �l{F*��Mԏ��G2�9���n�2�g1��vn�d}��}"�*JU���-�4c?�x&m��?7,n�q��c�"��^vܰQi֍�����ֶ�|xPڗ��?v�:~��=�d��U�����|��%~�Rۢ�gj��_Ib�@-�;z���
��M�ۊ�F�NWR�k0�"�x���(�9dm�����&��.d�e9�7�Fώ�M^�bj�����A}�n^i��{��(���]rL�����q����I���,�N>�-w@�9�]��ƞY(L��"P-�C�3�Yk�̰Q�Ϥ�-?�Sذ�s�+9?��^�m�nK�Ur�?���r���k�F4���Ҭ��tVP��'� �
�i�k2�
���_t?�)�r#*Z�}U�3(2�+�_檒��-��-�B:��PT$���:�"6���D��4l�+~qCu>���> LUZ�J�n2��_�$��8<]��V�t���V��2 �O�w� <R�+��:S��������v �J��T?��O��X�)��)�ҹ�6��5�&_�4�tAaN3;YȚx�P�	�-�ب�f���w4k׎b�J){�̉�|������G�a�5�����MI�up�`���7��A�FQ�8(�6�\�p�9� O]�l� _Le)�R``�~�jOe
>��?�����ly�>�T7����98�a��̸�<&�9ux���E�6�>%duE�"���)�X'{n1��ӥ�t�l� �\v<?3��2���(xA�`t��onȚ�\z�O��m�
���дX�N7Mq�2�o���5���Qd��,X����\-��R*s^�#��<��Q�K5`�L'��g�C��.�>
��z���ehC��BΘ���0 ����LQ9��fG�T7/�oO8��Q�� \�]&}�U:��s@x�c^�Q!B�~�,���5������Md�~��	A��~m���/�OI�?�:��6���nnsa(m�oK�^���|l�G-��">��A���W����>�5���~��#�l稴�I�!X͂<1�~-����@ c���m�����.�6V���d��S��{����ͻ�޻�-Ď���`��L��G:͜�F�}5*9,���Es�x��8J ���zڧm�)�m l�?�|t��a��=ݗx1z�D�A�,^H����1x0�F����.� ��_Ў�NU��"���=�O��:�o����X��z�m���f�1�R�'y_Մi[��s�8O�S�RySn�=%�r��rj��Lx���{��!1���6?�K�!{�}��]#������:�A���w�l�:Jk0'�&~���bNy���w��)a��-�$N/���
V�z��Oa���,���P�S��0���47��u�};�M]�9m��ݳ��du$�-�[��P��J#���w�u7x�8���3Jx�PzF�sj8T�������	<���ei=�����Pc�@:<hg͙�c����L�!Y䂋��JQ܇w�V!}���ˀo4v;�"�R#p$M����+��C:���L7���~rk)�>1��\��a2M9,x�.�Nm�#���H�����eoNт�rDQ��'eϕy�ÆW#�-A�x/z~LdQ6O-�'/z^"�i���!x�#]��W���ؿ��*���GFMx�?����Ѵ�CZ�TGq�\��]b�6v�4�kOJ�����NG:5%��#�@=�w(�x�Pf�W������,�.�&��I�ol~q9�����bd���3��q�	��d5��'�P�/�.ID��e��
��4wї���W���($�\B�ǚ�c�D$ď�F��@�k�}�[��7E���<�����: ��+7�+���&'I�8Ԑ~�;hU����N�)MN�&���p�D7��u6�K�`���9}V�
T�~���,�mrJ�h�-f��2| �����/z�������s/����|�9�+L��<<p)��?n3���9lʫ�ɚ\�w������$[���;���-/fS� �SJ�~�nx�e1?��I@�
����vz8jS�P�x ��8������R�z53�c�Ѓ�"},?J��q
Y���c:��4�u���vB��*���N��GnRV��r
�B�����y��%��@��ML]!71n�Xp�ͱ��sԗm�0���j�]�y�����w�@^�ٷc������߹�b%xʡ���r�1F�$ql��)Ō�����>��m�>�ɫ ^�d�)Gbl�"�4���2� ��O<)Q��=�z��Ã8$���.���PG@{	n 1J�1H�
�i�0��y��n��}xlJ�G�Ģ�	����L2/tˆ%����g��o5Ve�f&����|4L���d6R�X򞹕YLr�|�K�K;$��Ժg��9����@���e�O��8��h�v�i�A��:���YJ շ�Gϧ���G����B���)�j>9_s�`�V��vZ5�L�+v���F/���MR-.����I�!��VoG M�t�$~���:���IS�I��(*j�p���=���v:�֗���ɣ������{ ���>_M�N��DP�K/w`2y���N��"�������7z�l	�5zw&��N���b���u-�A����i�JK�����S(M�nd� 
kj�N���K��.��>y��{���T�������P����!DI�o6��r�u{[fz����RA�p�������	�LC5@�H�vH�B����)L@���{�v>m6n�:I�]?��ک��� ��rH�Ր�ƹ�b1��R���;d=����y_uo�P������K%�5����&�]��dmnI���Jg)�?[�.��2�'K�y�DIn�C�|�o���ٝť�E�:����1���j�|�샰w��������#�p�jY�>�v0��I�JZ_��$�Fyε�	��V4a�CN�����&B����Ej�/(���O�xΆ�3:�4���3"t
�Nҝ���)���3yY2Ń���W,ߪhjM��(�L�/�U�`WA/J� �p�u�.�p*r�q��������A٥	����'�8[������� �F��v�������Bx�S�U�`S�Å�o.�Bl�j�f�ŭ�~,����<��0ͣ��hyg���: �X�!��6<�I�b�H]MP�	?L�T5w����E�s�PG�� ����d���˘�Y�\`ltqm�;���>��7؁�%�"q��:�ZI�C5���)ߥ�OO3��sE��k�f���wB�*U�t�vd�y�\�tb؛'A���P@�XW�����������F���{ӨJ<�?LTSi�E�������<��:;]�%��\�H0!t�"�j���Bq0U�E��e�-���z�"F[9�'��Q�
�Wg�ե��f��� ���e:V2��NKWO�[��j��(+Y�sn<;�,�S3�:©�������2K2�'��8vg�����'���k��Яi̿EQ9�O����z���.1�{`ĳ�~��x���'c�ڱ:*0�x:��KF�	z�`��^ U�c���"`(1�ZV1���o�AЉU��(�c/����t�j��A�f�!��Լ1���řTG.���|u�3��%�6ZC�uzb�h�n1�tP�v����+,��D��J��v}�;؃�A�3L�+8E=���(l[��WoU$+7�Μ����/U���o:�d�9��͎�
�ʝʰ5�7��ҞW2�[c$�}2UE�/�Z��:8�t���S+ص��m��O��z%@l�N�~[���dn��@.���ʆf1�(N�6����Y7h��:�#EsK!���d�S�6;���W�nﮥH��;CH��/�rv9�.G/ ^I��YXs�0%� ���s���"h�)3�8���Es#��	4;딣������Q O��A�63}�H����;����}�N�g�� ��y#|
��}{�o:\=$���^�K%�������2a�vQg�J|
�����ͨ�$�� m6�y��7o��H�`�3��Js_/9eo��g��L�I�pɶ���*+���E�2�fä�D#�
�����z��*�C�}̳�]�k�~Χ��r0 `Z����W͝�h*6�s��v���aӈ
�9 �~�HG��нh�ƨ7�m�jp!'O�.0���}�̢u����.c}&'�Ab���U)�\	�P�92����P4qY�����qM�3���\%��+�2	�t\�@
q��>Bl��-&@��a;iŵ����TMv��ήHz.H���YrP�����.�q:��"~is��`���`�:�d���%55"�\0}A<煿x�!UoCNMQ�ia96�F�%u2�βF���3S �qK䣰�4���v�2d��K��;�ӰĬ��"����W��s폤cD�7a��m��)��W���v�>�&��=.W�Hi��k�p�w(X�G!C%9��8�7,`Sk��?Gzv���j�X���7�H�].�I�XM`��U��=BL4�V��٩�y9��w��c+R��;-_����!r�ü+z�-q�HR%k�NI���E��kA������c$n6�����������imH�=�D��O�3�O�"dF7��ܽ���ߺ�I5�.j.�Z�11'�zvT/F��0��R��y[f��dqu�J����hbi��.k��	[ǧ)K��Z��p������j�0lP��mi�kD.D���?k#�N}L�2����x���@"<}3"4��=|i���Ui��)l�=�zj�]�^���A���TH�h_����ce�3�|�uq�S?[�dԍ�t�f�:�^E�v���/���`���Bi��h�}��/*F�B7�V�+�n�& ���x}�Ó�ؤ?q_�]zb���Ȁ��]��0���s�?#�'u����$�W6秪�W���o"�R!MOe�d���e(�f�%���0��F����7g���z�G�'ܰ-h��M��qc��bH�����Z�,p&�]��G�m�KNI�~�)oHɾ2ۆ%����$����f�D	��y	���3�iF����*��Xߧ	ƈ�>�b�V�v��y��+�?��5�����\�P/n�����>]^_M������'"�D</}6���d*�+h���t�z ������VP}g��,�קI�G-�nHj�-�ƿWbQ��b9!m�H,eh�xR&�,<��s��z�����՟R��)�3XW�x��+.�oAC:��H����k�_<���=�2
D����aa�I�^r�k���^�X���@�"���v_�w,JAY�@�@���]^g�3}�� �?╍�'P_ ��n�l�$�����Ǥ�8uSި ��Y���O�QHm4���/��T�C`��2��3�]l���n�]�ʹh��	���p
W�C��3�����Q9�������;�
��(�|szL+��V��=�D�?ֲT�ꄰ���q����*�KG���Iu��Gg/|��e𮄬�>��.J+?������Jp9�P�����T�ͧ�����+NF���������������@�(@�N�9|�M9��b���cb�]�H��W�U� �`�/I�'v*b��__����y�ѹ��ŭPL<��p�b�R�L���dT���f������-6O�¸}��Y[����읅��m�v5v>�ﾲ*����[�m�/�������$�?��d�5pa��[���tM�K܆�qbjn0�+��D'++��򈼻��m[����5J}�� 9���=�vZЫ��Kx�%�꣨]�{�N��wW�B�f9�,������<V(����y���S�����8Ɠ=��<�N��L�'fF9�}Y��p黈�v���|��;����ޒ���1�7��7��+A�m/������@
ʇ)�����:��.qw���}��<|���B�r���5��Kb,E�gE�IL�(Ţ���_��e{�p~C2���N���V�Y_�_�x��4�zAQ�����d���Ts���o#yN�q�̨��z>�u�&im�5|�*�����WB��"��i�Y�Ϭ'AF���&�)��0	�$é�l���{��|(	�B��u3Q��i�)M\���	Te��L����tV�U�M�O�Z�vn�&x����<��4��a�K�w���F�k�!Q [!��ʔ0T��a�9��l�q��*���V��¶�>�!�7������S[&���K�D����2؋9>K��wa�)|*�K܈p�򶩨]�t�<nKFB�ahq9zy5��<���M�+"�04�����ln�U���>��#�T����g���������wu��r�S�ͳ^�yV�����jY�ޚ�S(=h����ٶc��[1�9^2D��`�&א����;+EJ�5:�Q�
|����A=�ӳ_u��94�N\�M�f(��5b�g�����fc˯jmbV�?G���oP��*?msGk�K(�=Z��u(:<�:�%�Z�rR4�y݇����|_���t�x������Leh�O (��W]Qd��e��)�[�Kߒ�1���cGp��[�C�5;ء9��Sz��X�-��bi�B
����V�?K�r�L����� �-аz�k�0��O��X�6�x�7Bg`�k^a�ܜCEF�<|uC�r�9uq�6Thj�<kO>��e�K�^뭐��ׇ�9�� ,d)S�ou����3�ҥU1���iȇ�:�A6Bɘ�>&M�̺���<�kQ"Ǜ��k)�ê���* ������l��&yt���Ẩ2O�Z��d�H���N���Q&�(CJ��L¼��C��2Ұ)�%(���l���Ac�AG��i�a���	���I 1]?K=?w( *�KG$�MmD���[Y)�{9<X���*E�K������M[ [E��3(��"�*w���'�����N�m �5싏�IH���#z$�<a4�%��J��چ���x�'�6�=�]	?7�Rʍ���IG�������p'��|�Q��Z
犢��Gɷ}q H*�3����(������回
ha#��>���&������^�2z��~"��'�q�_�°5ov��Y�U\�Y&5���5�TL��p�ϰ�.-�3�ߦ�?\�pK���<]��o�=g��h�=fF"Q�Q��˩�[�y!]ȝ��*\UE ϵ�P����H���U�Ń���Uq�O>�E7λ��N8Y&��x�$=����MII���'�)c1@xj�.>�Ck�:|���b�`٬����/����9ϙ���8`$S� �2�M�?�d�"��(7^NU8l�@k[�g��2�+��Ѐ��yu���
�F��i4&B��C�qm�����s+g���7ٵ���R9�0�5��h�^���yΆGņ���H�2�O�`�d<A��@���#�1G�%�mM,W�2)���2mz L'����2��H�q�'�����h׳I�XO�j�b.	��r*����ސQr�a���d��e��+��)\��
�]<�ف�BZb+�K}s>��ꐜrc����7 ,t�I3�vy��5�k��ͱ�vq��(P��x�n�2؇�'R�,��c�I��jN��Vr@ᤞE~�k�*݇���h��x�y���;��%/��0�C��2*S��:��!V�ڄ	��/��.h��F$��fAX#��R೷�e��L��-I�@]M�x���g˄�dgS�Γ�����]��� �'���(2N�!���L�"�M��E~	o��Q =�g=�w�M���;�?)X�3��_��ߵ[|r7��Q��9t���:��_>�00c�'��Q�&�*�Ťg/�T�N�JD��w@���61dL�\?�Ҟ����g���n�d��Ň�l���úv�e����`1�_�W��* Ƃ�U��3��b��}�YkB�1ql�"vC��%��ƙ'r��	M��� d����w5Q���;���� ���3�:9Pu��6���%X�^,��w�?;�)���mk�B����or��N-��
i���)��*�����\J�*�iu��9����^�6~��D�%$0�鐠ZVt)��TP�f�AѠ-C���Z٪ᘿ��Ѽ�$4��i�`���^�Ɛ�n3��ZlQ��_���.�ÁTC
yB��˄����j֥d�����	hI�Jb�����삶�� �I��m�D�Ndi�.?��Q��~�!��K楇��qQ_�2�k4\)b�7��ni�������/���Ί�r�<>6��o��8���K�D�d\{�Yu�	��-�}&f��1��Igz�D�_��+늙��{��@W��Ә*R��������S�
.�I���hs�0zh@<�߮�G��D��9��2����Se��o�Ȥ�M��v�^��f#;��� ���Y*A�@��J;�)�-AЏ	�y��%܉&�ZLv�i�&�F��xs%�r��$5�mC$TU�de(��U��ȩn�̳e�<w}SD� hUq��u���%����X��K�$LYi�d���-��-<]�Gcp)�4M,o�9��g�Y�����GƬ:�?��f��ȠO�Ւ�����.��,U��a;�y6�e�^�Ӌ]7"`�W��':W�Q�pX2��x����/�z^��'�2i+vb�>r[#�kL��g��VJ29��Y+]K���p�j�1�M@վF�+myÆ��#�R�6��$c#W>�vZ�,�Q� ���FLK�k4uMm'�V-����;�ѓ���i��r�`���:�DpYb��I����	y�LcF>��V�g�����f��j�N]w;Ij�U�s����8V-]�U���Ƞ�p��i�UAD�mՃ���u��������{%F����)�1`b)	���x��Y�);C�4��Go��@�b\N��	�R��ܟ�N�h@�]�~C�=ٽ���-�ɩ�88��r3�G���W?���~�lsSFJK�� �&��
�$�L����J7�D�'GB��#-M�� ٯ����&54"�m�!�p�m��D�sk�ϴy�f��^�����U1B�q彂��V��������U$�@���e�&��H�$��9լv�9K�ѭ���A������1;��疧$�ԕf��p�x�1Ffqt.�@����VRvS�M�7x��,Q��t�`T�n֬wM9�� ku�3������b]�;� �'�{��j���²��F�_�f�G_%��>3��?�]^�M(��^�78Oz�ࣸ������ �&Vw2TUu�߁�|�Ш]KHR��M��m��ՙ�&��9%&s�:+vʌUgz�5��C��"�� 6����2�T��־�E��pXR�	b@h
��낱�A�W����?�&[�bT��
F�ʀ�����+1KY����Q�ꈓ�����'�$�4Jp����Z�2����`8���QCs|��]�Y�wwsW��y{��' �gd��9ݩr�^{�Ңpy��Փs�l ���ڌ/��Vu�ȕ�Ɩv��̒ݜ�����i/��Z��NӾ#;h�pr��5'�0�����&22��nx<�7
�������gA-YCGO��aKbV#�%N2��Pv {[�:��8n�E?&aOQ�iْ��4�{�?��~��9y� MX�B4t��	�|�|�=������M���[pK��7��ڶ�jmڎeݷJ�����"��B��0�!�����f�*�[`xWy�Bp�ֱtQy�4������������ iG 3��������d���2�sUaƦK~�Y���P�U6�3A:4��s�Uᨃ�C���K)!j�o>�]m}�v��`A�7f�K�%�f4��/N�|]�K"�9���ܠn��n����ކ�����Y�7FbƉ��s���7\�`�p�nqC��6����[��MI�o�q�${�3�43�t`�c-�s���h��èx4�
�f@���)��b��T��r͚-�K�4�������/��2�90�����@Ff>中/�R�[\�o��z��TE>�����������E*��֋d��bނi*lz�+WCb��4|�_���������]��[�R����,PH/�[���ƫD&�1��"��/�YAӣ�ZM��fos@�xځPwe7�[�m(7��U*��DF_v�1'��*]����نrOv`��u�6	�:B-����i�-�	��	�n��r|�����4aW�2a��,���qM=��n����:-h�\	diȄu�-:�<`��6��'���#y7�>_�NYbD��a\򋐕&`_��.�22�٩������?��P��v{`��C�h�̿
S�{�$�nɵ���X,�����|g���8�������Z�iq��9���u�O������.C��Y�$TMű���u��^��1��aK�(Ÿ��.�:����.Va���Kz�1+�5	k��S�[�dE�߮��r�v	���a}m���mV�60�>�n:ܜ�`�;T�n�EM�3;O�M^�S�Tp�Q-t�K�=Û���ńї����]>N��Ꙓ�S��lJ����u<�c'r:�w�JL��)�,|��J�ٰ��m݌q�;oB�]�m�4a��O��4XB�=�bK#ċ�lv�)�����uwP�_�;s%k�ȭՅ�����56v�cQ����e{�b���~���׏���� U��5d����A��(x��4�W$���IR]zX�-��^�ʹe*�b� U��^3
:�ҧ���%�n����#0�v�y�L��0�Z3C�mG%����#�X��;Xr��_���>�a��Ѷ�;��hkY�|�@�GD�9n��{� ����(�=�9@&ݳljS���x�&`��"�������
���o�Wc�<i؄n�z�ğp*�vD��W�K>�nLYh��Y���#�����Zj恓Dw_�I���������Si1W�*/7D�^��I�Hv���w�� =����96,?P��cj/���M�I�q�i%��l RIs�I	���;ђr��6+�Li0'��S��X���!����C�_�t#���ف��_�S�����}��������)�~m�:����F	: �Řـ 6ׅ�Zw���޸��Sխa�sW��n�!Bh��)e��t���cڟ�ň\����ۈZ�U�O�D��.�!�2��Qߎ�RL�\����z n�ʌ�W/��	G��1�௾��&%\�]B��}I�!W���/�!�O� ��Z����6Z9�Y'gJ�%6����TK��B�f��TLm�{T[�7.�x�E���g���?Ŝ;�"4�t/f�N{�}�9u
�����Fi�f�!g�oy[~����w�ه)h�Ǟ�$�n=��W{�;Y�z�xT�N4�N�Τߏ(��Y��&V :�I�n>���1׮S���^3�8`�g���bwOZ<�Y���rD��GU�Kp��M�q�c�u��h9- �$1'_�\�3��x�Jb�MH�^���fҖ��%0�6�!�%g��Ko}���>�0�$��wi�l}�1�e��|3��G�:�^�'J����i�X�Rķ�h^�w�Α۫�r���{=Dq"Ǔx�����먧��$�aU��F~�u�B�A� D�=��u�TJy�"��"��a���x��aA7�W`���<@��+�/��%ʱ��Ec�>]���ͫ׶j�9?Gr�T(��w7�?ً;������3gG�+��M�(� ������I��_thv�M}�)���#�mW-�辶�U�\�]͆��N73����9���,T-� m��y$Y��z������!�X�r�D:�ٲ�Q�� �#�$��P��[Y�yN5�����'�/5_�BMՐ���f��c�G��5�b4
]H�|�W\���ސ�������5)�{s?��t�O~GA�}~g�Ά{hg�T�>Ԍ�yޢa�'���N�\{�����z�7*�$/��y�T�ǄDQ���Q���h�l�!���_��f����Y�[�IV�`���+��	��h�
�"#�g>��@Ց�[MC��uHxJ��*���] lr���q��m ��g^|/����G-E]Y�)yǒߧ�9�8�8,� 	{��`�E���M{'HA��j��.��ek����pպ�:�EܭZ�m�OT���������J��4
�9o��a��A�{'�_֍�eJ'��
�޹:�p{(���V�L<��͘��z�hz�'��A��J��S6=�Sq�t*�׎�?��y�]��<YR2��?)#V��M�UZ"�
�Ȳ2Ch��:6�ڐ���O�RD�{]e�I����d�tG��3[����,y���N�}�bR�n��K~�<���@�����'�m >���������<��|p@�k�����ћ0u�\�� ;=aF�21%*�@6X�:�l*�(��nG�
��ͷ�B�z�#끥��� <�����N��Y׌i!�U�F>�4r,��Xz��Y�n�0�W���W
��0]�d��`�=�U	�� �~J��j���@֭}����v�@�'���5W�(L���-ƌb܎4�o��<��o�)��N�ި0-I���Ы��q~9p��D$obl��k�A�Q�9���ɕ����G=i��{hp�o�@,�Ti�U0����t��� �ы�B3����|�l�&��#̥l@'��b�^!�*.8�ӎ��M`�;TO�g&��e�sL^J�����wd��g>�Xm3?
���L�D�i�1��G\��<���0�bB�uZm3�y�ݡm���	/�lc`&��Zp4�K�Z�|���d�;v�)�}�	������k���*�������|wi���i�jg+��>�`ٱ���'��ΗQ�pXO��S%9 �4
�^��e9`�����S'	�GU����h9=�/�U��-�^���{n7��q�J��F�\";Qocy���PA�0�"��ЕG�F�Q$���u���	%���缟�����Shxp���i^�C�7���̓��.�
\@ٰ��:�
*��Be��N���l �)�7��e4(` R�Є�
�k��l��?����[��'9�2���<���is�nH�`I�h�sq|���0EB���ϖ�������9Z9�k�k��b���rj�O����;N�:��Eﲔ��`mN�"�*��Z�)����\��%�}�ɓN��P�	P��3���1�Z:C�`=�%��l}~,)�~o6Px��\��Ƌ�݉�t�=�i�pg��"7��A��h����(��T�I�l��S�e�D��g
���2|p�}[/%&��ζ��-�<s���	s�ع��f�o�� :�O��c�B���E�oYC�-V<QD#��g���?k�J�����[�@9�STC%a�ҝ"r<w��A\O�#��K�%,��U�|���5"�l������LC.��(}�O�eJ]�]1I�,�C+�~���ƒ�V��9�9X��8^�<M�Ȼ.H���$G��v0hJ�l��um3�I{6JV�0�@%,B�GV�o�N��Pü��4d�-{�n-+k_9�/�L��@0gdVM$hY�k���^�o\45^g
b�8�[�0�`�>�tt{��A�o����|I���D��#�7���v\d�d��T��͢s�E�Ο�n>����`0���)�v�n�e#LuUrm�ź�K���=���a�B���v.�B�p��kߐr�/��!�@���
�j�:��o�j$�
Y��p����
���u�����>ۘ�W��e��4o�A�w�<���
��:�������
A�Ȓ�l���s"aV�q�E�� ��]*B�p��;բ�Ժ	�<�ft�ϧM�E뿈Dd07�qK#o�jB���$��1Bˌ�����������0�d���=s�a���E���c�@�h$x�\�Z��zŻ�����Mp�����<�:�^��@D���p��b�}d��]��^��J#'����z3d���|׷���%��|�Q��ģi,M��`Ѯ�f��i:����һ<��g������n�e���	��� T��C�l�G�������^:��Z0�%
"a���L���9k0'��U�,'��������9�:�8��Ni0�dT�)�**���_�G=�M�WW��t�/��}������C� �7����W��`�"@��ک�,�Pو�P�����S��W�3��:�Ls��U=�֌Q?�8��.��F;[`!��=�I�<ST��$�z�i4��=�J���{
���5zI(��D��M�8�]W���|��1�\�љ�I*�&H^:�o�9TwWe���H����#�R�Z��L��y�1�����'H�L���$G�a2��(�>�n_z/O���7
�}�k����~���.�Plm���Vm��3���mMu���=������D� ���� ���"
�N��	����c�aVy�E鲬o�ml���SԮ���^�Ko�y�|��<�Y����m@�6)E�����-��3
}/��>�,���6���.����bY�3�@�$ J���ܿV�c)�j�s�ĺJ����p�&�SfE�8�9)˂��.�=X2���|�����}!�RV**7�o�
���o�����e�K)�8'��o�n �@
��q���+�=]:ˁ�
��|(��X��;d]'�"�X�ֶL	,�$�'������&���=�Va��	O5��ސq��ͤ��|�P�$4B�P0ͅ0O��6�H�m�5��d?5����Q��Q�Սvb��I�j��S�?����U&Bԋ�V����v�&;��h����d�n *��[���c��)�@F?�!E�̀	��\'��gr��tĘ��y��׏�6�����EB3}y��,��B�����^�Y�_��[rU�)��Y�k=K�i�Őɥ_��������I(�Ϥs�U�r�ՅëW7��Јޥ�h�_�g��n�DhQqb$�u.X��Ĺm�xH=��[X0�OM�@�a����!�A�d7P �����NV�]��BuBx�.͢�êpm�rP�ڣE�(��K� 1��"ؼ4�m��AxG�k;�M����Ҏ�-Ӭ�sn��g�8���Ű��K.�����L�jנ]X]�d鳪��=��j�9ůa�ݜ)i�+��Z>���h��!�N��,����VK�
P���
%Pt!�i���@Pa'�Ȋ�e����W� i=�{��,�U'�����9�&Q3�TX�qp�ڟ�j��| ��e�`oB�#4Ջ����9
�S���Iv;(ܾ��؟})�#Y�_�$S.�k����Y��8��Z48^���85	����5���=�:�Wo��Ӫu�
����	�f�
K�틲�D��W:���������e��,rZĤ�0��qĽ�����]��i�kﰔ�L�33��� &l�:��H���&A�D��!Jj�,�܂�)�w��{kV4��5N�`TU$L$�3��]�U��3�x�Fw�K�U���k.�p��[��Y�سOLciϼ
Mke�p8�c[������	ͮ��*J����	�����i����>\]c�_��C��>�ˊ�췻p���g�8-�.;ƪ�Y�l� �JU0���_�$�x]�/����xyt�d�����*!�!����Ϫ*�l?�Ɂ�8F��Y]���/�^���3I��k���-H2�r���g�ul��)�����1K	�f�K�d`�0��5�GswM)T�I�t'x��>�:����n�.��Q[�b������A�;��!�v�^P	�C�z��/ ܅�H����N�v��>�HGǠe��UjO`��>-���>��Vx�1v
rx��!�a�?�`PEA+3+)�OB�5[��PkZ��7��[��?7�G�	����^�J�|�}[IVb�8K�C����j;��kF<�|��褃OOB�4��=����$���yrk��	i�9[?��X�}V�^jYN�N�Ѵf�.��p�m��fi&����4͆�S�C�u
�>��(�7�@b�OCh�� �k�P�v�+f � q'f�9p�J��:�;=?L�l%O$7����(i3�*BU��.ɽCT5�x��f�~k���u�����\/yT�☭,nx��ny��>�-�:���-ܟ�s������u���^zp�)m���:�NV�X$f��W��0�}�Ɓ�g.��z�&�KC|���.��\��M��Tu�\g���A���|<�b��X!P�`0�_�/S��.����{���9`% �j٣~���� )|��V�t���x��"����� ��FL-�����f�%�M����l*��e&��l*U��[���/��J�0 �|jĎ%���B�o?�E_��,�߄�%�sdy��I�! �*n�"�=: �M��	����������ZD�E���[E�A��g�B����B#9�>���|��OfCo���!m\B�J2��Y�#=�����
BDH<�R���Ϣ�<r]Oa��<X�j�������vNYR�鐐�+��?ߊ���Ft��vh��w�2�`�_Ҳ��@:
��� �{^����{������;��N�R��>�ێ��g�/�����|���ŀԸ��im#3�<�u$�S�7����,�^0���7<�����۪5ǎV�I�&�-�͈"��G���Nz����:�z}.�h��oW���p�+�J4��(��Vd���e��ʤ��bW@3�nM������H=kO@�?u�{8^-�����Uq��d����)"�m�5��X-$!�l����W�c�"U�.0ϹR���"w�sߡ�,�y�B	��@}Hͮ��z�3��<�5�⟏���n��iŸ�j^z��8�Z���E�P̙�b>O��Rkm�� `,Z��K@0�	�����؄��pr��0-.��w�!BAO6و�y��""S_^%ND8�	�I�/}��;rg&h΄�VZ��R*���u!�-4����w���v0.n��kn���96#� r��$�@�!ȩ*���c-���{qЃ�CP��me~J�\#��aI�Qa^t
�5p �̭�����ux��J��S\]�������:�J���N�u�b<��6��:M'�f��*���6}��]��PV���~�3uD@�{ZϾ�\��
_����pj�<@`�b�f����m�rv/���i���iyY��F;��ڀ��� Tw�}�Jx�a���9x�\�Ӛ�x��h&��oq�R̚���`6û$<vU~���0v.��D�+\��v6Կ���W|� �UF}�֘>�s��GwϨ�FzH;J����p:�T�����}�+�/��{1��C�	O�,��* '�M9�#v�5��:ް��T:��66<W8&���^+n,Ne�Ճ������Hg���r���aڢ���]��쫋�|� (I��4 ��=�v�/�ye��!�sT�g̜1Y�&�_���cK���s��چo��N�
�ot,*��y�K�Sd��Wᴣ �n�)Z�$HC�{�=��h��9��I\����@Q���В `��[`!�A0ܔ��]��^�4O������6Hb6������XK��}N����;�3�x�#��T���h^��Aza��Y�<>��/��:���A{0a��G����'̈́��ڪ�I�;k!�	�G�8��h�V����§��HK�����%!�Mˬ��>�BҴ�~dCl����\ � ê�[&3��f��#�����,�5�P	���~�[+�dLH�{�lu{R���G� ���-q����4��r����z5ba�&F<!ПzV�`
s�:Z��r��ߎ��C��������l4��2��kL�7��z�:�쾈��9�|xl�FxY��;���tAj��|�w&���h�,���UB>��b�.H�تSOO����s�4�w�b[��S<H˫��b���J���̢|Н��hu@��1��k�C`RY5K���`��n?�K�Ie���M]�	�)�A��Q����<����3J;�ˣ�r?��R�@��=��&Q%�@qn��&yL��8)֔�V�7�=*���w��[� 4}��(���4 m�����r�@~�r+3S��K��f�ƼҶ::0��6�oQ���e4y8�y���=��Yy%�ȅ ���$`m3ހ���y��	��ƨ��B�2ߛ*yv!?A�*[�/��	-<�Q��f�9=�����n�pS+�<�&7��z�ƒ>��I��
���;��]��%4���9}��wTԙ�������0.����]�?`S:3Pq:nێ}�ݞ"�0�e`Ż,��0l�^���٫#�z?��p�LsLZG�03Y�'gt"��ݦ�Y��(�P���l6q���%�ѷ�`y�ߵ�R&��Ŕ ͬr�4�Ƞ�4�hb�$��K���
0�B��dN:Y1va8|ٸ�+e��e,�PK�@����)�_��KNI 4r��]�r�d��׌��~�$Q��%�(`d��"}�;?ڦ�*�t%��;ha��[ǒ��DU?pJ����^���m�7'_�|l�H��o�
_C��d	��>"6|�3��q�.��1��7<�n��`h��%�����6l�)]>8u�aa���'|�V�M-M�o�w���!-.��x)@5�VS�@��Di�k̮z�۞%b
����Mؼ˸U�N��d2�Wt�%/X8�Wy:�,�f��= �pq4'utsi�=��6��+ؽ>�>�v(��oC�W��KS��ʦ�jˇcw�+����|�>����7���'B�+���"������",Zop7S������TQ#�0 +:�3P׃���%��ȡ*�i,��R��������*���P�m���N}��R���C?,HݷOb>�����B�w�a�<���~7Emߕ\N� �z1�mx�٨C�M8T�4�.��(��JE��+�3 ��L�y���ٛ)��T�����%U�<2Y����A�f`@�.�R���c/M�1%��z'�����i�p�]��q.p����+B�����*��?���蓴+����ռ*����i��*�0V,m�  H��lky>gG�"a��em�z(��gQ���b�7�W��U�}Я��l]q�F_��E�a�ULZ�Ej�j�|Ŀ!X�ѷ��i�{}}�{e]��U�2P��}J����ў�4���u%�tg�v�Ռ�Wp�����nE@���/�����L�2o�Ń�#���s��u��K��s��r��03���G���a9��V��o��,M��/�����"�Euʅ{O'��~-��Sn%���*<@�|dX����{�p]�@�����c�됳ֆ�ہ*�{�~}��=�����B�;84��<��u43
ƪ��4��n7\��6������e�-��ye����#��ը*�}������2QE_`�)��Л�FŽq'2М������+�:��lyU��ԁU�l X�wg����W�䀵���,�л���;�]�T�g�\��Ҙ�y��0Z�w��"3"�����S�0ͳg�)�m�[۔>
���5aC���>�"�����l)�W�q �\ xe�}�fW�}|Q~hFw��9�{u�N�z��B�u�Z�����F���7G��7�`�L
�
h�ֶ�1w�b���N%�/,(�ɛ70r�8�S:)%G��6e���E_�#��Z~�{"[��p��ݣ�=�ZuR�'� ��*��/"�ʔl���kdT׋�;�`���}�	Ik1�6wA��pФ�&;6�Y\�򠾺Ⱥc�FG%u�P������&�D��%2��0T����t&'�Xd��0Z������Bp)�&V�}<���
(=#S�����,�Qe.G3Y���""u��Jf�	"�5�����3�S���NU��"Ko��S�ǚ�����`�)�Y<�ǟ$1��82����w�,�`�,6K�@��0l�:��:���2J������,[.
]&��n���rE�R>�ֲܻ��	�Q���L}��v�?~%�H��4k��I�����^u��>:��@vvV�1V��^�P/vd��7�˵Y�B#,e��"�.�[^����%�[�Kn��~�$G���WtT��%A�v���I��<ƾƍ�VC��)=�Q9���-A^[��<���
���1�<��Ӧ�)�c�J �rY,<pl-J�pQ?�J�;���x��%7�C,D��g��0�HF�C�M�w�lH��:cn�LW����j>�̮��&,�L��yI�7�f���L��N/0n��-z����;p�{%���(��Љ�j�L��rB�/�6��&B�W@`��%�� ��+�k�Ŵn �dG���8@�^{����Z\�v���
_���Ӹ)7�c�s*>�>�w0��"R5P!���~��Ӟ�a#T˞�ѱE�1!)f�b�a$̒���ps$m��z��d�ds�*!�r���7su������n��Tc�/]�M�ʏBF1k�
z�U�����EeUﰑn��Y&��J~Z��ME��ݐc���N�p��*3��cL�!5m�ut�Y�C������)gLy�ʔ�}�]]'�H��Pwឤ/���0	S"��ȧ(H�n�1��*�p� ���@���2�p�e�n9����4>��L��G+eR�g6���G�`�N|��ڜ��~3Z�kd�ܠݨ�Z�7��E��3��`z����������~��u.�[�f$)�J��e}ȏ��Wf��aצ�|)��6_�����^��ָ�e����4y+�	mC���Z]x�&1q,*	*�d;�_Q&Vc��16&�`1����G�C������cT(�'.0}ʜբ����* �<%�5�4�����M`�1�~O���Aa�k������:�B/MIbVRr�!�52C�5�IK�O^S�m9:��ۗE�D�Y
V�d�V����?Ġ��c\SJ�F�aoyԾ��m.���K�gKI[2��2���|77�%V�>�Ӗ��B�nC�S�}��k@�P��Ǟ%{�d���-�5��Ab&MǞp�p��U��?�6���`˽+�w�?6L�{3����:��=�����p�v�ps}uh�Y�3�$[5�ME N0��D� '/L� ����>�K~�J�(��~���b����'�B)#��XV�X�H�:��>C *'n��QX��Gb�'|��1D����1+.��}gv��