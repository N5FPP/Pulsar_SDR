��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY�5����p}�"�,]<�U�5E����6�]G�p��h>vR�Ic0�ګo=��'��o�!#[w�y��(e;�����B<Tr}�bS�4��S��ŞR�<:)@x��.����ߕA�dcp��QO��QĥR�}�	��H�Y4`�|��ZdC��vB0�;Jw'oU�e��_��Mk(rx���O��Y22K�\�Le�ٞ��m~e /�4����m�!)`8����e��^����R���vUsU�\6�J�NW2^2�A�bª��?n�p�w$)^���o}r�4.e[y���G<so����֢ڄ�W��Nc��^^�z:����"�T��"IE(B/���6����f�&�:����#|.-�~8e�ϛ&~\F��i���jn�L�-�O�Q�Cn�Sň1�:ۏZ�m�y,51o-Wv
�i�ڢ'*� ܌�
\��?Dp��um���~r����%��
�+����Ҿ��28b�/e�����|[w,�2	^n�y��)`��5b�n���H�����T�������Q��HB���P;Y���x��tUb�]ꗶ�@;�k���V�6_�^��\��9i���h#�F�E_!���d�易puu��So������0�R�W�_w��֥�_\=#=J .I�I"�1�fR#�n�=TM�O�d�{�̣����W����y_[p�T�����)�nf�_�w�oo�W�-4OV�]���J��p	j��~��7��Z:��=̟����9�-w���?�}-��uo]�3�#�H�F2�C0w���Q�4$$�(\��Ʃ�M�O��]�]�Ӈs�)kM����~��l������WoL���jS��ي�V�tUsv�}L��+�Ƙ�R��Ғ#`��Y�^���YeD�^x=����h9$�>a���0��E*.2���G�U��� !J`0F�9��+�>JRa��u�n@�Ka��o5:1_�c�f:\�z�?@螽O�@����6��� �}[����j	E1���U�[��1��s'2��y��n�;'®׻.טGX�˙# �1ch\*gݪ�T{�[�D����u��EW�Δ�/LX}�9n�6��jSs r�inG#�?���9��U)P;�Tؤ�}&��T[�c� ��X{�~����C����FDE <S�fw4�},Nn�g2^��%MSE���Z8�JlWL�*x�XB��1aM�����#�=k�8oA�*]8:<0<c	��ݭݍ�����'�S�Z2�Ÿ��B���&�٦��U}�N^�� l�	��Hh� y���n	S\haYS<'e���߈���w{�O#�&�W������#��өGë��=��'5NR5�^(�S��1 I7F?g�wb���d���U�dc��D����F�y�ðT.-�h��$�ڱ���:�d��(�����* �
!ň54W446R|Z��q��>s���
4ʠr��'q��4F����^* 5H�֏|��`V̜�6���ĺ���!s�
��K�3��Ry�s������R ��;qt�8�gE�Ίf~݊�I6��Ь�!�!Ew\���ic��+�]蓟_]��oBW�~4����#x����Zfw��G�
r�H�%�A��r�b�? on�W7��zpA��e�KЮp��6)�y*�� <��0�y�W_W��V1�0��HK�H/d]@KL�{bV�a�.��=�MZ����w�	{�-���(M�9,�7�>}��c��ဘ8�����[�����8���f�)��N�|��������Y�O2��VgC��+	B�m��6x��Fw%r��RWf�s%Mv�ǂW���/�ZYI0xc�ǋԴ0��U�3�Z�
�z�3�_���~�>�¡�?h=;eک"(�lL9'�l�KK�߸�a5�Ǥ���)�Η9A�i�R[WGQ`yk�MmQR�����A�.H�
��<x���i�����a�Q�D�KT�,:�˱�G�9���ţ��H��ĝ��=.Ny\0�9��� o)����Q���u��?J�`C s�\_���4��^�[����'��A��(�����́��!c����F�H��nD�R��1����~�:^�^��^�R.�Z���gb�E�z#�s��i�}f|Ϲ��p6H+�=M~��fS)�M�d��osKe�x*�4�,�yKݘq��K�c�!5,�	�Ά�TUU�  L�jGmT��ѐx|J:��z��,���Xl	Έ���j&���3X�&p�<tP�B�Ɠ
��<赋}��,�\��H΅��،ರ�hx�R�B��	fD��������kp!�4S�rZ5Vߦϻ�0j���O����3U��dt,��v#�v��a�׀�<[�<�ƨ+�3���Ӯ���"p�h&�ݗ�V7b]��V �&9���f�@���iנn8EZ�]�X����Ŋ�\��\z�C5�TL22�z�O�-�	�É�+���zDpM$�	�v����b��)q��ݜK,�皨�X�CwS��U�s��>C�� ��I��>'�f���ڳ�-���*�/���yU�116P��.K�h.�,!�Ŷxo�H�P���ʈPn��zj�2_��ΰ*:�ݿEx�+R�փ��!X)�4:IlX�9,�؉�ɬiѧ�4�Lnw�}��B�W4��ܷLS-�٨و]�u����zti��{�Zn��E�����$��bݰ@V���+U�8�T��`'�o���H�m��(���)���m/`;���?��7�����W��K�H��{̊�\iMM�)h?/[ɬ�&C��T�G�&�ɏm�=A,�k�1;�rն�-���'�p�jV���׬��SqR*N�*��|�ݪ��U��u@p(�g����uE�06�kz�Qiu���3�E���!�I��V8un��u=�.k�m$�T{-R��=PS�B{��p��?�J��"�VRx D9O���B������ �AN�spj)��Z�h��j�˿�x&�ϔ�z-vj�YK�{�-Q3�I�m�
Xk��[e�̻w;�T��P�3� ^=:��B���fn��Q0�ǿoe,MPdg1.tZ'��}%�M��݈P�2�W���H�f�_^�Y�pX�,����zwT�ڇ
!�a�G��KHT���*'�( F��;�K ��p����e��#��a�%�vä�5N�Y^���#w�<`>�!t��ٮ�q�റ�!"����vl|�I��i�i�~��J�nK�����gK��J��vI��ia�+=3�t��#;D-+aXX�^����ˆп��˲���+�vl�����Z>�b�1�SNQ�&cs_�'���)Y^��%?o;H�����ѓby��X�Y�K�_��0�«yW f}6�������Z4�^[�=�?�e9q�p�3���+��<9N�m���[6Sw�ѣ����J(�(Dx�b����u��&�Z@
�:C�~�����bP��f�2�բg<��U�l�ѵ@z�sV-ۥD0���|�����P�a�q�F6��T3H��dJb�6�e=�:�V+�?{P��I���
[�>�ܾcU8�������^�$��u�C��V���d_��.��[���r�h��XI)Q[��ͦ�n�7@1��޿][�>G�?ӊ��l�9J��.F+�wB��\C�ދyt��,�u$���`w�R�L�#A ��uvt���	���W[�̰:�wG)ƪ�����c�D����7wO�Z�q���e�ԁ���l)��t@�V
'(�Ry� �$m��<�0��jJ�lr$�I��+$�tZ����T;�����^u�E8�Tiq�Pr2&������4���i��B�N�9��.=T���(��I]�g��x�������E�}	�
T��K&�����Rh��2W-�$�`b��(��3�GFN�5|�����*��}~�zM����V�=/u ���d2�G����^�pQ���4�"���VD��J�f�w2sA?�&e0��j$��|zmN�n#�����ZV�V�IR�e�u.��"�g�$4����Zߓ��ho���a���.�G��A4��2��1U�:�p!�����+�MK�ʍ|�a-SJ��M�Gh �qٶ83q(�c+�85�yR�%�����ʚZ�ʩs]�X�y���+�w
 ��D�e��Uea.��:��S9� ;�)L��-�5�5�Ic��-�R�RUi�c,��rٝ�<b*R9"�@/kY*'��ҋ�d�xk�6K��`�}�� s�t�A? G�c�Y��32s;`������C%B�̶qRyʾ[>Zqh̔e�RH��QrB朚���2�58x�z�ƾhg^8�H�/����F�ߎ ���c5-A��=G`�*UG�4TO��*�-�.K��N��m��H.�!��w2&���
m`�&�K��u �F�B��"'.vTJ�=
B �1��p�u�v���,T�U׫���u�]�S�F�sek����7�9d`��M�$ґ��7(����4�$���I$t�yn��.�#KD]�WI�7N��CR�k.�@r���)����&��T_���`'����;�\��]�:�I�\�Й�jP���"s��w-�T�8�{�r&t�5��.cl���\+<$ú�u���/�o�Qh�xD�&d��b��հ�㛄�^'�)a1�.�<�'�#��FfP/�^31
�BuE�LN���	��.*������e��fڮ6b9f2\>��jo��<%?��$�dC��ЬX�^��.� Xۘ;�����glM6�|N��'߸�p���=.�v_��bZ��s�ަ�F3��%�����;��!�0ͣfG=��Ӯ��ᖶ�G[m� ˂���%v����ݰ�",2�~]�m��f���s{q��ƚ����6L�ٿGF\B�6�؄,'O}ut���S�.�+H�^�R=A�J�kw�Z1���8��hŢD�&����Ow���G�j_zx#��Y�%��P���r�5ܐ�xP(����ߠ����L�ԿuϬ�*/G5�mb�q�Q!��W���O�M�i���ݓ�a<2W"���� D����{$>��0a�����"+N�����h%�g(��w�2�",�n���f�%JK}Fn}�7o�#�a����P�Jc e�ڡ$��@�i?j9>d&��)��#�] ^.���uz�5G	�b�o��=c��R�B.�V�QĚgA�,9
��L�r O�cg?ȇ���|��K'-&Ȋ�7�z�^��_P+�&l��'H�*�?)����+��}�suK9���3R��e�P�����XN ��d5�o,NttL���SȰ�
�{ aY���� N6�Nl�;�s�W���a���t!x�i��<��<
��/}lͲZ��&6*�z�"D�� �g+k�/ዶ��6*����A�t*vo�9iY~Q�g�ctt@Po"�ܔ�Z���y�9��*��Dm�:��%#�x��yq������WB,����@�n8�e�ՆȜ�ծ�o�sj�nLܲᥙu!�H׈7|
n�cM�����3|�y-��XiWaz#�VvH���
�����8�Q��S]w��or(�������2G� �|
� k�m��J��̀���u�I�VKOsK��М�o�Ss�cA��L6�a��w��y%�Wr^]�h�|m�|�8>f,�@)�/��������m=���e[!FF�37ʹ������O/�M�X��`�� F�;�E�"n.�Š�ɞ��Ҡ�Ï)����ra�(\w���_/Y,,c-r��c��S�;l,`�ٖ�P������µd=8㊔�*:��g̾����`�����d�'-v�oj�
��ʲ����H(��)n�}ӹu�7�Nɿ�ry@��׈fw.҄)�nK��hznH��o"]r,����1Z��q�3�oݧ�A'����a��V�5�0k�Ώ�Ȓkzy*94ޙ
�FvE"mas(��Q�/�[y���0'}�'�~`Jdg��/?]��ku*����Nࣶt�,F^�����ÞQ�0`���R�f)�yr�����"�q��5����"��8��@?hR�u|�m��G��n����2�n]���Un�X��.��㚼�	NXqx<펁�C�{@4��f}h�м�#�ݮ�Ur]�ߡ����*�ODy��������Pϰnj߈!rB.��<��WrBX|ո�ؤ�˺<z̡{��
��sl1q��Z�A6���z�J`�M8�%�ntk�R.G�yi�ʊEn��?	�#��:ͳ��O
1��
�0���F!�Qɵ>H)��L2��\�N߱����,��c�`/�T��o���G�5H�d�����P)�f����m��-�$�e���5�ٚ���b����R�a---W�COV�V��n���V �� �(�k�sJt{�ӎ?#�-�D_AKh.�6��0+'�WjO��sAcS(�:mi1��E�n���(�x��6�����2�2��5���9��/��'_'�%��F%��>��Z��I�,W0�!��o"�H�DFpw����O�ή����务��W泵�]0��a�Gl��9>/��W�;M8�4�V��c����p�ȟ��������6,�����t-ݳŜ{q�c[�I����MZQ���awVk�,*lmA��+�z2o}l��+]���<�Q���y��� G^c�O~.�&�IX�SVܜ-5aX�f���Ҳ�43�<Q&��o/�6�
!ҫ�:�B\�d��(ԑm�^7�[/~^YJ��Ks@�̻�+��