��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY[U4\}�(`+��s���k��T6 ������z�<{(G���l��{�C��M"$�����1���4�*$##]_�w�`�AK͓�oek��%@@�h������ހs�����(�U�̋`A1}0�C�I�� �҈���~��(�����ZT;�����E�˧���I�Z68�C<A��D�NI���LUdLlTOk~��S���-��n��Kn$6�� ��>��#�$����kt�*�� :6�5uk��%��"U�"�~�>��I��%pc�uFm����YQĮ]������'�^�j��LC`犀��J6�����]K��*�����bϙ��6�p|K��B��<����H�Cc�vt>5��$gZb���9�#"Y�	���?$�/'����\���M������h �h};��k�ff����-��5B��DDΕ�l����V���}4�I����Y�vM����;ān��ž�ۊ�jcg�����v�� 9��5v� �/B����V�^��;�@x�W
�w|�r?���4�M[�0Y�M����:�*k̇�/�B��U� F ��%��rζ!��i-D��ʜ�r�%���q[���B0_:Up��P#x��݅� ����r��0�H�}�'e�*n�WzWB�ڸ;����u �@�xLw)@�'w;�_��U�[����U�I�9�����~Ba��X�3$KR$}	%}{�=L|bB�3Dzk���o�J����@$P��az�˝��g��ԫ�{�AÎ�}�� y�UR�a}0Ny3�G��t��w� �%\	��4.�\����N2<E��uY(�U��~L;��]	�}�r	p���]HjkG�C�?�-��u)��'s�hV�B���9�u��,�6S!�f��
�.� �Z@	t��Y&�>�.1@�	熏s���HŽ��i��/�>���m<�^s��_%���`a9H^�}��U_fX�����e��m��)~��VW��8��0A��4o��ژ��[m���y�\b��2������@��e�`�,�%��5+)d(�ҕ��j���9����n��P��K��e�`ǹ���C']��E�Q��舻���c�����d�f�ئM�J
�x%���,T�V�0�����Kx���e����w8��(�2l��H���f$��{��i�-��x�,��W�A�8c�4�P�M��d���5�V',)B�~�$��d`^�Q�!�8�4'E��:���z�_|ocM�#�`B��跩���q�&�c��<��AR�Lx�@�ێ7�ae�Z�qiz$�U.�Y�=�
e����;�%euTHQaD�1���ukؒ�1�4��3M�����88��$ {
`ъ����&V�m��"א0ר�7:W��6�A�p�{�Mg�&��Y�.�E�\�܅��H-]���p��'�#�Șv�~�8`����6��Vւ��Z�t�M�qg���.��򚮼� �(��� 3)���(1�û���/����
oiV۱�<���Xj��g!��$
������5l0HZ�is0SԘ�O���?v}����ޒ��n�M�'2�]���U[��l;�cn|7�R�,u��Qά6.�-f�w��)��㏜�v�6�2�a��O�P����U���,Is�O�F;�4��@����)C���͗�54G��EE^����s�t���̜sz�I�1/E��ݰ�:�t��a�
���k�AL
�ُL�u��Ɔ4�Ԛ����L>���M�]m}���u� yW�>R�E�D�Bv-�{�8��q��Y��zfG!(�l�r��\F�&�N�C�g�nE�B}<l�:)L�j�����v���y��>_4�5� U���Agآ�j�p��\�:x$���o._����硦Ȓد:�=[Թ_���?Θz�5�o*M��)��&�E��[��Dq�/���L3ส��d,p�#!K*a�o����4Ё0bx����)a�uV,\2�h��y1��+,��͂�b<���@�J�4����B����O��qcC���$����􋠗b,�/��,�ks��T`��a�`J4��\���֌>�ocY�
����Ql����(�V���Um�f ˞��-1�S��aǏ�'K�H��[��w�F^��
O��fN&g��@L �|�˿+9���VAEy��!���OHo�ə��a�r���}��X�b���v倝Ou�EW�\�f���J���OB}57��ܮ�9�R��v�ɫl(Mވ���w����C>i�&6��~e�t�b��O���{�Z$���;��w��0�p��o�5�1�FW�M��*��i*�<�}�h@GN@Yj�e�̺�<���^i
�~�7��;!�[)L0Kq7�[aN.ϒ?��5`�xq����|��	����M���8���D����ip&�qR�SV�u�s]�P����"K�fCԶ�����/��H��A�~_|��H8��>z�{S0�:{ї��K��=�
����L��t�[p?+3���fٗD�@թQ1Q~c��ǃ`	G3�[m���|i���U��F�3�gK�ŗ� �F����9.r  ���;�s�̶���	Α�8]�+06cZl͒�6��� $<=�r����yC��F��	Q����l��I'Ub7[���Nmr@wT��y\j���	P��V�R=����Pٌ��czz�wo�b����#����0�;���	��!���{]v�+6�J\i�������'v3�����Er٨nJ���u�S�B����p���g��T�T��٪եrG�)kFVOu�CG
���t�`�[K�3�
�׉H���ҩ��x7�j���A1ԛ�}�!dA��9�q���"��ρ�qyT�R���z�DzV�Igk��%� ���v�<t�#E��>-Y�M��34 L�������X���G����p�1�߯%�������&�ֲBZG$/��A�"���׈���ib[1��I">բ!<�PlH1�?𪱺�D!�&�^n���G��P��t�4l[w����d��@�	�ק�����x_�����R��H��T1v��҂>mܱ��CJ�A\�	je�iv{\2����f�1�����n��H��PԞ�nW0g�n�g��by@���*q5	������ \T��VE�3�х�ֶ;�屧ݥ�1��z%�~�n��Ѻ.
�(o��ʋ}W��ݓ�����g>ݲ��e��{f�MP����}����P�uo�I��׫J1Y�j�|�� �ܪGZ��A��X7ٮ��R�M�Ȫ����d��Bƹf E�bK;��s���!���O�����}nZ�?	r8�=�~�R0QP���
��g߃ӗ�P:ry�}�Y+p|Y�1e�-
�U\��(�R���QnR��/OM7�Q������Qcb�v�)�������D~����@謚��D�A(�x#w�E�t(��[�y�̥7c����X�0@�$�C�f�q؊������a	�,~�Ѫ��;x�k�a���@��4����7�P4gA�Z>b��W�1����<���r�����P���k�sD����x��Q!�]b)������\�K�:AF	��D?��T(�U���L�j8m ��k��ms�%m`��U�8���~sD�I��!J�oB�����/����$��_�BV��T��~�la�R��*V�kT�﵄�v��;�Q����rڔ�C
Si�\�ZyZ,̰�5O�y��E����/���̯���D�ª�4�W@7�L#w��F��XP�P��N���G�q�+]��@��j��):ҴZ�Y�Q�]*�sbq��菣VhiT0PQ&BG�&	��;�4 @��V���-'S��"�Gc�,��*����U�5G�\*�_(J������M���w��D|�P�=���}Г_��u�� ���_G�?��۟����{�YjIߓ+՝�~�l�!�B�
�0��U� ,�u����
���ڊ�#;�F�fTX���I�>�c���!g��<�S��`<e��߱i�����Y�G�ɵ�Rtֆo֢g�Ό-�@��<<�/�]�y��?�jB��	�c�$���l����.T�i2w���T�D�05�<<|��X���t��}�NA��&�4D#��ciM�	,��t��#jبܑv�P�,di��Qs{i�)I�L�[��R�"�Y���_b@ž0t��lޞ�Q�d�sdR�.��Q�4��4�P����75I@�nJ���B�i�����;J{���Wj���|��I�EY��P&��Q��c���w�� gʙ��	O.~R1��(��ߨ�2��)����H�7g͵%"��"����H�:,JhHw�08kjZ�ǎ+NL��0�N�i����5��-mF�E-�ⴍ{8��������-���=%ī&n�)���]E�zb�5�.G�Eڟ��l��G<յp� ��?0��*U	u����(��/<����+>�1��������H�)���5��t %6���w�B:6�`	���hgE.��Ak�J�p?��X�>fO����[[n��7n�KᅗJ�t�T�[#R?�j4��X96�H��Y*2�if�m-x�e�|H�re��N@��\��F��7 �6�ao*�*����}�"����bG�O�3��j+��O�:~Kk+
�����g`������(33	.r�ґ!^�������}Ǳ�Bꗣ�X(�D�=:�=�
�]������WFɶ-��ԗ]E ��tE�^X�0�՘�)0J��p|�k?(T�����0lP������� 5|���-��RCkF}c���?F�
F�|h#�������`Y��R�'�c`
�&E��D�tx�1~���)l�\:�U�[SBSa�]c���t��PTV� ��Q�)�)?���>�<e^<�V{s�ي���{�VD�U$L�.�T;P��Մ2��c�ZGW��	S��B����7�����"���϶8ql���+���.J��6�\v}�q��5����{c犡D��Tj)F��qc���dU���H\��ax��|dp!�����Oz�ieB-#���߯�����$0�ä���{8>{3��P�ٱ�J��61BfV<��7 c���@tЦ	�4���O���4=��|a��q����j,QS7��{Ҭ�8��<��>�; ����e