��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��e�ik3�������w$����g|��J^]�|&�`��3S�1I�	Z�����Nn�:f�*��Ք�:���o�s���Y��PVc�O�|�B�f��#�����4��u�C��\ �Z���C&��b�q��f��P9� 1���k� ��G�6Ci�%ʃ��}�Q�<��ZRi��ڪ����E˔H������**�5V��"O�U�1PSz�g��(���G��QYFJnZi�S�M�@���[h���:Ƕ�G��'�8K�Xj_�81t��LE$!p',���= �XI����$U���}��j����*�B���]�$�j�,�J7���n�j50.S�~!yп�g	��X��0Ȩ����m���%p�E;�[;�Ι� F�(_dzW��K	�)xĀ�K�Ѥ�>��������)�!��t~>��MQg�ͺ ����3[����;6T*� Qث}@��ď|���B>mҀ����4���P�b��ӑ+Bl�^�/>0�
H��z��h�,��\��E/�9ФZ?����6k��.��6��}�{*P�<8�р������5Y��_���������4��+��b�[H,�����Cg���˝BX\
��ڐqB��������g]���Q��_|�{��ћ��mSX�z�i�"�(��]X��l6�j;����i�&�eU$�S�	��i���t�#��}X��dF�df�b{�{.4ֺ_�S�_�t�䘓e�G�	�N��슓Ʒ�_vo�B��30ܡ	����{JUZ$_d��j���p���"�*x���w�My{%lGR����o������diR��Gm�aaG�1#$����ُ�6i��=��9�ˍu�ˮ!�t�� gi��	%��%�-X�_�ԡ�"���\�)��7��+���Z���@E��D�v��Q � U.��=��\�6� ��D��Q��Xtg<ȑ0������C]�-i|]Ӫ�x�dWȢ<:q�a�Jz��t�As��W�wP��95�/�X���K1�>��m9�x��������`lNC ��".�|��Rk�Vu{I"���n!t�c�S�5;�o��K��S�V:&c,���������|Po㥲��ߡd����y��X~���J
�E�������0�O-��	[8����H�v�͵��c��M�'ʪ�ӡήzl둭&����+{(�5e�R�7�kz���B:6�5�lk�r&�!��7>�&��t����jz9��O6��i6;�#k�F�y��0l��F�m��h:�6�������|��?��ם욻�|NW+��*l]!��a���FkY(�ZP��3��S2�rU�Ӎti���HB�ј	�X*��N�K�N3�!�'D��g'M'9E��h+,����45�$�:�I���}�]b~��wg1� 	�����:�E�%Ȩ��x�+��3�,��͌)�)��4ZU����;wh����e�է=�G���ʾ0��5g�>&)�	."����RS(���ީ���(���Ts�-�!�oTY�f$�C)�8�T��7y`�d\o���]M^�*(�W��M��!*��$d��/�m����>|�{�$���th��#;<t9�x2gG=vި��qN�&����`*�z/_$�H�*1��殈�O4��bs�V��?���
3�Iʬz�dW"�ަ]`�q��	�E���n����:�zP��auN+�Uv�{ql�\#i�t+�GoK<��ř�\��E��n�=3����n��a˛�|��� �ง�r�-�M���j*"$ͷ��-��6������_���bG�]n{Y��m�����'�m�<�Ԉ�W��R�������a���U��C1^��k�2��>`��r�7@<�GBc\��������?76��>�ޟܼ^�DR�%��)ZͲZ�� nk�Eu��[ w�� Y�7q���+�P�Ix!��!6�Ѯg��v�S�]F~%��K��=j��[�ʥT�#r�H�g��m_��\�9��9q}��X���V��xO�|�dr)v�D8o���O�`�1;|����?��dֆ\M�����nSӋȬT\IR����Y��oP+1�B���:R$E4�`-M'�lRE)5���A���>��#cW�=��r�)��U"�.�?� ��EӔH�nIثUPkX�O�G�k.;!:͂D#�	���n��"�5M=��pT5)hW�Rx��ن�4��2�C4��o��}��هKfqx ���o���+��e_C�~4Nփ37��U�ʧ��K�FBe|�G}�'�4��Ε�8,�ʮ���B��=��B �$y��FG��<~�T��T�*��fIѻ�v������m<�M�	��Δ����8B�
�X��t8sS�M�����:�(�m� �߄�5��)��
B\�l�Z|:�fF��e%K@�ȹ�����hZ�=ٙEL{�O��a,Tx"�FM����gJ�G�!)2��?�`CR*�U���s܀J:����S"�Us���tF����-dP�-;q�]4�KdK�zȳ�E��쯛��Q��!�/�m�3�=���H�C|�&xs�
֙�aeA�]��A�1���|��;}W��J�u9>q��q]^�XB���g�?=�X(�9��*�(�ۇ;�/q؅p�rq��4e�d�KcJ��O���<��v�O���/T��DV���z�Z,mq����oX�׉Xլ� ������f��o�˱EԑMU�Ɵ��g�[��oѠH��5 g�D��T�Qc��Ê�1���.�ɪ�U�:��YhKҍ�O���ReT�қv]\k��'�Ğ��WD��1wh�;�����/&G��ia�-<�//nku�Wc�>�Q<�5
�<x�#6�K�6��u^��P��Ί�c4[��=`�]ݚ�
����:�n��"��D���Iv�俦Wz|����'9wd?�z�xF+!Al]��q>9�V�(ԖM��~�D[�z�lLCn1�@(����ȭ�V��c�t�n(Ds',&��ZZ �|��ؙ�a��d�b�����e���"��r�3���<%���~|bb�6B�P���T'��c�&ZC�L�L�R/���ʟb)����U�=�K䠍�Oǎ��,ķ��*��O��@����W�7 �~]ALs*g3+¾�^�k7�R&�"� �Գ��=Mb���'W3�2�e��/ȿݫ�Xтт�A��hItW!o�n)�/~�'T�B`�Y���P�̇Lھc��3��X�HI����p#}�ٟ��Wh|�b^�៰y�~�w�`�(&Q�[8��;����"������q��~�BvL��Ip4�R�0��!�J���������e�a��>�Rq/�q���<n�\ۂ��!�7%���E��1;����K ��
��V��X�|�ԙ7m�`�֫�I͘� (+�Y$���۴�hGع�x;ä�u>��zO��A��$s�@1t�GڋK���~����&)�[�H��x���l���D,I�#���a&jD1潠��X6ŽCt�ܷ�>&4�K�k��:M\� sQe��U��0��Ⱦp}q��b~���N��罊U,��O�v����|�+�p�5PA�$×��oL���+m��7����a�����/=�t��ot��������#���$o\|�p�N`���6m������2��o��y`�i�-�?{ˤ��ʌ�2�վ��rUҕ��P/ͳW�X��>�mX��=�&`��?�k�k}I�z��ϢFU���m֍�Z����k�:�5�����ͧW�(Bm�*���DP>>�#X!���fy�Y��/��ĳX�	���u>��Z�{��`�/���M4թ�6�������z�?���j��_���a�������{���0T̚���Mo;,��u=&��q�L��%q��b!17�&i�6����l8�W��A�.)�z7�ͧ�޾������Č)�h"r�֡ox�o��^҅���/����Ǳ�JaX����{oX�N-�W& '�����t9�7����NR���|^E8������#�i�
�َ��V#���O�h��@Xh��h���Y��>��o�eq�2M2k�'��TxSq�J�Ӗ�ئ���^�U`���E�`(������:��c�<M"X"^N�Bڒ�*nM�!3��o͊����p��2�'r�o�Y����Y��;^��񈓤�(��ˆR-�8u���$TG�P�!�A�K`�vg�U���+�T"���}QbY���G�J�,y��z���/�aj�8,v�l�wx48�,��BW@�Wa��懻�ήvv�5y�W��B��_=-x�[�Vs`g�#��_�
'�/kFz.&c[n�X��t!g�LJ2�|�p�!�@S<�(An�kVӻ�2�}��Ϭ�D^B1��2r���Q�meZ�J��������6�i����X�ld��V=�B`��a)�dc�`�Ju��Ǐ��ҿ��)!���CF
.L����S�[�6N^����x@4�Ǖ�0�h��� �tL�r�+��=@~�������9�;�X���d�ÒP[#u٢�xh`2�xk����a����kl@��K�Ca�	�jG��H:d�힍r��z���
�� ��Q���m$+��վU-����l�QB��Z"��� G���F|��zi.��,� ya-�������V矜�Q1N���9��Ξ�~k}���i��c9]E�UOtd�7�|��{r1un��t��F�M��F
���K7t|�g�o��8�x���l���	���"+Cל���S;N
�^�>7�\��%�3�$��A��u�U�yNd%-:[.��]��*���x4����� T�3�f�cˍ�%��-��m�ܭ�J���x��[�4���Y!Z�DU"3%�񒽠��ײ ��	E�6`���?���t��K�#�μ��ȷ��r�/��a}v刧�u���##Q[A��Oj���ʐK�c��;�]���T�AN!M���=53<�����J*z��I�QD��4/�CU����h���^��jg�i�^���bJ ��j\]�8����]c�>�z��?v,��Lrx�X�Dna�?D&��?��V��/�����$>�ɶ5��Z��g�%�eQ9��
��3Z�R���b[J��&R��'x�}{V�-B��xnk�סL/A[e�~�.UOdb���M,��k�����'N�Hv}��d�> W���n���N:�(��U��X)��K��#�g��C}����d���ѭ��K���"a#����^��������W�W��R{tX�E�4��O�ݾ�+p����s�É
j�E ��7ɯ��@���d0�Vx)m:��@�m��Uet���	��f�Z��b7� �Xб-5ѯT�C��B�5�M!G=��x��ɊK���6ɒ�5��	Dfe�������΍�d�@����
O�p��vm��]vIC%Ԉn���)q��#}hvWc��'��K�~b�	G�ETTX'!��@�!��}������.C���D@�:����g�`>���^��e��)?��v�g�'�ш��y׺��i��g��Eδ7B;°�3��e��7J��C�k6�����#%���d��L'LEQ��י�/[<�U�$�AjQj�<$[� �CB����(��9��E��~k��#�񹺨Q��>>�Un8����如
��dL��
�_�VN��MG�h|유�ՁboX�P������v�:׌e�S����f�@B^�sNS�	h5
4�h8Q�L�]�\�p���	�5{ ��=
y�G8�����ndsh�����}�^l�!ij�Iֶ�Pd԰�.m���,��!ja����ow�1t���k�����%g��%r���!ƅ��]V���gueU���?����U�{0�N]���fߦ��;>�w7�A,���y�#��J �sp(~�q�e��1��6����W�X�$p���� ��u���۳�����c�a_�8��ab�N����g�'_�\)��I��z�c;��=�����%zu ���V��A��CZY��̞:������X��H<�����zx�����/6�;�`��%c��c�b�P	��tcoft]/���Q')�ۊI|����kk������4�A������Ό4��Փz� �É�ʵdzF�=�4���@��uY�b��>4xY����V�B���q���GS�[�O��
�e��qaB����5AK-=�Y��yT�>!��X�lW��]�-��D�15�ׯ���������֓*ү����T�쫜R��z<�F��lQ������W�(��<���0ٚB#1w�~�f&� Cv����N��wv���j�~���	6�V��-���g�S妞$NP�!K�B2򋀉M4�(o��a�pD�a�6/
�=I���"X�4�f�u�M�;Y�=|X��V����ud�\�`tc�k߶�b�?�
�+i:��X��Yo���)�K �9G��>�놚�i=�i���X���tSU���ͭnt�����nקDN����g��{�m����X��-�cS���~�����s ${;��7ټT6�;
y����������o���e飼��Ѕ]��gA�e��}ww���F��`$�M9�:ڶ�����-l�����h�ٷU_,��`�~�lS�1h]A�5�̳��yvv�x�~*Ԙw��P���sTx�գ��'�Y�ePq���BA�x��9��d$M�^s ����;[,G�#tTG�9�C#��"�a-�i��^�!V�wi:���e�I��YL��ڥ��׉;�<�C��t�'�/Kf���.0E��W��)�z� ��s]]܊*�s1�!Q��Y}ջ7ڴxs0e+�,�e{ə3��W�YJ������/Y)K��4	bn(�*��:��Ʌ��үuv�A�GE -r�*pƣ{���Ŷ��J��T��i��W*��"���Ϣq0�o�^p���7{C>-T�-vB�Vu�9�\�����w-7J���N�L �:�j����_t�f�9"^˵*�kW���d�O�h[��yT��l}�@�S�Xʝ����.�d�m�I��w���ց�n���)+�7��%���.GF�`�`3(�߽�^��a�hm��<� �H��qf*�t�^��H�Msiz�T�V�>�U��	D�MQM��*Ѥ<�V.�}ՕsH�F)Z��U���ŴB�3F��!��B>�x�r���x�s��-t��Z!��/�%r�W^Igz��g�����RX��]�秫B�b͠�#6|�G�˱Q�jń'"�f��g�}I&�'�	��6W9��R�8���H�b���0���`s���/�)�b�@�J��Q���(}���r`N�|C�2c��4�� u�'�c�͡*l�%���
n`��=��Sa=W�L"-���"����a힌*��o� �P�1���T�`J�-k �R�ɽ=U�nu8��p ��]� ��,z�𕄥O�	X��goǄ�ja9/��X|K��k(i�����膜-��ZSZ�`� �
@N`G�d��<���O8I�J�t����V��ny��HĖ��C�����rc���j9���e�{5�$	h#��.�gĶ9:p�Z[�l��E���Y2K�X�"c��������r�rf����WY x�IYTٚ���R�n���kܹR��!~�9Gk�V8��]�[⠗�i�A��T��6A����	~B�1��)�خ��|�4䫋[��Pql����	���9�䗪�a.i����kE��mY�K��1�ie�o4s[�r�Q��D4:��s>���.�׉¹��+2o���[)a��n����� ]ߺƗm����}���~ikv�07�~\7�O��yŭ�[~�8�)[�Sq/�5���/S�;����-Ф����:M�T ���_�$'Ft {�j,
p�ٸ��w�zY��9��:flR������-���u=*C�"�|����k�ֽ\����M�)�Sh%.��'�y� Y�
�t:�[M7Ϋ��V�a�5��ڢ������X7E9&T��G��Rh��Z �@µ��j���(�A�m��<L��P�E��8�����\c����T�Ő|О|$l^J-�W3�R����+�v��S������ߩœh}�=_}�<kH!t�p�so�kuDge��a�1D�[>���elw�/iYKDe[q�f֗�i�Jx���Y4 �Y{�;Ɲq��{��K���MA��ccL�|�sgu"�������C�L1���t�X�}�Y�s~H�|M$��U��GН�� �p�#J�z���R�3�(�Y켂� ����o��v7hOGw��#K�N��w`��B����	%�βv��e�On���Ru����̝�G���|Y1�Ra�N�mI�y�V�y#�F�v{��*8��aI�P�,�g"OW�_�C����n0�Y��%������~U�6���h�a?r{�x�n��ôƣ�O��\�	��/+�on��$�1|g��ްH7E��¹X^���YN��iؘ��j�b^I��_d��?�ɟ�������]���^�����ssKΕ�Z�8fr�M��1�'�Sc��f���$fM�j3���U�|.ڮ`�_�,���9��X��\�ZL%+/�:V�>0����vdp;O��H.��8o�4sd���K��T��s�Ƭ�(�Ρ�0�����P.�Zu����L1s�&��KhA������ճ��J���5�������H���;�����V�2��&n �cI�u
���XDyZ��ⶌF����t�Lr���@P]�Xsꍒ��3��*�����2�繻�nbRrS��S�X��I�ͶDM^�����c'X=�)��'�G���p(�5`X]���+l�g]h���Kt�����Ӯ ��{N��C�'۱�N[$�v�U���I�i�IJ���4�Rj�8�>�5������,��@��z��7Jp��Pn�r ��q��zE��'�Ud/�Os��m>�sS	�4ΝH�ݢZ��xTx?���M#e�6V0���pFT���J{ih�aȴZ�6� �&��QC��k�`�<��JjH��kݦ�7�3�T��FŁE�T�sұV3i���4�y�bA�]TV�, �L=v��ج��q,^lӬݭ��P����ͤ�}OɅ�J�
���,��ZF�1P�����9pd�͸T0�.3�c�0���"V�w1�m!7�>���H&�]`s��H]>x�Tɬ����(�1�����Զ�`��E�x�D��N��z�EL���� �w\���0廰�̸���o�Px��
P�U7����Q�۰�,>F�</P��)��z_���S����
)��tk�ӡ6}�x��""�*̳ۤ����ǽ9ױ�s������4u�q%c����A�$+��5v��^��&^�k�"�� �, �ؑٙ�u�����Hx�l[�h�<�_�H���J����,r�r\C�{ iɬ���;�4>�4����}?��٢�g��F7���q9�-�Äi��0>�7y��O��M��ϔ�>|����F蜃'�����8X�pl8���\>+�C5Y��1����_ND)	?K*p��?��� ���ѣS�DBC�g�����S�D���߂�\+������z�~kKé��r�l�iW�QF��y^IT�W@�i��K^�ЈpNf��j˕�&X��b�2�kB���� ��0]aO�Sb�Y篼v'�|9�2���d~�t`�1D<�G��S� �"��h���q�5�^a��盪��,#IQe���n=�o��^B��n�JϗFjy�q�v���a�e,W�!����1����9�$�翨����̪5>�02����MT��é����E6��e���\(���+��$īU�dQ���{3VW��J�8��W5<'�4?�^��<|��w�~f��v4���B��j60�烠����0���ܥZ�R��re'����O��a�	��/-�Z�8��ۃ���ְ͑��c�=�I��L�4�_�,��h؊2i9v�����#K��r1�5�:u���u��J�tߢ<�޴;����#��ʈ��L�"�E��p`�j���{�<6@���l8#�_f@O����m���ӻՒ%P	�p�Bf�z�7j�8����ʯ�+��jY�l6#'�s2lĜ1jt�R�v�72P��
�����,�^��e|�p��t͏� �P��]A��F��.�[R�~Jy�гF�=�W/�]�z�'��Z5y�H�r��fp�It��^�YK�*��N4����ܓ�P}�u6�֢���K��g���y�c-�P{0�l��;%2�<-���j	�4�CNG"��d�<I�!G�P�ɰ��ܷD��$h��"W�\ƹ.u��WQ����e���-ڀ������h�%��;)��0�H��
υ�L"(���"}���%Ս����m�]؛C<���8d���Y���y�[_�U1|�g��KF�g���>�`��s6.��=S�0ЪQ\B:^P3�ҕ�|������O�=$N��r�* =���sEƲ�X2��JRǰsR&��+�<�kD�w��;�p?����1&�ݛ����n���m��RY�G8�^i������HK>X@h7b������nf�'Ϙ�i�L$����-�vnp��<.��	�R���d���m2�Lp��Qk�,y�^ �IW�2��l�L:<9p$8�Knj|ߠ��+���لj>_�a�Ӂ���@ ���N6�M��?��"&�|Ԍ	I��)���j�F�Ʈ|#����	,�������/S���:A���3=c����}�fy,��"
����}8�Z�\��A�����#^�B��9VN]3i�T��8t74���S� �f̓�Yp:�`<�H���
%�Wg��z���{�fj�j�/�g`�JpY�Q{��E�8 �.�xՌQ����L/�WPV�x �7�h��#�x�Q�^9�*ߜ�:<,��kֱBW��XX\�h�v��Q7��H:hrԸH�d����b(�5f�r�e�A\��=��x\��
g���p���-���n�j7�
Μ���m��X6�n�#"$��o>Q�^46Y��]���_�Q,kmH��h�T`Ȑ�H�]�qE~�T�����1�e�N"�?˙"=���u���'�a�����q�6 ߛH��	�Z̑U`�cl��Y%K��9����l�ٰ/��tE��v���|4@��  .����~�M����m��8D��g��wJ�uс�BV����د��P9���ه�J����D�$��F`�%Q�*�̎�@pY��]�>#of�� !���볈�\�v
yZh�]�}�U���cH�d��gϦ���+�D�G~*ڑS�ޅ�sD[{9G���+��{,4�n���e~��U#�e`�tr/��
TF�1�q��v��?;�eo���a%u�	��v���83�OQ�1�Ń�ھ��IB��g����`�D�@��3�>
�b�48���,�-;�?7�?�"���XVe�K�D�\���U,d�U�P�&��z�<�gͣ�W�]xd�D����DT��a� ���Y�\A#�����%!z0`�,X�$6�UU`;B*I�U��z����I5�X�Ҭ�0x��l�ʖ���cXZG��c-M�k�Bfb�2�fjs�!{n7NX��
P��c�����)�{�]�^�>v��2ҽZf:�����Q�?"���`��dQ��)̄� ����y�������2���W�#f1R43oU����K~kb!ˏ�Hz;<���*��*v���M��Qqi��Z��v{����!���_��I��b�'>Y������vX�� �a�I�q3FXl]�# �67��e�H4z �r-U�|����M�+&�5*l��#������J����;� �;|9�>J���v��u����4'K���i����*�(�)5�g�8�ߜ���?s�&�cf8��C��P�(e�Ii$4\n�.ܲ��-�����p��N����S�r�+$�ZF[�S� �I�˚��&��=�\�!UM��3��&r�X,B���?1�&��~����q�3��	)������t��Opnab|��]���󂩇��5�8[�����<��I��>U4��!N]J`�5X1���(��T���Xz�4&�0���'.���_���v�0���BkGK��;���x�=�-���t��(�E����h�?�9>�J�4+�h�z�H�u�a���Y�' ��0��Gx��̅�O��u����<ʘ��Q�E5$��S���c��o�_-�\���/#`G�V��m�%���U]�re}Gk�9�I5=a���Ō����{_�fˋ$���2�����y}���2U�6�̜܎��·;�Nw��Ҫ~W�pX�s,��|g�b����/(&L����b���x�C}i$a��e4�c��Av[�Q�\���7"�ӃX�E�r��d,)K��Ca�2�h{�m��J<�X\��CDB}��|}�g��s��@�w��+!�A����R� �+�ټ+L5�Z�Ξ5��qkn��fA �;���g�A�HX��跧�tkx*�KH�0���{���o����H
(r��=��0k�)�(���U�s^��[_���y��5�<�$C;i�b"ЀT3������H\��p��>�%��ꚕ� �2CE}��E��cB1I"j�~տ酪	�R5˴�(��q7��K�*�y����PjN��.mM����w^�Σ�=�A�`ޚ��n�@Jam��=�����3�
8z�8�������̈m��^�/.�A//E���[�|��y����b�ڸ��a�"���]����drݼ�wXo1sJ@Ե-�'Rk
׈�a&V��͢�޼�px�"���{��m�I�6f����S򛃖	�]MT�QϐK��AV�C�4��R�%0�[���f�5�rj�y��E�$�_�)��4�����5W�X>cϼ�p���;0�[�$D�/���EB::M(���7qC���;�}�g�&�e~X����3�S��R 2i~�+:��Ԛ*tL�@�-�~b&�����R���΃A�ע2��Ƅ\mO�*�ǯ�[1�Y��k�[sk;@M��L����'���t��]��
�x���^��3>-kO��,�������E/�!(�6�� �b����^6�|�K<��Κb@��4���KTb,z	�}yS��<�j��W�r_�Y���������Qua����o9��#)��S���ף�䖕Pg�\����{E���������Zc.;�=��
����f0X@Y�׵��ޭR@m�|���pZkC��T`I�&���#Wɯؐ�3���&ۃ*�'��<sm�ͫV���B)�F��AA~pK��(+����\����!�/W⮙��b۽�P�h�r�m�_9c�WғPN��6]��u��F(��z�y��{�T����
ҧ�;goI�ݐ�~����B��PY��y`� ��1�p�Z��Tt6�l��;������Mnm�ب�����%WEed�'�7���_��d�%Z��3����?��D( z�*J��:�g������o*��JX�5&�oj�q�+3��Dƫ�xN�9��w��S��uc�[p��_�2�g�����n��1����^V����U�_!�&Ԅ�fĆt��4�#+H��W�(����3��╫�xcHWn���Dl$�Z8�/v�Z�Īy&ȕ���[?w�d9�l���� ;�������e�H�<���1w�u�@��&Oዏ#��0d��/��><-iX�VeĄz��o,sx�������Y9iaCK9v{�g�O���Q[��q< ~�J|%xF9�1�}9�瞬���:YW�����r���[��1����3��4w�;�e?�]p�����KJ����ja�h�ӷ�1sG��2cZi+_;�����.�vU;ٯ��ƫ��^g�ڰK
�����|�ޚ}~�y{�CQ���>XiI0�4�2���ζ|�]�B>n�j#�{c�3 �:ӟt@���昚PQ��0�,NOC�'�)?WWg��>,�v���y9k|W��9l�lP@��.C��ɡ��[��}���t�o���VD9_(�VxA��bzT� ��$\��-����$X�x�>�rC�pi���2>��;�iU��.�:�$���e�m�fW��*!�[a�qwƽ�6���f%5�Ւۇ1�8"L��NR��НS\,�%���7�* �ˌ�{���_R)~�f�I����u�6n8.�s�~���v!b�`���쉚نC�At�ˇY�Z"q�S)î�ꂣ�Y�φ�9��Y���m��W%����U� �@..A��ĩ!@ր�U�s�N2�xj%�@���di�ᵶ�C9YDhJ�?���}7%]w�M5	hTMՐ����\�|0i�%�d5_�!���( ��B�ތ�7ڷ_�3SG m(���*�./j�]�*c����R,�Wʹz4G�����bπD1�;����oz�5CM�ګf(����Э��86��`w*�G���by��N�����Uc\���p�q���5QYtʦ&���5�4CQ��|��Ԥ���4D��0	SJN��n�NcX@���^�t҂W�Nl�N�^���C�{�{� ��C@'��˟��JR�)G�v���U5`=��+� x��mC蚉9Ի8|)��&qи�q�#L-
���f�-�U��! �5�)rN�w��i�P*���Š/c������28�Tt}$I��f��A����"����<����/�<�1|#�<��*=�
�Y��c���1���h��~/��c���]^;�eF�5l�l�5i�J�����9}ຨ�C#]��H���;~�X �P����/hq�?�ˬt��`�¡���)������Fl,�	�(�!�Қx����=���:Lg�wW��,��t��DN��i�
H�"��d��#Q�8� t����V]��,�bd��y��h����c�ig^�&]����w�L�������SZa5�6$��m��~غ�Do�/r�W�Wߴ����뿒�t�C��XHk��B�}y�9�B�mdܭ~W�7u!2P٭:�i�C>ɞ\�*r��`;�yJ�Sܮ�f��Q�:������笺P��3�3�~(̵��U�8�(��s$Om��1ό��>�G�]_�ܜ�Ӛ���*c�m^�6"��E�3����LΠ*���B�Z�	t�v�烿N�?��zڃ��N%�T�yDFȺ�+��`����8z�Ð�3����b"|�W�����{�NS�@��C�7-���'�{�I��e5 �����P<�%M�U�d�t���O�2=�	����d���KW徯���bY{Xŷ���.���8�,
H�!�mj	�=ps{�,c�_�~RJ��O��4���.~:M�s~� �*�H<�`/\-�	��dyw�$2�6����pm��_	-�AZ=�`|��ʝ`�qB���$��@G��U�u�����̎Mn��!��CqE�ڻ�>4{��ߧ �=%�-m<�ݨ��5��;�P�	�P���/�	�����K&�g���E��?���(�,eu��'h�m []W�+5	$�;����$ȟ{z���>R��]Á(���$tu��	���;�a��l��g)ͬ�=�КK���kN.x� �{N�6M���P�Κ,�_ǆ��Bj��|/�S��`rk׀J6i��Cx�����/�;��ݐ��i���K�E�%�?��f44w1�i��7gA*`��S�Sa����˜8h]G���K�c�����'#|����e;�fE�6яkG�M�U���u��)����6���Ġ���1&�&�������QѪݪ�=���|�#zu�3�uw��?'u������H�y�h����̒?Kห�������VX��J���fX���.�)t����y�"JV�-[-�-��8N�#�ǎ��q>Gb�Tu-����p��4E��9�sK�z�CZk6��ӿ/�W�p" ���[_�?��s��hK�^0�,��Nk"W���շe�џ2�$k�tI#� ���؅gG4�wY/��}"ǔI��0��?1�>ϡ���pW�P񜲱N}s�aj9J���W0�(L�$-�_���(�(�J����\B���/Nr�]��a;�.DFV�ZT4lrg�N���I��@/���C(����/����� b� 	:��;���E�#�<��d!���7�r�
T'�%��fU�:�Ll�}�g�T�X�̖��N��`)�_<R�:�1��Ĉ����, X�w����,9�t�D�%��r�l�^�X��݄������^�;�GcJ���[�r{�g-�D,1�G�B`+�a����/��+���_�d�W��@�s�(����:nj0�� H�]�D�7]�q�s��4��S��d�
N̻�Y��i��x���H]�����+�a����-��C��].w4D�2�������3fC!�[�'VtYb�t�L�>@�Y�{Y_?|x�}Y0S�U��/Y� �;����c�(�?FGUB�ɩi�dDs�YyD�]w�L�H���k�1�<=`�}N5K������l����.;ɽ�&w�.T� � G�=B����4����Yc5�Z�d`�z�Z ��H�ь�J�aWJg����uc<�˩���+/jv�ě�<!r�i)���1��$|e�lU:�\I֏|�=�6Դ��o�L���͐�V��Վ�
ɺi����{���")^rڪR(��9P���T}�X]�^�C��g\�6������h�pjJg5K��1�s4g����f)��6 �;�>���L�I�6�F�ۃ�~�$�����W���@��O��_����R�-����7�p|w�0;�r��֖�|�w.��n����tsI|�6��!m���`�L�ۊ�R��	ۺ�`�;H��?��V*�� Sl���*��R*<���`�8 U: }�H�.s��TR$�2��yAb��¢����~����W�r�_������e�.�B�Bm��/���,�*6	�xv�u��I�{�h� ���\�C��A):-Ln0ߞ�Π.�w����RIb�b��׬��Z�;��Y�H��D�̑��D���"v5w�VuD
�f��-��e�Ƅ��5�E�8%�
��I�}:���b��:���A��t"t��R��Df`�6Y��Ԇ��.���:�nI����� N�La��2.oj`�(g��A4 ś"��&PA9�v����lPl�okh���Zґ����w�(8�,��*�ȓ�(�A����Y��g ��x�0iH����ԣ8t�ة�QX����]ƕ񠰚ͷ(x��@,l�ur���G���T`jW'��I�W�������͜4��N�@j��r�`�H�>�ɀ�*1��3��e�*X/d�5l�Ңt�QwFڍ�����K����-��a�f.�-�5��ך��ԸXY{o��M�-7s�+�Y��t����{����� �v�c�)^koM/A�৳/������m-���|w�]��uX~2����-+�{˕��W	G��ҭ��G�9P,�E4��H�5�v��J��Rz��I׹?���E���X�v�8�=K�k�<O=ҐÚ=���\S~˽���B)���^O'Q��#�z��7� ��h�I:�\m��K��8��E���3N.=�M�bE=�C��0�y��-zn�&�e ��!I�L8��\���2��|ڣ�-b�ʾ}q�L����}�᲎`���*�S6R�6V��o�N;(>�?0��ӿ�[&��Je�oqK(���[��K�7�ża~ZIs�>N_��a���DS��֟"���m�s��aሗ�%�6}ק�5�=�B�g��h1��0Fì�)|{EE���(L�_8x�{��
����>���O�����][���P=ŀ]�5�2V���D\���Y��U�:�8�;�L�ŕ���axZՖ��b誾����Cxۋ�of��R���kP O��[�Eی5=��$/X��i�,�.��BW�����>��d6�d��O�يa_�L�@�\٤lP�3�VG�F��1�n
���w���LG�[@�.���MtK�����E�!5ª�q�����i�׋�vzOw+\2�ݭ`gYO��Y���K��'�ZHM,�,Ax���{%��n/�-x�t������|�x�O�T,��\N^��C�Lz�g
 Zɥɨ����I��A? r�9�/u{�h��Es.Fr�~]����Ϝ����[�ˢK?tF�4v��erEhWH`PS�UPn%Tզ4��p�8RN�<բ̆ΖO�3Fʾ��B�y��
��edjĮ�+
C�d)�|��K��a����ߋ�Z���,������<HR��Rw��&�?be����,K�@�T��X�_.��CD:�-~�c��Q��i蛰p{����CA��f�[� ^���5��}��g�UM�G�0cZ�2���}U��6:�A���]��%
:�����1��8O�F����hT�]�zT�G]�u����jF~+�`����ﶓ���a���B/(��`�(!\h���rڔ5�q��l��N�dnK,t�X��� �0�<�~�����2O�4'�!����!���<��U��z�⿢&�2� �5:�!	a�((2<t�(�F�����*�c�����W��:�:n�v�;IG�^h�(�AE�7�R!+���JV�`U�5��
����sY!���!�M�aL��v^$�MT�}��*H��5�v��6�x~��.�z^��]K[N�C1�/:,�E�igAW��+��%."@�4�@љ��=9D����ʴW&��s�H��R�%Ef��l��2 FP�0��Ng��`Q����@�r���n�`��Z�탳�ȴ�-�!84��T�Ѷɽ��VC����h�#�j,���Pe�͎!������ɪ�6�/�*W��7����n�8��hW��Ee�,O�4zF�y�0d��8�ݍ��*v�ʂf^�}��Kb����y�"��2Wr̅�E�4�.T�Ї�s���D��hB�v,���ƾ4�Ѵ������J���@�׬`,�{��(��(��m���}��vj��oHp��Br�;`\=�:=ޭ��5j5a���{����-|&!Pe��K?mԭ��ż���'2pg�;�H����C���<�n�m�@s.��t*�R�p�U�X�ܾ�����Ѿ�Q�yM	�2��l�lf�Ri���[=�W�������o�}J�s���������j	�PK���Y�@,��=��6AH�؊�����1�5P���
P��'M����w#�t��+�d<�&�4g&�	К��O�fY)R1l�G�v�A۰o|��ŉ�E*����q���g��u�{ȩ �y��a�X費-�����{���z�W6Сw�����k{�nuɖ����/��d�NKQ��{ -���dFuhT�K};I��:^��"|V�p��`�J��B�؄1�~R��^���PD4'O���P5]K�^�:.��i���	y;+���vA[2}e���AR;��f��+|�hqLT�O)Ro	�4-��/�GPϊ������B�i ���T�\�r��Xp�H�%R�mD�q�Z�x'�j�z�{8b\�q�r�7�R�.�ym��9����`�$�uF�1"W]��E�B�rQ�0ǔ��x<kG�kV��%�6a!;�G\�}��IZ�r����h�ͯ�f-�Vt��5��?l;����g���=^@��$͓A��N>����!4J�IV�8��΃�L�g��SQ/�Df��� ����e���܆�Ծn�˄�@E�E��>��}}BA	��4ApՎV��c/iX����dļ��Z
8eZ�T��Fhd�s)���@]��G��!���ۧ70dK�����Ե�G�4�KM��=ZT���1�>xP�F{���~N��L�9b�3-�=a�Ѩg�<b�;���W[���"���^�u.�+C�$���Ipl�o�z���P����M�&^��A��:M��~y÷�-���qf(Bv�z���9�4xs����x�h���@���B���"gr�����Co�Q��@���>tġ���,�F��z)Pל�`RTU��#4M���~O����R=S��4��;{�[�'As��zov�0�����|]&�1b��+4]�-�;A�ՐR^`��58��sڽ��� �T?��!���t<m��� >���z��/y�u���BJ?tb61,��?T��mR"�� ���ʹ����{u��s�?��~�ơچ8$=��(a�je������݋�&�c�K����E)�<���-^��k��ڐ��X.r�?'IUnN�zi��������B%K�z��E�ìYK�����b�����`�}��Ӻ Ĕ�D��v�#�hh�%~y�jG`����J;"Z�2���|3�\�jOwY�Fө92��v��8R��JsEe��HIY�w��Bĳ�4/��t�*��?�]��sF�{i���"���'����;i� �����Z��Q� �F�B��b�K������3��f�G0��,$�6���3`/_N&�*ع=�`
¯ԗ�az\{/�.���N`%�u58ò�>����g�I�Z�4BE5�����ψT}7�@4ZiJ��K���(�e��N� ���~��럭�)Z�%P�0Rk�u!����eF����ca"I=���r����5u�7����va�}ZH�@��f4��bcU�^�'s���zxJ�/p9������{'����Kx���*�tk̕�镄�0]�����V�u���N���2#(���2P�e��$pkJO���Y�Y�A�X�?� �x.ocI�@wpN܀���N�ڲaMQ�5	����.=��/��[�=�4��[�9R� by׷��C���RFZ&eҢ� ��{	��*ï���E�\q2����/�ls�4�S�Z:��c'[�>1�_I��ܧN�\vϮS��C(nl�7W�Y���{\��`���~��p�F7/�E�	"VwM�c4�Ac�	>��5�U��z�P�N��C��qW��%Q�SM�7��-��Ō��>F-:�y��2�Y�Cxp�k�P�7ɩ�૰E�h�=HP�-&6x�u���0P,��=~�/e&�����..��:��������u���^=8}<:��7�Ժ� M��&Ҷ�6d6gs���>
��|}����%X�R&FVM}�+&�OM �V���3���2����~x��ϷC���4��$�Z�mO\���U�{Sf�䘶e;!sZ�!��0����(��ъ�@@ۮ�WN�z�D^+���ڄJ�d�ī��5ӧ���FIw3v���	J��1��%B�*���7���wN��@� �G����AZ�U�öз�
�L���y4V�z,L�ރ2�3�@����u�*g���(��	�2���uZ:�@��3��N����d��T��m���CF�P���Zu���h$����!A���� ��@/��C���Ұ��M��.��?b��}����ټcJ
�x*�]�3M1�!e�����dx<��J��uS�z����NĞ�xdFS���<8O&�:2�xz����3ߤp�-�D�x3�QW���ބ��}�)O�o��u��>�L_#(}���Q��Q(	.�'��A�`���
�s<,�*��\�(��E�w���~��*�V�[�z���$V[�[�����8���Q��S �Dl�#)1�����g��7�\6}�bp�rU����Ҙ���L����a?8�j�������Q�H��5k%T��d�ڛ�*��']�P|&�R�<;V$�C�V�D��V�"��L��Gb�����},���^��6O�v��IƑ[u�~C���&�>Z����*R���r�IR�|����>����?�rh��w3��$7��2#kK����)�4�M�daX��W�)��AM���)��:.f�["�QDâ�/�˅�Z���]�/� 	Zh]ô��I����̼����#�"8R����K��V�w����^è~Ӻ7���p%��6��H��}D�z�4̅CJf���uⶉ�<��O'>�;D?�?2���9�I�[��7�a��Յ;��(��NJ��������n	EUс��i$��AJ�GP�QR���
�o��L�;u~Z"qm��؈�\"MP���M܎q�f�Mi�D��1hʿσ0��Dɜ� *8N���^<�Ӫ�V��8< ����F��w��e�5FM&;!YL��&�i�G�K����a_t����h��,��rTȴfh���?�#a���t�}�R�I�>�MJ��^��(�92*a}���#��gT���]��M�WBA���<�<�h�^G:q�?�$�T��P��X�P:�8���π���'~��<��7��SA�=/��x�ER�G�,���]��Oɾ�0��USC��bdw���
��u�-�G�&�O�m��Ӷ�f*�U��:�xNAq��,��m8U� l'��?0Y2H�Q::��g��̶����ax�� ��>�ai!���|��Dϑ���w