��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��e�ik3�������w$����g|��J^]ؽ�2h ^A ���'MJ�<����g&���c��VD��+�e�YV�i1!H%K� A��&���{��,Ê �|�T�G���t#k��ڢxt��=�%�ԗ��x��{]�^����{@X��Q����T���8�8��������	g�MN�s[��o��bR���Sv�$�52����K-2�,@�q�d��Yp�zM�Ɏ K���WP$�h��9B�2�����������\���b��Hڈ�n�B�����ڒ�m��<�Z�yO��d4�Ls��O?cEcrm^��ݷK�K�FWA5�u@��wQ�������XH�/ɮP72+uwE��k�pu��n5D�mή�V�D񤈅J����dB$�{���)�J?eۦ�K(K���C���1qpx�;�	k����d�����iZ��DF߭t\�����b��gs�/B����/�y�ڥ5O�g�O'*I�6�O$E�d8
(�V��G��h�k��݂ߠNa�_��o<CRw<Dk5��'hْR��N�x��;� �k�LN[���R�H�X�ֲ�:������1��%�H�H:1�i�G��Q�mQ㤿�ٴ,�X�(�z�Z{躯���0P�?�
�z"U��(����c/���p&c�����%���M�+��?;�R ���kq%+a��q�T��}�{�K��֜�=�юO���8����\vL�T�>kR��Mrq?j����Ø��=�I�ƕrzr&�qdA  ������b���v�;�eNø�CK(@�1�����p#Z�1%/�~p}��Jj?�2i��VK|@��V�k�#�dhq	�3䳠C�(�>6�V<Љc��z��{e#�JL��t�xp�ߝPP������Ԑ|7B�7�#��ʽ?z��R��.(�VY�
��N)JJ׾����Cǡ� �mt�9��a�jpcs�7;�YQ谤�����=9's�|vQ������˼���C���ӕj􃹍�A�7�e!�6+�K0�!�������v��L�c?�7b-$复�� ^_��DRT1眅y3�|"ĭ��5�do?T���,�'�Q #\��#y��
mL�4����4v�ᑀ�U�)���IqW #gK�|�c���G�RK�q1=I 
^R���H�}b��X�(��<��ٵԱ-�/��e ���#�r�'|���Ur-���E�� ɒƂ��ɌiU;�� f���S�d%V<��C��#�}��/ʥ8�0d����Ꮜ�h6���Ӷ6���[�9��4����3��6�I���a�tł�Э�h Aq0$x�"W���!_vi)R�S#K���]��B{��(���(��Gv):[Y8�n�L�t�tR�?;n=�`?��E��4��U�`�q���K���nK92��X�Q�<&b�Du�M_��0���姥�[Ec�v�1�;�� ��~�ʣ\ŵ��t���`�����K�k�,�$z�}	i٧�{Թ�����ɠN�&C����	�Y��_�CQkƄ�1�u@m��H�P�8ׄ�u�X�K4�L��ɽ�ch���t�O�M�dī�k��\h���n�������|Pώ�5�a��5N��@iTŌ�jl��ӵ�d�ts/���/��/���d̔s��>���!iS�md=ʸr�9*v�H]6�W�(�^ٷ�E�!^?kJ�i1��^���DMߐ��&#2 �l&(��H&J��G*��)r�au��ۂ_)��%�Hj6�[
u<[̕A"�0}��w�>	���w ^��uL��e��N���;�y�}�w��[`����M���8����Su��"�ڎ5��a��H�i���}�O������*ܙ��GT=ƪҹ�J��!��%r���7~z��*�Î�J���Jq���s��j��)�Ҥ�)";�L�s:�]G�w��U�ruO!Y�~T�M6E�M8�K�u~�5c� �B��"���������>ZɨP���̥�8!}�[�?������<��Ez�� � Ņ����ViR�s`��e^Q]�l�~�l�U��븥B_�Έ|El�֌�d/����'$�ߩ��bYZ�(� al��m<�Q��c��G5�G�K�}Rd_w
(��5�8�0��\o-�[���<;�iq�[nt�pQ�x�#��U���9�}�Ze���� �GN������D�_m -�lj9Z�� ����	�FV-C���ئ�8]h��/m�W�~��6`�kh��O��Y�l�S�$272����ݒ�?~�O�� ��;A�~�Ü]�m�7ND��-$�2\U(\�V>�k窡)<G�����V�Ы���1 ���m��q12Dὗ�K�� �A��'m�h������+�J��n �1X�4��67�٨�WX9nN�_'�	�� ����~M���2�s91���(¬�v,�	V�L�&��L����Jgz����ڗ�ɯ~PbCӐ�EV2S!z�Z3��("2o&F�D7$P�b��`�E��Ha����42��G���	��
����f���Y���S���/B�8�G�����x�a~�iv�)j��J�M`Ņ"�[�ÄG�9��	"�\,4XZ���}"�,[	]%�P=0W��0�;\��U�A��c� �c���S����x��)� k��D���)�#����W`�-����)lSks�z�q�V��D<J�y��Ԑ��>��}̸R}��MR��'حYB���S:/�;�1E������Y��BL�	 "^-�u����;կ5�Չì�+,�D�	��[Z��J�Y.�A~�q8'�5��)gyf8�$B��fUmy?��{�W{yp+M7>tb�M���Y�y/w�F��mZr��)���|(U�۠p������%d�ځv���Pn�����Ëk$a�D�عp.!f�%&4����q���;}�~D⮣$� ��&N�����֗i�:�
Yf=�Q|@�
�������a�V����=^�U��訔��0�۽j�Pq����r��>�Z�rBEl$F�=�MJ��V� @w;>v��W�g=.s��<�L��4�>dYG��y�s=u&�Eb��wo��֖��HcI)Fv=�8���zd b�ǨR^O����:7��[��h�KYl7�>�s`����p�R뮊&3����У������f?XR|�E��sV�U�ʬv�v��1�=7f�ŭZ���W�Zt2����sB���,n)��bzo\�D��w1I���跑�Mx�R�1��g�-�VP1��M���C�"�pݮ�}^�}A��� �i���������Zb��K�:ou�m������1ʹ;2C��k�^7�Ðj��n���_��1���%������XU>}{�,X�^*d�!p���u6��gn����Q�L�_&�2ʹ���"�H��#8���m{�<��#�p���J�~� �>���Jv|�C���c[�B���o뼯���F<��r�yj��k5�� ʩ�\�y�X�l2/s"��<l�j>t��A���y@���b���(�Y 6�8���s��[�vd�̂�o��-���}Lu�!�	XO��b��`d|a��G���D����u�ۙ�t4�,���2cy�hؼ�`bf�y������W ˒̇p����$9J����@�ƀ �Y��_'�/tYm��x����nb��G�]ޫ*X�㛕�]8�:{TG�C�@{~a7$)��i��#����֎[��]_n�d��)5Y�+�v.}b�4Fr�(��dah�t��I8=���dJkY�z7��D�NA'�����P����7Z�V{F��`7��d_N~s�*p��h�ަ_�M��^���������D�ɔ𴓗?2g(=���uѢ>�O�qE��m�{�?ϰ����x��7�.�m�"��i�XXeC:_JP�F�(�ự�3��,,]�X�+@�'�)zu���+��06���:7U
�e����|=����t%ah���g�|B���c*�;W\1��g��puA�ͧ�q���!���l��a&⭁_	|e[p7z@]�v(�Or!V�
��C*g~c^Wϙ�L0���dV��4Ȃ����`Q�'է~S��S?w�i�t�Z�˪+�#����}�鏓r>��]Na�j��G�A�HٗM���_:��dhnd%����2b�m�8��!�j+~  t�c�;y	]M�ӭӭ˸M�+���W�"B}�1A�%�s�v(c�p+����M���Ak��3��ܼ��L�Z�%�K�B�r|�@Fk�r�aI!uqhU��at�`F_g����9$Iƫ7�?�����_�h�rI���90�����с�����Ё��p���V�gX�Y��W������}�B�G%��tg2�FQE ��s)�����e��]���YsPfb�������0\���[u�{��``k�g�#- >PE�v*��%V��ɗ#�x������{�߱y�^Y1v���w�zŌzũ�Zp!`���`�z�+��K�p�S��I����s�15��]�/�?�kr%�A����zN�v�{���� ��w�	o7�@�@�Ȯr`��d��Ǭy+��z�Ɉ+i�>�f�A7!
���1J�?�P�P�]�2؅	EC���CK-���#��n�'��[*Q���+`�H��"���68��E����{��@���n	8c�J_<�|��%H�#7�������mM�t�t^D���	�[�j���T˸9Y��h�f������=�S��g��@���� 7���ޙ�ntg�S}�����I��/�1����Oo���r�c���n��䉹S�L#.��`�M܋��o�*o3� ���lQ��σˏ�ϓ�V�Ɉ�]��&���I�C;n�U��k6pq>-j��T����E����tBX́��&I�>��f�W�.���1y�nľ!��	�b*��J۩��ڡ@��j���cԌ��?��&:��>��I�o8��~4�5�����:(�����xZ��Uu�)4l��M,�wG��0S���T�oj2yqX���}I�h#��Jlf϶�/��mau$=��/��K��(��?�-Y�Q������U2���u��{�Ɔ� ��*E�1�j[�7q�O�[O����G���Q��ƍF�3T&��x�=5��Ds���^ܺ���I ���d9��LؿAU�	Z���-�OWO��t�4܉z}���v��Nm����Y3"_��#f��ɻt4=��SO`#"�.2阅#�5_.�g�-!vx�c)$)9#U�{��p��x�g��(�p�*�A�^6~�m����v*Pك2e��"��5�K�SZSW�Bh�z:���n���������
��_���񊈁�a�GzZL�X��
�x�ˠ�;���Lׂ|).�Yh�3NlY��{�(�Ə%�>l��?�Ų|l�Z��L�n�k3�����Th�x��AجQ�AYS�ޖ��4"4Ԭ� 	�+Yv���a�p���f-5�
l�%�"�{���v�H'�k\��	>�E=О�,�iV�EƔ�e���0����˒�widL5
;3�Y�p{1�Ԉ3^k� pU�.|Ċj9�>��ý�f��R���x)�lU/*����hU�ǉO�ն���u����h��U^�}Տ����b�R���!��E�e_���R��Q���CqH/{�� ��_#�ؑ1��yk����Z���!��L%~�#���d�"U�F��'� ���a*�Y���\ D2/����MI�``{�9��?�"l�s�v&��&rc���=�;�6�BA�!%'b��3�B��RZ��������W"s)�r;��=�[U�&�������	�����Bp�"ܦ>-KDH�c03�6b�~�����*=u������FQ��e�[?ь��,�j[�|���a� ����_s�~fϔ�,�h,M�v)$W\חb"݀e�{K�y��u��g��9R��c���@��*k�Q?�1� ��+0���<w����ͭ���䎙"�i�JO�
$���pgԬ]��W8z�����?�
�8B���Wd �;_�R˕����(�Nv
ZmA�i�&�ub�ށ`4n�g�>�:)(�=k*��
�A���v}��t&�&�)0�1σ�(�'��s����!P����g���d��u��W�E��,_%�ʸ?�3����Kt�sF�������A��	��ɹ�\;j�ϠQ#�����[���6��j �����n��2	nUHS\�G�s09�r�D'8�s@=��*�;P%Oݚ���շi�������3��;�K|�A�`Ht8�"	Y��g�^���FP*DEm�ص�'���ν�Lr���O8��I�#��k��bl��{6 y1h),Q2��ɜ��8`�=$��h ���~4��6�8���J0�p�D����?�>Q�R'��/_�Y�kýn�$0�Lsh�/�k�=���x�Wza����K��@B�)��w�=�@A�B�M���U��w����!�2vI���i�jV��5+Oh꼉e]�ў"1Z.�
�~��	'a6��ėL4��B^���㛱@�m��5�w���2�u�!t/=�hّ?w�(�2H�)ڍ����I����կ��E#�㾻�/8��nժ������{���-�-�򈯜DcX=�x���΃*��I@c���z�$Y�CQ?5��}���CBfƒ�ó󞊔�(�q�/l)�{��&,�����[�E�}?�M���Q#�@f{��6���߀�"?�0�������%/��ۃ�T�e*�C'lIaU��|��ܘ��|3P��K��o4E�J�*��&�%�3<����/QE^�9e�ޏ:L�9^��n=��R�#v #�B�9���6�K�0���<������՛���K�ۋ�	�UK�v�ڝ����=1�_��jVǶ&���5�oxH����
�k}���}��i�x.����=�r��a��leR�h�ఌ���e�{���,�v�z�u2�m�7[�g�Hc�0H�wg������ˬt���~:�o���IM�K��9�u��vA��S��mxX���\�Ĝ���}=>*��3�#�٪Yt��9=i���?§�Ba���B
���K��]=�4�x�xk������0}*��x�I�����8��<�]1�9��!E�Zq�����.�ݩ�R,��g��E4�m���wn���(�[�pRm*#�SK>;��I�D���͐}�� �