��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY[U4\}�(`aL�ܬ`PT���I��\I-|p?WR�K+\]R}�SVI+%��F�7����^5t�݊�F�����*��R�)}�Ѭ��[T�g.
WiC���wΧ���_�E��:'�ɾJ��Y>E�B_�̒����.ݱZ�?���cҨ�J�*>>}�H���D!���&�Mx�$%�����!$�I�W?\�W6V��Ux�U֢�g)��rX��ԯ&�P�cƌ���{��P�Ȫ�zPcYU�³��{�*W�Yb&z����0m9Q��S��OVf�}4]K�$���5�x�h�j�=|��U'����g�Hӽ���ܠ�	f|{���4���b�e�~I��T?��D������0^�ϭ\���p�5ߗ\%)*�����@�$�e�� y92��Bl���vBA�/�C�m�'i3�L;�Ǖ^LD���=��}��ֵ�a.Z�����$hgu ���|�\d�\��8˾�D����q/]%�@���{�Y�71������Xk���Vd���Sb'7&%�(���m���n�/�9��G)n����a�W����i�}S�du��pb��1��6�b�F�I�[.�g�q-%�<��E28�
yq�)<�?��C���!zE$�.��r$.��\�r�{���	�����w{���h/�i�Ox�E�`gsd��a�^)�*�qEȁ��}r�r����j��_�;��nS�R���w�	b%+��s{��t����ύ��������C����3�+#�Y�� XEp�zӵ~���8$����&���2�@U9�#[���`~^��aQJ.Nޏ��	�j-���b����vl.�X�0����͛ �!�,mXk|�������EO":�V�1�1���}O�|zdfH̰�\�>}5G ;P�F1���o����ke��MxPV�*�&��4�Jix����$+P쌾Я`�C�E�������<�D$�R��x40I�)����a���ߺ���`�����)�]�hȕa͔DA ��H�eɴ�;����}ķ��G;��u�j/]Ľ/����)�7e�_����1�XS;��Z��b�r)�jA�t�c+�o#�EdZ����~���ueO�p�h������X�!:�vZ�I�a���O�bD�H�a�,��`B�#in5�8�6n��Q�J-��%)m����`��joi.-�h�:���W���zd;N��q��w`�"�~�o���rT�PA%"����vMb4�Y�0�co�8���Y�UC�6�H�h�q����ۡ�?%��67�ϋ�Z��蕑J��,h�N���>�ht������! YU)�趹{��kP��+ 7���4Y
��/x{2�v��E�,;�Bq���I}J��/k\��Q�P���=Q�c2�(8�҅BD&M
d?-{H9�p,�j�iÖ�vA��?!�%H��C��:�� �٫fu���p0
H$n�Ak)ݛ�Z�{�'H�;~㧪�mG�p��/�6s�ƼHԚ� bM7!	?�=gwy�}	�&c��>�&��?�witMQYZ��\&�b �Qa�PF2d7&Ո���e?/B�Q@�.��7��K�.��N�}��n�_���S���9�E�ڵ[���0Q:R���z�u2p*�[ұV�ruq?�LmRf����OZE�%�U!P�P��<4����jU���j[�h����~LZ�����_��ˌ L�W��oܸ|���6���W�cOtL"@pn��t��������OԳ �OxqOEUɜÞ� :}��*���Y3���.3��<;����UWoX_���=u��S�+	���y�761]F�^���n`ܙ�a���"xs#o�L#ө�6:h1	q��e�!vr�'yJ�D�Q�t����Z�@�F"\C��ʞ�{cl���MPع!�z�����:h��,iT6���S�����?$�G �p$�e��#�w�3iM���:��Wj#�jt~*�,��줕����Y��,@�,$�ի��r�W$i�a�Y����
��FݥT�<t���79��#���e��q�FՅ�wXF:�0;�x;F����|�[��0�5mۻ%�0ןf��s������#G�#I	�?͐�͹ ���B������8@�N�@��~�>����H�"qC�ē����Rdb�r����&��) �lNU�ڱIn��.��8��T��Gy2�������~�,Hg�D��U��Z��y �Ef�~��aF-�+��w!y�z�0��TF�XU���_�Na�"���YaF�n3[fi�k����q�<P�����|4�pZn��Xu�Mq-�A��]�F�m#zr�@l�۞p ?Q��$���5-d`������n)��rڹ8�޹OC��5kA�c�;Q�i���⦞�8���7��>�G(��ѩ�>�����@	g���� �x�km�Ik�.�-wHaLU%N�@�s�1/P)���r���*.xq�C�y�e�)�W�֫�1o���H&�^���ƌ�-V��<t��W�2�5r��i'x��xRN׿v~)X�Izl�5dMU�2���=�'�9�y�X�췼��h���Vi����6xE�n�!�,��Y��ؚɓ��&�Ĭ)+ �@�dCdT��A���S�(����a%@8JHqb����q�r��T��X���zK�J�9TZx�3������Ο��z/ߎte�Z�ع���n�?�q�	�o�l
օL�ͺ5n>�4�tzc!�|���V`�4 �?��~�dLE��hEs�K����*���\."�K�b�P+�ӆ)�#�N����RXY�nw�V��*�2&WpD�^T����(�I)��a^K�ba_G}�����rI"�z���99m�@��4Pq���:`2v"�Ь|7�KV�/�t:����q[v�3�9���܄!T06`%�A��+���K?��/4^�uV]V�=���]H��oP_J���${�+_����co~7�����`��J#OL9�
�(�<��6"CH8&6k�_�|�҄����|���~W\<uqC��Ҁw�}���@�,3�~%�k|�&,-�l�{W�j�Xp�؋(A0hd�y�1�¢sF!b���&��� ��GYje�ƏE~Q^�A�i��B�F����:R��|����kz���G�/��eB��^��	�)�9C�2=XRD��(���y?[\���L����op,c��`��f�v�7�#B 2�6R��ѩw,A ���Kk:@(��pw�>��;	�������aO/ �\��vZ
dnӧ��;�&�k��ٱ#f�@���ox�5^����#էb,�W�DD��0�b����ݙ�.}
�#�\�8���q���}��]¦+1	;�Y���3�#�4�ќ���7��fR�B��</PR�ua@�C, Q�B�񾄕UB��/t's����Fz"S�ې��)"�Z7��0�a#��ޓ-��GA�Rh���TԼ]�Щ�`�h|sc��)�<F�iw����"����x	����eX4��Z7#iuY���G�,�u]o���\"���VM)D�ҿ�o�]��jk_F��my��u.l׋;�N���n�q[�o �m���������˴�W��QF�g��r�� G���T�5���E)8����36l�#3���� 료�춁�B�LGb��T���*�2�ւ�|]Wb��V��q��[�4�Ԛ�K ۤ��������|�W��OQag��
��ו3��%S�p<;F���:Xo ��S����av�_TTn��1/N�sJOy��%>^Q������#T;�tM�)�?tʤ	��| m?Z�c�Nw�]�S�p0ط�5�N�	]�փ_��۳�V��}��կ����3����M���c ��2� 	�F4V/=��ۛ�'��|�н%�[St���F4���@E�1T���f��p����v�>�ncǑ�͹���pI�
� �����u��>���3�t|�TD�L�{�rwM' ��4.�Ea�"`5�ό8חfK󠟎c�#l�`����Z�o!�T���f³2w�0�m���̓��c��Z�F��V7ܵ�k��]��ۂ�4� 'x}�P)`9���7��Y���Yy@���6^릻� }���>��4����@>H%�+�`��T�,
�̱@�+}]fQB���(B=c�q�ޡ��)�k����N�Wt<�ŉ�o�_�f\���.n���ŋ��z!}�`�	�j��f;�����(8�^yؑ�;���s��0�HS�4"�!�&OO˺�n�v��>)�W�򱖠��=�2�^�ˇD:�#3��/s3ĝ3��N׍{�w�Q����cK���R��6�#�7�%w�=o�ʺ�#��<�ͮ����i�W�'���#q^�,� �˽+o��1�S��^�9���� t�P��v*�	�y�=jG����%�9�%���/����P �_��ٟj
 ��'���R�u$w���ײ`�9"ȩa5~K��V��I�L�T�+��\�c�W����i�-��1�T�u6ڜ�+���O���֠��;�!�Ŕ�{���>�F~gO�J5�rB�3������/�v~MY����9�xd��,	����\�=�5�	q�����Ov�^	���b.#��A��@�ğ҇&��<�;F
�M�E�L�[���}eDEJn/�.��ԋ�`l-�������Ah��qX���,�`��X2X��p�A��?��H����7? ďɾ"J+���x�c�۸�I�D1V�\��T|�q�����NK7Ԧ�����!��%�^G�@6YI
[.�[K|�D(�C*�iOƳ��=?AЄa����1�a2���*���|g ���+zN���s��0Z���-�=������<T����oT?�N�K�M�օ%zz,hj4ɷ$�o����G`��@�����
-ֆ�N�EM��6�e�<���>Z��	)=��nI�X+g�C��݌Ȏ+�O�gcL�Ǫ�d�s�Ŀ��-?M�!��m��;�/���J��+M�T>�[�櫮ꁃ�#/����8qi�����퓨�j7����"��k/����e��%���y�����W�v>4�ASM �¬�fs��U�-��	�h��`�,�V�7k�7C�"�;�X�8��/���=Xk�Z��B��u"�E���X��Xa7�Q b�>��Vo:�'@���SА���<_(Y�G?m�^m�Q/�O��60b��G#I_fL���.C�d}`��};���S�	B�;�16�*6C�Q���Pwדi�8]�}�A��N��/�T����H�N�3���Ef��Ly�q��2ܑ4Bf��HyL	�#�����5I�\����Tb�(�/�GU�~���+�.r&EQ,ċ�' �B�"��rL�	o0[<��V��w�룭��^��D�H����n�2�H�漩�h���i߄��4�7hT5����tB[�d⪻J��3�0�DC��g�k�֙,~�	�:��T���4?���h�����(0�ZD=4B���`|�����Fׅ��q,|�A�G��ۃ쑅�Z��N�Pڪd��q��`�����o��[t�C��kXb��� �K�ʹ��s��a�=~��a@.e&����#����l;�ͨ��9Ka�S�;�C�k2�Iwz�\1��m�p6�;���3��"�9�c�cgy�dG[���O��MAb��W90-&�I��>D8�?�d�%�@S���P���gl4��	��a/��Ӭ���2�E���w��G�����W�"Å�Җs�ٓ���CY�s:
�rô]����#�V�r��gc��>�F��ؚ�����{��cSi���>=���ȫ�WH�Y6,\�"�TF��Y\3���c=%���R�������+Pl���@��:>�G��ݤx1�7��zяu�9j���t�;R���-L��ta�.��"߲�6# �L��A޾���n�%i���Z���L�G����-L=��w'���,�̮(�T:i��X`Q"i�ٽAQ������`P�W�O��H1u���ۮ���ʴF�*r.2=�8��cSw�ʖ�ٿ빖-���i�buⲡ,�E�S�O.��ʉ<��S�x����hw����A
\�^��b����W@oA(�:Z��1J���vn��Y��eHQ�*��kS�:�w��s�}�����~�á��К�Af�WZ���py���e)wc����q�G)W�
����V�t4S�bY�m���k��޶*�|!F'�%�����( £J����eȿ��g�wrO@z9d���t�@Ю//�����Q�v����%�������k"�f���q�Q��ד_L?7߆�� �jU�qT/�Z�T.� z�n���0F�c��)k�niy�ͽ��[CP��JW�rl��[H�3���%'E���}���u�Y�054R�m�)D��ٟ7 �}d���4��S�����j���Ӭ�VF��3/��+�̉�]o�.q���n�~A�q߹)�tx���s8�����NbN�qK��<��8|���h��@���,��N���`At@8����ә���и���m#��K+�����ۜ�6:<o�ɨ���en�>9�硩^���sxG$%��VG�r�>H�iB�]s�&*��kM%����RF#(�t�a�~D�95�Q�g��P4>Y�V�\���\��wP�|j�n�9�(�J�E�����N�(�B(��(�*	�7��;(�lt4J'h%���y*�8�@b���F�k63�>Q�}B�z��ۻ�,������vϴ6�ƈ�б�ã�JS�j4x:�\k/�Ld����JhlE"�Z��%]���5Z*�Fr�-sP���-˓<1���%���ç�p,�P3U�Nvӄ����|���qɪ�<N��߶�z�F�G�i�K�]��.�W��X}���3n��.,�j?��g뗅�T�X�r�sf�Z:Q��7�Z;?��o�q<L�Ec-�3��~"��;C�32�z.��[v�W��ާ`���Ͱ���"�(F	mCcG4x19q�Ο�a��� ���ڳ�þ��Q�_��5B=Ԟ�6g����W�g�F�����`5]�������&n��"�V�Ř2�.h�շH��H��D҉˫�c2:[&��&1�d��P��[A=%9�= 蜟@a��������?#����T>�բ�"�.SVt�׈�L�\����	�.z���h���ɬ�����������u8��ҏe�h2�n�p����m�i�V��Jvs��y.{w�E���Ӡ����߲jjѺg{�>��.�E{᭘�`�)�\�$y4t>��7����}2;�]}g0RJ�L0�"}n`ZX�GoE	et@!E��4�|�gJH�uԑ���#L�W��0]� P֫(SM��6��R�h�~d��6�0�eᲾ�f��>p�Ⱥ(�	g^v?��1�c5탿*e�ʄ��� %��G�lj6����07*Kۮ8r ,����!v齋gD�3�.�����"(�S�Ck�T�KÒ�4К�CSbD�\2-�����:��X&�a��քE�RˠO鯗e�q_(򰣓5���,�y���xu�4gT���!�UQ�,�:�$���c��1��8 �#fE}�^���q�זa����Q���#X$���$qZY]XJ�X<�\�Z�%��k2�}g���L ��]����-E��D����M+�Z�&b�*%�̹|�}�](����7?R�����u�����(҅�5��O����Jq��%mBS��Bt'�557�K�vv�>ܯ����ԋ ���_I4�Q�5�:z���w�@$ccߤe� �������9;]U���*�g���pqb[	�+4Z�9JHQ5�]�L�ES�\�ɚ��K��3� N��ɬ���)�� h���r'�=��2x�HSE�t.^g��8�z[�ؓH��W�"Y���~=�jTLڔ}8+hZ�2��*����F��
>�7���}�!�;ξ^Z��C�G6���!���e���2�ïqI�Vj»"KF�鸉wy*4>'��.�K[	u\m[�eLGs�# �	$���E�y���S��q��S&�E�n0��;2�a)��� �B��|�ăz���%H.r�8�$~T%���Js���m�b�}u�Q� t9�@��(P�P���2�K©ם#�'=Jdz��@I�p�&��W�58S�G�����ښ�"�(��a�`0"�o}� s6{��	%�~�[Ńtu.v+�hk!BK�`�W����ߋ���hr�
�JL����8�ؕ�u�Ǯg�hM"��F!8�(�K�*��Eq��,`�W3�k� bO�Ed�9 ߥ�O��iF4�?���9��U�.���zPK.T��ô�*D���Ԃ5�f�9F4�6Us#�=zv������_$��2��U�LG�n��w�A�@~~�g�$mFDO}��h���qT�U�KUm2��d�a���ϫ�ʯ�ӱ�ߛ;�3�.I�ZS���Ml�����թ?;h���ߴ���v^j�eT�_����-;�Q_��gu��q�'��E{�6�x�H�a�����(��j�����K��1�ݶ5�/������%�7~C]cJ�|!jkB��5�&��.+�P,����x?�΃�� �S�g�	|6���/��A�b+-x;���{(&T����"�"&��o�;VA�%  �,)��Ie�Z�7����r�Vg$�j 	�����S����l�R��r��]�~ˮ��`_��/z�'x��X<�?�0}��h����D�t��}�5q/ɒ�R[d4�Nl�є`