��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VYjf�>ρ�f`+?�H����tZ.ɍ�g�9�>T��������������e�똬@��h#uyN$fq�fa����Jwe0/VZ�
�F��;�d�l�H�K˃gɩ��!J��.ք�������ǡ6S�gA�,��>�u�b�}	����P��d����^JΉ!�?x����صkz���\ B���ݰ�sf�KE.R�q�fL�C~���5��oG�<�+�X��8�v@9�%|��$r�N��@m����>����b��-u��J����2���f|�c��Ӹ��e��>S�:��,���胪�ů��n���1��ݍ��%�\�ɜ�{��frPȸ�:wOs���1V���bC� �GG��B�!QM��N��RQ�Be�(�s��O��s�)n����)y�ǟ�e t��Vv'%`!�Y����xU�4R�^v0�N�>�!�Gҟ0�Տ�Gy�A����YT����Ky�ɠO��b
MZm1[���I���M&�E߸�cG����� ��?)}����7�����\�-T���W;\�s��P��:�BYqc�?b��YY�4��]��q��Ӓ��2��j����3q�:����+bzR�p��$K
��㟡����*�C�` H��$��UDė��mq�}��s�Fs}���w���~��\2ǹ�l�p!]�����N/�)N������"� %��q$�򈂖.%}��PB��"����21�π� �,��PpLlC[�2�"�#RH i��+����Ѻ���0���$���r~�m&JJ����h_��݌�R�� b�Gfl���
��*K#����e[�L<u�A��vFg�7��TV�N;M���ܵ�a9D_pb惙��1ܲ��	��/�3�ɖ|G���Ӎ_�;O��F�SP��9�vD��#�ض�AW�#JM����T�uBXQb,�)����{T��S�{+kE�x�1`J��/���&�"|R�u\�&�0^]�a��ϧC�~?�'��sg�,��i=�,�%:���)�]'�X������&!��{��N��䁣�!��^:�֡m ��I��T��i$��{�:5���'ܮ�����kV��~G�ڃ8�0&�$�QtP��a��$�.&������t
���3��^K��}`�i^�sO�h�`��7B��Ie2킮B ���wRn�`>S�57$Zp��z��f��
&��0(�zI`t����;��ԕf���	HZ���K@�,^��� GNع��2M`Nߒ���B����é����q�,�(9^��(�ֈ�Y�Y��ٿ0O1#��.X}|%�+l��w�T��e�Z,E��9w'�Kko8��^��PA���3T�uq!�k�I�kKi7��IS�/�k��|�n�sޢbq@�<+���ib`�R����:��'1�4u/X��s�iݗ,_��=��/�L6���[y�Ԏ��QR�}	A$������r#��# �*U�[C�+|��ra�Y�O^�X���Q�9�����ZW�^{��Z���힗���T�[��oWa��wg�����RY��	�|���X��nC����fa�Q3c6�'�B�9�N���Kᙒ�z[�ӏ@��1����Cn��t��
?�C�D.��I���42���\�c���1	S�XC�J||�g4c~HFǸ���� � C������Z�OQSWzf�DS:)r@x�n�^��.�Gs�f���R��嘸�����<��D|w\��B���7�M�\��,�g�#;H!$vk��}�e|?D}�b1c�Q�q`@iso�vE�� ;��)j��G@�4Ȭ:�%]*_J1/�Q�h���Q� �^ҷ����-��
���<q���p���*p��];Տ�)g�\&n_E�K#��u-8�����VAO>��e@p�;-H�t����LTصDsvn©)�{7�R�p���7��Jo���Sǎ�
B"�W�ܝʖ�p}�{?��t2��W+�����9m%�G�{����P'����a�쨰����(fz�\w��>3�ʚ{���,�~��<3�+�;�ܘz�o!�� �92�o�d�B�V1��]$�K�g�k�˻��������qm��V i�里|q|�0L"vT��)��fڠos��Pl�+�N<��?f�b�Xa�"�O��O.��F��Y`��+�\Q�SJ���χ����W)�h�u<<b��c�ޭڦ�}�2����mh�.q�> �?��%��'V���S�U3������g�ۨ���.&���p�H�u(`�y��d�tT[5�|�H��fc�$F�ڙ�8G��ڞo�f��b�\�g��Ec��>Z��L�:�)�\�Ϭ̛m�M>���'�����C����3�#�"L`ϱ*%_�0��	��Je���w�����8�:S�e��LG1����3h�=�0����.]^�l�thk�r9����rkyy�{|�Iӳ2ԭ�l
sgT b��{I�}��]ƤP/�c��M_e�9��U�%�t`lH:j�Gqwئ��.�L01����9�-�xU?l�
��}2�<�JzXV��g)�O'jp�➜J<��<?p���󼴢��'��۰(�Es�1�(KQ&lJ��AE�MjB"e����� �V���N��)�2֙�FU~+�E��%�x|Ԩ:��XS����0���\l�T�F±L��X�+q*�(5����xg�M����v��{±V�o�?k�3:&ف�=��GH�d ��;�C�{?b�[�e�	�5nb�mB��Ӛ�A<�x��J�'*���?L	�zvJ���$��h��Lc�s-���ا��ԙ�[�b�>��+97����hsX�8k0��濑m����h�\��5THz�����4����dQW[s�G_�R�خϣ�m*� 7���,��
Y06�RTuQ���G�z��D2�@�7(M;jǜG1��Hj�H+�	�H�J�2�&���fm�JR��1��<����B�;9{�Q�n���~��d�%UQϸ��~��V�n�q^���:@��	�N����ήfaP�3�'��%	-�\��U���R����W�����`ݤy��>՗lnv��暚e�y�4�i��J9W����U涏Fݵۛ׸�� �%���M�bӬE�>�ڈ�hy�QG��cwUm5=��AW��,���^��%K�z4P�m���m?}�IG�z\0c����m{Zs�c�5P1���ԓw���g�	�)z�ףN�Y&�����J�_�y�j"!s5����!�_��?��eEj�)��)��\�0���v�l�\+������k�U:ّ�^�4�n�dQ�k�$�NW�
f�|'���R�Ζͯg��P��W��]�>ɔ"tF��q�)/�^F���Q��E`Cz���H_?���O�7FK�cf�@Zú�=�1_�d�#˜������l��=ՂI-����e��mE�j˗�&
������gp���7��;��
��^��=�*6S�BmP�Y
����d��5e�PG��fx�&'�Wn���G�.�d!}l�*�v{��A�l�	3�V(�'!4����Ф�;7)��fa���{��Qp �S@��Eس^w��j��-��ܤ�,��-s�y��ˈ]��ɀ"��5+�-ov��	�#e��Ru���I�{p�n�"��ժ�/�?]C��Sb�Y�"O��ek���|��x>%�9���e��>�Qq?����4��qX]n��n�#��Xy��C!8��q��m�	,M-���ZY43��4�k	�Ǩ�&�2�q�
eFlx���c=��bWeJq�Y�>�Z[K|3]@ok��Z�"�F��A�N��z-�i;�Jy�A%�GfT�"�*�����=�٥����S�����6D��eL}"#�ܳBFԻH�b�{5#���!tk���_�� �+��7� ӝ�s�:q�C+K�㱞��0<�&껒_$d0T4/��=c��ր���C���A�C��_���4�5�W�J��r�Z�.��'ț��B��a^T��������%��������a��Ñ������N �:���|�������ȅ*�y~w��
��KQyz�5��]�tL_���ު�Lɷ�u}�f�����K�r${��6q���#>o�+�Z��(#c����T=ᄵxr�%�пV�7;�٧x�p�>�d��k@��7���6�r���=��Ʉ�^�c�ØƇ P1�Jf���M���̍S�!����y(��# ����OY-�Ԥl(�;'�@G��w��tD�$�]/�?2 e����ɫw�|��Z�:��?��/qꂖ-L>3~}���e�L]ޛP'�.-�����d�#�YiyVX�q�bI��
�n;��W���
�*�_��-{kϞA��j���H��>�HXiR�0����f�����)5�(�+\GŢ�/t��T����x@����(�]�a�^����t��'%u3͠����aK�_i��p��^v�e{Ǔ
�����.�����Kq���U���o˕P�h� ,�o���8�sN�4��u����(��S%>L�'/�=�^a���B�1�'�1��c�$���K>4GE_b��Az!���/)�N���+�_ڸ.��
K�^t��T�����܃�s�}��V������A׮/>�9/�Ӎ���l,�vhK�*=�	�n:\�s:H���n����	MJG�σM$+tf�u B3�
-P/!�w��g� w�َ0��p;�O�֫��T���9��FC-W$,���[�	ϑS�8)Q��	��G:��YF�"����B���!˃$�v��;����3c	�>5Ls��H_+��m�v�Sg���e�2��r*���;g�jX�dE��@(��)g��W82�x�$��HE1�����/�v��L�U�D�tc�>���ٵBϢ�Q3���$��ɇ�R���h��qr�v����B�}L�� ��������@����X8KO� =�`y�E!s�� ��~�"��g�$I��z�Ў1Q8��>���w�ٲ�8l��͓���(�_���&��(�p��5����=�.�� M䁶���ݙ�����Y��/��v�ë����Q���|� u���4*B��3P��������c���{���bP�Cȉ��C1�͸�q��<�I���7����~P~etl@������B�R���w�)��ˠyf`d��yK� ����4�Ӈ鲁V8�X�-Q�Kbkm�~+{�>ZZ|����t*��|;��n[�(lf�kC5U�����k��y����lVD��/'%[t�������I��~8�7��W'P��пb(w/S�2���'��%Y2ԥ�ׁ�&��ŷ+˝��!?N
=I~m�tPW6.�s�;�|U�����@��`�b2$a)GӅ�Q�r�nc��]����*�@�ĕ�n�!�md纠�8c�b#��!id��K6n��"%�$������G�p�2���(oPI��["���� E�B��-j�W�OL��eqh�v�q�,wE�qW��`<u�d7���fo�d �/�xl���5�����H���h��$��2�<�:�
��{�'�ͦ{�q& ��l�"����ۻ��Yt%��·+r=Y������;[}��`B�?�7�4�h5>���nf{!|n�*���-G!"V���ܬ�a��}ë.ve��� i��_C3B��s��WȢ�XLE�M�?����`��QHߨ�I�CJ�O��g9PX=��;S�*!��@�+ɦ�f�\��5����Q��� /��WD]@�d�A�O��B=�ܴ�Л#B���`�4���MIi�Щ�����m�����������-��W�l;�?XfL����u�C.Xyn��o���*���W��^4�O`b�*�05Y/^���+���G�H��D�Y�,X�B�i���.��JD7����1ue��䵺}�RY��� �8������|�e�կ��
�K��|��p+XI\&�ei�u��f$X��]%�����ua��37�kPTm�X��{��D�$[^�y!w�_,��G`\ri&b����m��od�-��yyup�����:Ek���ñ,�/܆̵�ԕ����{�n��7+��RV}V�F��м	�5s�����n4��p2�^��'����J�-�V,�Tt/��"�M�&�"t��{�]V��2\~�]p��1ag!��v�9�γ�!��)#M����řsV4~��"'�@Z'�[^R���h��eG�)#8&S}6�
�[w�<.��~�RI�C[�Iu�P~�x*�*<�%��py��S�#���#H+�1�7]����JRx>	���L��=�h$GX{�T�QUQB��T�=�]�P�BOf�	?��, S�t4#�g;w���6�t��?a�čNp@o}A��|~ZL<�k�"�D�~$�"cyr㹰�ֳ.��n�=��DM9���5hZ1�G�1d��G3��J�PKdf���>vJl��}s��z���f��,��[��'��"B,�큼�JIT��@��H�
omwR~?���:���:<Y�s��*N�{��N�F��7[*��t%���PBh��7pXVϩ��0��v;�-h���yWF[;J���JH8+c��cٮ�h�y�l�(
桓��+|D{
>N,�N%�����i�c��.���������bb(	���߻���3���X��[4�$�|�7D�cwe�M��:G��z��Y����!��&�1��"�y޹u5Z�<�<F��'�?l{�?3�cV�����_	��YW/E��v*~C���C�(ʚ��]����|Ji8ZO4gt~�<�������K��z�(��@R�3p��M]8�qm({`���!}�lo!"͓ǫ����Q�:��xW抾�v�y��vc3g�i�r��R�74�e�V��2BUq�[�� ?()ɢ��|�ܽ�'�0�Qߩ���H��k��{�_�W�z,:8˜9�I�W���c��\�=�XܧY��7��<��X�/)R�������Ï'0��< �]!�t�R�6��}f��� ����,��}��vxC��G�tg� ���
	���O�G1�;��ˀ=V��� .��E�y�Nw��UT~ O�Pc-F���~�<�v�v�6d��'|=�H�`���B��P��}��/8����,��lID�V�a5E�m���(�c��>iOF�-	]��Y���vf놓�B:皣[ф��Frɱ��:�8킧�����B�YlB+���9��^��`N��ۨ*2�B��� ��I�᪅C�{uÈT�~��(F��E�P9ߤ��C��N�*��҈^#��#� i�'�@�[x��Û�^�W����l�(�.�a�,3r�05��&�U=o��v�mԋ�%��!��5�s(b����zU�&Ɩ��	���s��b�ݫ��3Gm�S�z�ަ�un�\��J�֎�JZ�ٹ��hy����T|DZ�ԇyE��}��mg�6��{Q��n�B�3k�,N�p�����FB�������Y&z_�*���E�E5�|f.Ԇ�e��Y�YF��4(�0�'�٣��κ���{v2����p�6�
��3m���\�Ȗe�|��Ԕ��E	��r`�<1dV�n'�l�ٳ�X�A\#�z�w����^
x���=�\�b�dx|�����]��S5D/���B���J����u�-9!�����]�۶��s4�c9א{am]��U��|ĉ;�i�1�=~4աZ`q��3�͸�߆���æ�f��̛1�[e���%�������3��g[=C�N1��M�k�
K
����p��bܱ���P�{b�]��3�\6v���r��(��p�2�,�	�X���q��[d�;�]7�(�CX�k�~/���EPn ���"��
�TX�=��<�\0�|}�;oO*i;,�P��m0;u� �6�����ޅ���"��kp�9�m��ϵ�Ʊ�ޒ~yu�f�p�Q{D�>�`�B1���f���(N{;Q*Ϯ���d�'���9��X�UHP��k��*���P�z�4�T�2�hz{����]�h�H��\0�ݽE>�0���� �l"k�^@�p&�pdIio�B���_3E�b)2�����e] ���׍���O��C��L��O�vI����to�+{��l�Z�,�4!�	�f��\�}�;%�q�B6
�X0�����j��0�h�[��-P �/��K�׳2�*p����@G���'�&��eQv�&	x�.2��� ���K0V:T�c�!.i[����Aq&�YRǠ����S�@��Z��������*)��c}�,���d�=>v_�̄��
�	�T?1$L�;�J����I [h�yr[�n��{��0��AD�iq�~`��Lf�0���4�|<��Ĩ?�3�~��뼀�|QA�M��FJ��o�g�H��/ֶ�`�H"鸥�<G �c(�w|�/��OFg��_�� N/�`y�B �+ hY��=Lc4�W�ȉ��_�,�&����|���/4^P���L�$��
H����VOW,bu;��'��}�I['�3�������\�c�p��R�1�E�t�?�$r�G��Ծk�A���7w�Q{̳�!0_^���Zh�u�W�然j��s���訏�h���:�L��9 ���I�D5#�x���q��D'|���EF'�":ג%7s�h�'��&I�����'�X:^^|NlRu���Moþ�~��܏�2��yW�m̛\���R`�O��N�x�a�� ��@�+'c\�6�-�5���7����MA��ҀJ.�Lhnvڡ$�*'�blͥ�����bc�S������P	@��/�om��RX��N�;�P��PJp�Y��vXn�<��W	-d�,�d��	&�՟�8�67'ƌ2��ʻ�m`c���F0z#��#Dg3ܶ�=��a&KK$XU�A�m�9z:�#p��6�:m#��5���s��D�0X3 ���B�mU�r�ki����7ݾ�۸Ӥy$�%d}˭R��'&�rO�3q�we�W.s���zLF�Eֽ6����wV2b�b5K�N~���U@���C�kVCf0^XN�4v�T3�Z��V�J�8���<�F�z�O��jYU��B$��$/Z� I��ʭ�j�,�YAEP�6���yB���=>:��cGtc�0�*vhϧ����$����?dm�O��ͻ�P��O��w�k db��J��<ȥ}v��3n~��n���>[�.F����r�pw�G��B�Ba�֎��#p��N���T��4�NZ}��\����_�ܻ0N�$���f��Ku3ld�_�c��y�[呗��bFB��v&�ňiZ����_�tQh����B[�N��������f�6ӰjΙn��$2�f���Gaj����4v��oy6�(�o�$H��%Vۨk���B'����*P,�'����=#�qy�q6@9Ƿ�Z�Y� O�X���'��ΝW��\"��nC���",�f��E�W_��N�y��|˥Fg�pM��[��7����U7TR���Q����  ��*�����׻�
A�NI��Đ-�TC�����R��_���$apl>����;ox	��h�{X�'�Y���q���X��Գh��D�U��Tg�@`'�� �f�B�ߟߪ��zb4P'���# w�g��$���h(�N�I�[��걼))w���\�A��
�?�i3�@��ٜ�jG^r�X�:��Jw�o�1t��1F��h5mK}�4�Q�^��=F��~�c>>s��bNi��`���B���]�^�M��F�YӀ5��הp��vS�h�.��M�u)����-�g9�%auJ��O���������W8:�iZ�3�kA���k^�\����‪�*�Jw@V������ŘN�r�)���w�f�fGSI����!m;����ѷ��ID�n�2K�Gx0�ͮ��]m����.�oю嶀����J�x�Y�=�&�[��=F�R+�`[5�!F"?�ޜ�=r0�uG��y����1���=�nt͉;����f����e�
���?���,50K��Kw�!zF2�Z�I�]���z�$�G﬽���.*��j�.�o��-ec�M8���rOVV��W�.j���j���J������_������MGY\�RP�6��:�s��8<alO�q�NJ�I��7h�kte���Gv����͂.�)�V�`+";/q���ʲ%5_�@b@%H�F��3�m�f��^]
ʹo}(=Io��
'�ǿ��~%�oK��E���bkB��FM}�2'�w��>~����A�G���#��	���6_��Q���h���7�#�IX.@��d���l�Hʫ�4��(�{D���D��Zm�Y\]�N����׳[+���8��ۥb7��*x8�ܮ� ��\J��PZ*~�56��x MTg@����kA���K-��c1� �Ȩv�p���z���G�\@YqM�A<� z�7gg�/��|�"Tf��Sx6_��OJ�Т�T/V�ckA7a�_	iϯ��4IXM��G�[�@�&��;韛	賍���v����a_ʲ_X� ��O-�b�p�<Ш�������]0wJdy�s���sX�>QE Q�0h����~�TױH*s�ň�n&��1���@Q7�mG�aٹ#���)0�ߛ�6��'�	7�-�1k��/������-r���&^Kt-�N�%M[r�p��`ή�ᄗ 7��Cj,�M�\{g�5���h������͗V[����7�L���گ���`��Z�q��To�
{"W�����ɴ
�����9L]��C�T�tyy�Ki!�n��]K���j؉�>H[���X˔��s�S����w�&��N%o	�f�3���s���K���B�������t}���5��s���N��J�Y�Nx���ƻ�>��H���nJ/,�aغR�kn&?_ҷ��}J���C��Zs+%x`�{<��G�Z�Q�q?�DH̚�R�K�v���¦��}Q�Yw�׈0&�-k��{���EC����D�J��q'�T�#��MH��w�Mf���3�L�C.d���^�4sH�i�t���e��̈v��?��A��[��4���w���1�PX�Җ��U�hF�cO�TQ:̫���j6���a��/�4	�yE��rP'�6*e'�_�#�f�J�O�R�^<�0j������8���S������8�+�G�����rM�jH�)�؀N.�P��V��`��M�C��S<�*=��ǡ�?����I�h��BY�`�[�ީ����r��p[��Y��Xy��NX|��jɠ�٠�ɗ�I	-w���J�G���U�LΗ&iŘ9o���&aU�@;���ބ�A@o�*��l��TA��.{��n:-p�Ǫ1�R��x�æ���:3�~]��_�"��7�}��\~7�|��"{�H�,�,Y�4Ì	�-d]�5�U�fU�(��G#Vђ�Z�8k��/W�O�Ws��CP*u˴��O�����a�{�9���A!� ��f.n:�@�u4"�n ��j8�D���Ї&��7N/K���\aN_]v=a���+M'���Hb�5��	֎��� ���nf\U��My�#�h�_ay��>,��dFfz_����A�e���LK�HI����I�EP��J�j��Sx9�Egy�,����V� �o���-�_�*+�Rc�Ȼ�9=�UM�	ݥ��t'3@�KL}�}����B��*嘶�����A�p��Կ�F�$��a�I�-yv���Sj�/vl\�
� �C�O��M�UI������ȵt���핺SK# �6L�Z�<&�٧�£��?�Zd�9w�N�i��Ԝ	��v��]?���uï��V9.8��PI�?�b��ˋ��~8Fp���3�c\M���^���w�UZ��D�	p�I��c�}�s�&�<~|���7�&jLnQ,�c�� X��9=�ecl��.Ҳ��瘶���e�z|�y�?�9�q�*���x�.�oe�A���=�7	����އ�tzj[*�W��^m��]�]�|}�z)���Oo���@N�[�W����ky|�7�.deS��#�J���7zQ�S
'EM�e�|�\~�3Pߕ�Ԣ��H$�X����r����1{�IDti���>U��!�ϰ	A �%�t�~/��W�x�ą69t�_���u�\N5[�abHf�6lUW�J�a]�I�y07Ђ֣eF�=����8�J�Z �B ��W�$����+�� F�%㾈/���p�ޅ�)7��"&��h)_�<+�-m8gq�HƘ������
�8�(��y`_�����i�9]TL�PkJ�M�0F�����J���.�?��-{#��f��:P=���O�r���)�)�����R�fHh�_MHG���h[��Rev0X�'&?�e`%0e_�3AT\���5�З��z?�r�r�vg�h�^�Ц�s(�Q�>�rA����a���^�mt6"W9��T�LҤ�Cm$�k06؂P}���,�/9|	���E;
���w���s���_ Q�V��h�|���G��_\��L��s���o��Եgs� �n�1��Թ��,���|�@/g+�I�vA�L��.x�����!�'�h-}��栞��?2]�[��7�KS��l���e�y6}*12��^��ɇ�t7^�-���J<H�?R/Ŷ]#�-e�G���~��tS0kR$ug�i������xw���*`�>�WSiܬ�ԖYTYA.�	�w�����S�Eؼo�;i!x!m����o�]�K�hd'U�T����t�����)jg�a�p������8ESkw.�,�;��]���.q㿛x���~��M���ߪ�b�ʙ�&^��O%�3�V!y���B?l��.������	�y�u%E��䤎�T@��N�ѹ�U��i9�_I7���_��d|t�;�7����
�kx���)S	l)���bJ �����D�(��qqW�9*�d;���E���Vw�$zt�ED}��o��='x�W3Q�7-f<8##m����P�+�+4!t�����*��+"�)D�(���b�hd���x3��A�4wW:����$Y ]ĶӼۇ������s����-�d�w�t���0C�̀�_8�z��}[�r�T)���ew(kn�8BQ2ۥ��b�2F�gB�T�X�M!^�X
��(�?+�<0��2��uH��X.lSڦa)eo�+F��lJ�Z�r%Y@:��Y�$P��扫?qvk�(������	��t�Gn��0���w���7q���Q����=8�15K�!��F�uk�c`E�^�B|����iXy-�_AZ\ zb�E���H)(bb����(���?������u{~��떠��4�Z	Y+�D�N�\:�ɱY���M5�fv瓕`�K�\��6K!2c�BO��lFdE��?b��p0y�q���6�c�}T�rެ����x��K0��޶�^�U=v*3<5�0��(�=�* k��ӟ�u@{Z��Ya�%8�Z"~y{��'��k|R}1@����t��G���#��+�ղ)�����*`�gxFq?C��g�7i��b%8�+f9QxmP�(�t�-Δ?d؆�_\ ����:�Zf�7l�km��E�}�P�\�8!Ԡ�E��&,�R�\L�N8�()���4�o|E�N�E�"�mgɋpLo_��0�=\/�*�� �~!�^!�?�q�~�K�4>�&w��d {�x�I%W���GFUԐ����S�/�4�<;�𾕍IF�G"��Y��L\�����-q�'���o{�x`��=خ�'���ؙ�Z0�V�c)ɜl��PH��k�u�O���`.�l�������+�x������+��7�;�M$�4z�1=�}p�'�J|\T4�.P�f��BJ!pKo���=-�^���sb@���[s�9�ާDW5�C=>�#'Tȝ���8|��JR�X�v�=b&o�uE5�G3h�J�:p�b@<�RY-��D��\���-�CY�����/���j$z�������	s �5i$�\7�s,蚟E��.c�����\��>�y³��o�n���؊�'[Hˍn�2��Y�)������K�ӎړ�\fG�9����,s����-v�9�J芫�f<�5
�3;��t���o�����oa�?�5gV`!Jn;wO��D�|L��yY�hs6��c���=o��Ϩ+蓗K��=��u���S9��d�����X�N7��ް��Vx+�A/ף١�ЁB8{��E��6Uk�ռr2���ݓ>���5囨��>��B�~����E�z���	��=���j�7�B��F��lZ"�Ʒ�\B�e�����r�ƣ[P++
i�r��h�/��7�˴{f}n�x.��*��,${�h�z�����-��$D����y�P�H��S�-8l����4�	dt.$��y��s����H�먓�?h�C�7�6�ʨ�۴����7�ǿ�Ƣ��8_(��g�=첬_����M���=���w}X�@�O+�+8�Ӳ��Q0�^ ;����>_*��:���N�l�I4�޵ �h@��G�׈"��W���ؖ-�d�û���ʪ��lyP���{����������?���8�w%b��'o��wU��T�-k��-)����W�&A��Ǖg=y-�CJk|���]�!�,*�aB�I�`�&ӝ�LDkh��\�(d�"�FXB h�8�>5r�lj�����t%�RT����v���t���ߌ�ǯ�u
�MJ��s͇J{��"���P�fI-�@އ���
�+�Rhf�1�b��9��bf!1K� �5T���=��C"fp�sv�N\=��=?`�ή��kF�'��S��uF|���C�G�A���?���QCy҈��'�teB�'���U���թ+:��4tƌ�Z���D�(��t���M1o�����~3@��&F�S�4!|?�I�tΓ,1��U���C���9�0�l�q��{N��%y�>sx
�F�sZ !���\3`"�Q��A�
YƎO�8�2������_~4Q�?/&�����Z5͊��8kp b��Y(cr��7AJ=wJֵSaa�jPH�^�It��U1��[z���O
<B�#`��ǂ�lG�2]�FZ�KG��9�%qa�=ܒKy ~��ᱤrP����1@o��{o��km�����3�u-�۷
�Q���P�!n�M�2�p�'��p���ȌQD��Z�j>؄�H6$��K���O���چ0F�8ΎC�6u8���j�mi��o}\@ҍ*���q��WJ�k=��"�Z-d.���>k1�F�,���6�?�"��NnC��Q'�
���<�o��6���p�#u	�:^+�`[��Vw�zBvK�೻Pd�8��~��:L��tU������IG�/�T�!ښ�͞�3�ʔ��?H7�H���L����݃�q�sn����ɬ�CAF��M�|���_���Y��Q��y�2	�k���V���s�)��\ Cz�&�=	&��[Z��¸.���E��'4W��.��W��b�}m��A����3�^^���#���lX�/�ǆ����'(h1}���ϙ)*���<e�{�=;�"H��UA��qU��EK������G.k��Ya�`n�%FuO|�/����?.�z{�C`�3hMw�T?Ǚ��P|l���n7�g|�V��m9��.���9_Þ{��ȩGUf�HԸo��9��h��2A����`$9�^��������jcq�N��U���}Ӭ�6���پ���u^�I�]�er��CǑq���;.F�V�O2��"�}F֜6����2�R;mG�Ԥ���S�^��خ����H0����h���ͣ$�S��@Ok�'6��"���S��B��H�vm'��7|�Xd���E��婍}Y�V�,-��U���J|�V�)2�,2���	]�+Ji�����m��j}��kp|��zt��;��??�{a��@>:o��IE����y3��~^����{�C}���G ����L��B���gdeH$�;TLBh��j0��`qh'�ȏ:�Zт7�����b8c�c��|��>%�b`L�ײ6�W�����Z�o��f[4p�d����>[�K�P}�xl���M����|kx�t+�ʷ�1i��/uʽ��m�-i��ؖk���9�c�A!��1�1���#~YvM�hw���x6�s5��ޖ�jbJЪ#�'�Ji�W���ci�FI�������P�Du{҆���r?�#i�^n"�q�Dr�z!,�'ķ���'��$g����k�g>�}`�QI?Ȗ�R�!t��ۢ��]6��pO�opR_��F$E!��O۟e��������1�Ѡ�(]�Ť���E�^X���j{/���&T����Փ���~E�@Iw�ߡ�ޫ��=�����?)x@��m��6����~8QFYj:Z�P�PUn(���p�Z4ȯ<�^k������΀%=�I���[�ݍ��<�����n:+Ui��cm�k_��|�T�¸+�,5�ck�sI��1�ĉU٦2�␳��E!H񠊬�V�%�%9/릱K͠���ж�)`$���qy\�xlW�����,��afnk���ْD��|W����T44U��/#��jD�dg����ך�8�w�|װ�qD߁ӿ�yOT��d���_B�k��������D�d�W�XK���_S��(��0wd����l@a6�A���xd�)�e�� r]u��q\�nq�QRh�"��t��Q1�ϙ�2�t^4�K�;���G���(��4D���u6�|�җz)!(.�7�NM�1Ys?i2 	)24��yᴐ(��)u�]�h����f��e�ʒk�\Q��&�Q@`���o��k�k?*t]�0�iV�o��AV.GB���ҡ�W�CT�<��D�W�Wro�Rr��;��$=����?�ZR#{��,;�:��be�R�D�\ږ��Ѱ�5Ӏ��r,�j�z�
2���~�X1`2����RZk��Dc}�����
hkH���#H[�o�a���t�h��~�x��I�|�=a �<<���
V�s��V���]ؚ�:4IN��y
��` "����4j��#戱0/w+��6��~�)QxU/U������$O�'��H�V�]up�k��2���BK�B��Xq{nr�w�l�Y��!�Fh/�s"h*c0_�-#+�w"�}\�](���M���b�~=��	���<SԒ�t����x��ZF��_�V�\��e�l�J�ūzض"c�������d)� `V�p4U�1�s��v���� �[\wUB�mnV���v����<`�b8�E�U?U�Vȋ �������Ԁt���
֘Z�H�RsL+Ư�'�qFU�����d�d� ��ߐ��bS�.~������:~�v<2*�XOz��Sa��!rX�.�
��lc�@� !��d��+tErT$i5���=7�~�}�'YO��E�ߥT��RD��yiq��DS�}�δ��7���}��<��`�&��_���N@�U1���:�)�� z�?�������~��C\}{lf�~oՐ��B[����01�Æ�8;�Ϭ�f������.�&)��Ǻ���Hni.R�(%��q��z�aJ�f��;��-BMv�I@����b���b}ܬ;i������oo�8Φ��J7P:o��p^���Y�
�V�BR�����p��n�I��t�0\�b�����V>��Hv��2��%�nb�s2�߿E�ʽ.QK�j����0O⽤������Nx{�������a3����aȗ���8H���_{�ty���9���P^��y�z��,��U�ZIYe�2t:���v��c߇��p"z��l$+ L_�3Ƿ��|R����AJ	�ϙ%�-���+o�b�T��)�c0;�Bu!T/�pL(���)��gk\!o����/����d��Fw��4AT'�Ud�Sb�`;��!�k]�=!0�Ȟ����N
�^�����vA���9:��� ����{ �]�U,���^!�%�%III��#R��}�#.��)Y)<�������TQ4�"�����eFNt\:\���E=;M�6��d� KP�=����ᒨޅk�?�ת�A�[`ۇ ��9Q)f����y#�$sN�w�Q���:�f5σ���C��p9��˼^�M8�O���p�a�m&���`ש]k>׆οZ����9X����VG[,�ڙ�_m(F��{2R7�n��������d�Q)7��{lWQZ���}KYcQ�]x_'�E���
�j��!�g,D�����2���|�+<������˫	Y�@*J�'_	�v�G�n�w�TUDAB�G��n�^cⲸ��~9��:������ͤɧr�+!}�#��
9iIӜ%H��6M�>�`Th�g�W�sݏ���t�0A|�������&6W�"���b��VL��}^S8f���d�u�r�-?�������*iM�9]u�c�ݷ�w�H�ɋ���c�ʂ�x�&��aR?�$�Ԉ��:|~Ɩf
� ���V����ߤ�[w(�7`@Ow��U26_Wbʀ8�+�-���O e�	�J�@�h��3���{=�?KM� ��Ͱ�4lc�@ˡ�F�&,@QN/]ƛȂ�b�U�����`y�Y�פ��.��:%��u�Q�;ec@jv:v�,�>�B�H�b�l9�->,�9�y�f��w��۳��JS�R�r�΢k^Q�8��0�y�8�Ic��T�2�q�����J��@����C�`iR?�QѠ�w��ῶe*Q�L��ӎd?
t�Lꚺ<ةݘ�t@ߓ���H�en�qu�ߡ�'*��f/�C�P$�������a"ݵ��cȱ�]
��U-�kes�0%��4aLL�t��r�E�o�zG�3�1�����gc�'����)���
W`NHPl h�4��±d.P�cgR�@F2��'xC7����3C|�P����Z�[~E��LF�	H�(=�\W�U�x����]/�P��r��%e�2MzPSt�����1ۛ���GߍX�)b�ņ4���\������<��ۓ���f��p�"���p"��z��Y0���\�|���e9�&&�ֈT��U�� ��3�v��!A�O�r�p|�jǟ�݅
l��#=�ե0C�u��+]P��)$�x��K	6���� f��g�����'����4��WX�"�g��q�:�t3b�� @w��<���Uk�����D�V��F4X��Xx:j�J�z��m���.�ol[��2ɻ��+ĉ�P��7��hm�k�_QJ!�S9Oс"�3L����7�[�j*��p��Ė1��U�n͍��!h�3H�������^��O��m�ς�F
�O4{(�#�1��C��C��}e�`[~;!�:�G�O������D=fbв��A]k�$��)�[
@{9z�b	�6���Q�3ťZ&Gp�W1`�ؚ���V�zø�;^1��2 6��~�I��ؗ�C2(��;��Ū���K���b]I�Ά-���R=㓭B(G�N�S���z�\�0����%���$o�k�� �ϴo��!�6 ���:Z#n�!��daZ�?F�HR�}�3'ȓ��4.(G7�r\}(- ��,� R�����D�>����b�1E,V+*�_*.o!��:ڼ��C��(�d���8	���9��X�Veι���1G���NF����2 ��	��KW��z��9\-�g�"*�5�7��l�H�5j���
"�BB�d�`R=���(�g0���0Н��o��.X4����>�\K�&C���n
FmzQQT]=v �Q/�1��4k��������(&`v��q�:T��0qtV��Ѡ`?@9!�3�ˁ��}|s���r3�P�������)-���v�]A��[�������YMQ>���S�P�ǰ@��/�т�㐼�e�4�r��.��U�58�X;����d_�j��)�qF]*c�WO��l�� |�4zs#��
p�D$��1�	�4�B�hA����O^f/��#��:-O��JO��BaEa���8M��xÃdf��0�([j
|���Q6X/��A�y�=��1OǢ<%e&���vI�rR<���Jw�����(1^��3

����7ߎNcSp�U��ȷ��-��dN��~b��R����Y~>��0,�B�[��0�Z庳 &	�+&b0�zS����G��oL/S��xf��V�Ƙ�6w�YR�}F��^n�]�y.������]�f��4/��$�߃��#K"�C����~��OF��N~�ZQ�:�S�:���>':�uG���v�:�4@=[��Bv����V��g���a��Cb�Q�'{�%�ki�<qg��$�F]c�a�a�k2i�ٔ* Q��A%��`x��ƫ6؂V����m��`Dxz�B-Ηkc^5~�/F��煺�t���'�0v}���\��ϭ���J)mb���#���6�L�6��E�מ?�/!�(�񙙮v�w��2��Z���Ҭ��c�R�M�^���ER=`���	�]���Y���i��|*���TR�~�E�lM���ߎbJ�1��M��h��E�q�cآP�������Ǭn���$]�0԰��N+:es���1�vN�����R�|c=D���L{����qw���at����Kp�Hr����έA�L�뮔�s`�Q��������O��ٮ}��!�	�#g#��=��ؐ���х��P�.��-VP	����%
���x��,W�C�ކ��l)bB�F�C?��"�������ck��v���%d�E��t��R~�EZ��m�g�_M�[���`'���T0�L�5Q0���˴J��*��ruUx��>˂�G���}�2��b�QB\D����I��;el.�K�f,	*�P3�XD�;�n��.@׎�<o��AՑ�"߼�}�+Y���oz`s��O���h*��)�OTO(�)�J��$�o��:�~��3b��$�	fj��VdU�$�s@C��ki8T%��J��9�Ɇس�&nZ�$`���S-ƙ�pw�<�!J�ʳoǘw9��KN�+�Olig*����G�.v��rޛR����q��s�M7{��yB(Avz�ɸS b�h�fZe.L�>yh�ysdm<r��.��7��v�;�U8k:���U��^Yf�t0��Y '?����T#>N��ޒY�H6; <q"z_\P���E�q|���E��\$��?�x�����H�a���� <�	h�%ZѸ�m�L�D����@m@>���.�|������N�=����ޣR�[���q���`�*��i�l�@�]��%]�����;�)g��8k e	�D<>���"��H��D�7^�-�Z+�F0j�9�[UZ���(KA�
O/��$�h�GG�����n�B�T�he`�;�?�!]��^�nk'���z]�C<����F�����f��-�)���ː3�>e�ޮJ��+o`5�G9l$�5�L�3�*ĭ0h�> ��7�O��T�L|��P��v�ʚ�y͋��A�	
	�!D>6�a�o�s�s�{s�R���g���'q|����9�Vi(��q���۾��ųe�%zS����ϳ���a��J�k%Ͽlb�xIIi���zqћ��J`�}�ZW��+!�똣�L8�R9�D�Q6H�Ԓ��D��<`�����Hte�;�P2@#~B�iؙ�f�}�|L)�_��{<+��H��:�+j39��q��͡�E�o^������`5ž��.�QZ)t�o���	�����>U�9���t����*�¢C�e��(A��� J\���p��s��)���[�W���Yi��_:�"���:V.�R��0�m~���z�&�mf�/)�7ƃ��O%����\,�vqXx�>P�.����u�E�Ր!v�1��f!^��� O����f���ڼ!:ʏ��������C�/ݧ�ٹ�d$�l�;r�29`6\kmc��!��<	!�Q�a�����b;���Y�9^#���@�Q��϶��P���r�)�6[���6�	����i�������:��nAq����[$���i%�,5�DS��<�to��-T�����uL��2�ĞI�rD�p�!U��`�;�tׁ��)�Kp�/!���gΫe��My���7$����
������Ւ�@�(5���H���N��Y�=�\���."�Q*7��S��$�^B��W���L ���%�b��)�#Zݛ���MѸnq�8��2��(��E'��u�2��޺J�l��IC6���H`"R�6�Oi��ރ�
S>B�'�]:�-��c�@�Y����?��+�.{�i��֝LK��7%�O�\J�����E?����<O5�����Ç��C&&��o�
�d�our�F}Wӿ��Q_	j^�sJ"�`�YG�b)Q�XV��}@>�$}4� �M�g���C��8X�?��*�%�'�9B�pp��g	��Bg4�.㹿as� ��擃q�J&G�O�vW��|�K�38.&Ua�	->L*�dQ���}N�%����Ҁ�nj�������� h������z�� i�	H�nj�g��ӭn."��8���q����N��I����	ED�X���W��h	�iO�	��e��PLNGg��	G��W�\(Ȫ���-��S��]��#���B䔖�olQ]<�k>u���L�3U4�ID�MM��ܽ��hH��N+x�%�-J�w���C)69u�h_�TVOM�CF�w.�~ҐY��ۙ���;P92h��5�w���M(�E���Co�19Bn�
�h���v���xC��W��y��L�ꁲ�-H��"f�]�m���UlQ�iz)1,�"o�,�l'���(f�zj(�e�iKW�^��"U6=ť\^���r0���g�!h������C1n��c�`3(�n����3��S�k��J���=��=�&�y<�x��wl*�����l~E��BVr
�FY�/,y�����.|{��[�����)�V��0I|���VP�s��M
���ODRU�*�=�?�4U�c4�Ov�| i�m�������\�ג��AʇLj߳��\sJPF+ ���_ʹ����?8�9�El����}%?&[E}�����n=BH#g��5F�o�`6#����V~3S�z��}�y�.BKZ{��XL�l�$+_ ��Z��Bh0�ć% �����>��K�a�u�w��/�G�'��i>�)E���/��������zK_�w�*�3�A��s���\M���pֵ��_�n��(�ǀs��D���-,�Ȧ(L*ü(̫�W���Y���0�V��a��v���ċ� ��e�y2[)�V<�1b�W���p�*�i:� �����M����O�����`Z��!MH��RW_�oO���N\=�4�/�8���٭%r��m���4�H����dvg
Ӏy5��b�.g���ߡi>I6�A��*��2VL,�v<��PS����4\��z!/G�!��g����TӉd&s�x8�−ߎ��Σ$�k�?�� I���6�T����D ���R����)��v}&$H+mq�t�A��Uaɦ�v9GJ���.�{1[%Ʈ@�1 py���i��_2Ot�=�Lh��t�n�YqӮ�����j�CdɿGw���U�s*�@��8�Ң���C� �+�YS4�Q��W�J���mP�\A��O,RL�I��g%��H�0��u-�L������U,%1u[V������R�lπWj�Gj�,�Dkr�w�0�3�@{6B�~��w��O/,R{J���:�&��	��0_ۋZ����)K�PL���ل��r�+�/�-0�	u(��%��P�
a����nZ�=������]��%f�-�����u�3?S\/��^�`��K3����KS���{��5�"�c��~�k�wc���|�2�PB�1��9n󺨖�?7�f2]���w���֋�B�(��T���{�L��xt4W��P�qL�@2����4��ߎZ�h�	�m����>:l���������?k�_ϕ�M�a2��t.��"��Â�e8�ʏ�����ll�s�q�����ƭ�AQzo��R�;aK�c�tn�M��D��nZ�f��!�d�b��.���ᒢm~a4��x;�dzeMzk�y������(TE�d#Ӊ��F�Z��ל�,��N`�1#8�rKPvE�7B7�e�y�?�C��Uz�F�w6��&�;��M0�:o�HDh�	�I�Z��Y{?��� e.�9�%hJ���Q�1�Yȳ�w�_�`�f��6�4;[�1ڷ���S^��K�8r�%1�a%���-��(��v� ����U"�s�=�3CsP�j=������,(��k	5dtR�[5��u���S(|�j�-m襲�ˬ��\�x��mT��F�9P�y�$��dx;�8!�>D	Vd�MF���ا�h�����|���,m@�Ez���0Y�²./r��Gl
V�mt�۩�����l�K�P^��]�Y���¿&BW/��9���Rq�vZG���{��i�a��_<���|��T���W}x��ڛ��-�1�t<5&l�!�AB�o2^���I�7	�������Lp���m��"���1�3뱪܆N��$���R�dƯ�^N�V���0q�� !n������]�"=R���8�c?n���Gifya�Ht���̷��[J�*����R.]	��g:��P���?����2�$�pX�0���O�h��Ch2�>�X��@F�+�Ī�ћr��H6<|}��"��K���6�Q:�Pk�����I:��v��C��:�D6����a7'�m�7O���[M!����� ���k�d5��U:��4j���բ�U6"�I�=~��6��%U��%/B�������29��[z{e���ؗ�W�H	�p���sΗ�0��4N�7����n���8� ����U��+�l��&K�?#���q�.,��1��z�S���J�~�G���t���.ɾ֚c9�	�6�o���Qݬ>ק|B�뼮e
В�G�r(���� �̡s��(S#�&�h�=K'�睩�B��ݥ�>]�;�x)�m�[p�����
ժ`Ɨ���<=�҆4;!�� ����kTKЇ%w��Rr�����ɂ��)�Kn"�**��.��d�'�9������5E?�,����4N��AT6�U�~�RO�vq�j�,��N�4��9�v�E*����k�_be�\�Gڳ�/�����<�H�:��!&zV�.P�9+n��{�b!�k9��{:��ѝgi����(���<t{d!{�ɪ�ot�8vD�ū�-��U@䎔M�*�ffʓHf��_���_�C��O����P�=�u�V�NO=x�YB+Յ�u�95�ko�ЌqM%�U/y�Չ�N!�hejQy���n�S�R'	��j�6r\���OU��:�;���#��Eā<3�_��۶����k����>���(;/�@�����KI�-a�z�8viyE#a�$o5��}�M���\N��x.XR�a�/�3��t�bhV<���?�zAv m�;Rt!����b���p����[Gm%�!�����r{4�?�9X��D2��oH-�b}{�Y�5�n�`8�HAq�g���k��9f�|�B*��xVn.���7�+��F
�:�����~2���(�hU��݈=0�}���1�0��7��޹���L�9)��~�?�E�p���t7�9���I0���ὣx����h����b�=�ȹ�L��ݫ�����~�?��p����y���=Y�+��<�qc۫[<~�i���B���U�����f�5m�G�+��1���k>��Z%J���B�'���o�b������C�&L?�g������9��.Z���[q� -��q�'���������DKY�'Y�*PV��Ð�AY���=i�Di�r��p_�@�Sx!�9����!�7�z>��=����I�$��!��t�~Wxh�k��!̭�t������@��RnW>���[Y�tdO�s\Z���St��נ����*��z�z7&Z�{X�H�H-{Du�"pDP	�`:+��tb�G�b<������zo�{�r�'e�[�N��������� E�l�X�`� pL����۩SkM
�t뀩XH��Ny���[��н K�Ʒ���trv��f`�;Q�JO^�_��o	�;6������F��Ai���`,లJoخl��P��`[+�B�U���v���#]��zx��3��kb��N��U惪j��d3`3�E��<,e�

E��8�bZg)� .ہ>�}V�x/B�5�x����d�ڽ���/������^��r��s�K^��oE7��>p�'�ß��$�'��Y���g��N�6ބ�B{���أ,�5nڤ�.]>�zf"�e��K@���w�n�J1��/6H;�٩�8E�}y�A_���.L��*��G�3�=Q�:���nU����e��Օٴ��V�3�S8n���l�P�����smz���Q�B��lym�;ꛢ��u� ��=��F�H͚{*d�/���o��0�D�ʸ�;ɴ�o� �z�|���2�`�7��O]k�QT����o<�B0�x��j��=�~�>���튾?��j��>�C���/(l�Čo�JCԡ����e��Dl3(���<��Ԡ�<2$o)G�?�^�[�(u�-��c�y�￸l�X� A�����G�ۺ��q����A���9u@���05��bs�֨�=����y�@��'�-���Iìp5ZZ�U6B�d����;��ZjN ;��v�ͻ}qa���B1�J��Y:���7����B��I���?�Fu
59A�̕[�.&��M�w�����4䐘	��Br|PW�Tl廙YH��)�q�y��n!<�]%��Z�l���vX��\>G�x �Y���74l�7=+e(��y�ث�i�c瑨PN١;�#�l!�Bj�����Nk�\���b�A�r],��ٙ$ZЈ����J����^��9�
�q2��J���/kj���v��!as����Q��.A�X���0�Li�P �K�~9��Sb�y�6͊s�`g�Z/��l�A���􍐟��:�{r�x�,��hy�4�����1�K��7L����}��K �
�Yj��#b
X�~����Q�S��a�n�&��˚EV���Պ�n��+�.&�ő�}yk��[�I�����`]���K��%�`�������D�QI�,=��߼g[OE�S�K$^C��[����g�RM����Iw�f���py�hj@Eo

B��(�X`y;2<X4"�r��f3��I��~ۼ�q�u��m��mTd:���`B�&�����]��|�m5��6:�"�49}Th4�GG'�̫�p�$��v��KB�0�=f�c�+:�{l��Z�F.T�谉b*�+�72�S�[1�l�>MV����Ѕ�J��{�mߑ��}?B�e8e���A���jCR�z�%�!�w�J��̗.Y��A�D���|�nR�k���F���A0����h�L�?�H��-��S�c��ȗe3�,�N�ˌ�w3��梐p/�^_���k�U��v����`5�q9��U$��1��:i�<��0��	k[{�pӷ�h���т5�\\d��^g����~��3.D�א]˿t����(@L��:�ƚ�ـ�L�i�	GR7ǈ�3�Ф�i���>i��_����"��J�^[�e��i���l��_���1�s�aGJ��E'f�{�d`L���C{p�}�� �^�'g%n�,�\S��T����>��K�~��*W/� ���i��
=ܣ�,̞�z��Q�[�����ֆ������L���G:��Ą�1��;��=D�I����F���5dD]j��p�]�9�b������D�����_��ivr���r���M��-����є��J�6� �+�{�{���)��i���7����z��
Ъ�8�Z2�F<�RRY.8�J� �^'"�ǭH=
�wDc@.f^e����`M�e�<0R�����b����-��vV����]�r��B�ôΞ=@+��-nw<]��z��>�s(0\�����i��~�>�L����U����Byi����I�B��a�B��^5��2��,i9��׀g��.�����q��N8�·y�9Ԇ��`n��˟JuÐ�
�WH">:�u�4���"��7������x)_�8�J�7�1�+�+��~�8 q�����Q"x͑1�b����
�3���հ���h������'�=��Ź�}���H���`1檐��JāI:��S<M�}7��S��zɼ�bZ�aZ���b���?��&�0n��\԰����n/��>�s*7��nÜs�U��&��f��;E!���co����`�b�1z��K�fLH�A]������}d�f��a�������� ��,E��#�t@�wT�-zY%]���s��8�ס�Ȫ���][h�e�F�m�ވ!�I�Cs��������>B�M ��P�mD�X��~yJ#
��Ǒ	E�����^�L�)��Ub3�,̓Rӣ�ed��B/��VG��Ĺ���Z!*�Ο���a�'����t�.��1m
9EY�t���1f��qQ�N���].�����lԈJ�/Tψ�5���w����\��LP�׊gq�#�"����]�	�IO�%�d-�R�%Kah#<Q�H��E�6h\��N�{�+�E���������������������L$π8�',��2�[)�{(���R֙Jc�f��&!���T�\C�a����[���!Qu��]=����\}0����a�ei�rV���`�a!�ȵn��$���[&��7\3�(��BqaZ���)Jr�t���E��~#�g���T���kaD֍�I���sD�K	�Z�b�@���&4��� ��FsK��D�`W	������r�>��|l4��>f Xa'.����M�Z�9qƟ��K�FX�P����F�]���$����u�2�˱�5nmC$D�ԟ�E���28�������y����v����薧P(�j�H!2�+�i�	e�m;g*�٫^'�P���d�`��y"_u���u�" �ӣ+_���2n�	��P�"Ӝ�o�&e�p�-��i�ފ�NX���Sݰ!���4��c����S'-��&�E�}H�u�����}�L醇Obo&ݦR,PѮC�g5Q�	�EX,��~����Aw����\�t��y�&������Vb���$�b�IM�&�Ou\��h8�-:3~��a��s���0����׮�����}]Y�ZfU�m��,�L�=�K*k[�}՚S�d����׵���!`�>��\��3BXW��� %���t���vtdѶ��=��Ѵ.$�b����5P��(��#F��F,d����u>�}��n%�=:x9b���v)c#�7��H�Յ&�U��щ�^�v�>b��_�9��P!��i����dbUj���3�j�ɀg�\��kp�Lc��������m�?>�����o����?{ێM�W��՗5L:�z����/4!����� \\>���;�l?B�I;�yٱ�ޔ��I�a��������mn�#���s�L@�\�IK�8ZV�������%`5oYN;��r���,YX@����AD�RӯB+��?�S?g���l7�7�ڈ�SWYl*7��af�/�N���)��;"M��x6h���Y��vj)�A�Aڥ408����qk�B�-���%�βsj�w����k�'M R��ί#i��K(���+�2E�߼�j(}��G�v_5	>�/zAk�� �לBs~`�Ό�j�A�I����Ŗ���wQ��E@�@��S3��H�H`Y��tJ��y�0�t�eԠ�q�.� 2\�.���-���a�vi��������6�P�$o��+���U ڃ�j ���/���/�i�<�JJ�����{��I��C�m�/�+�mP���i����I�i��1(�c7�?��#�38W�+Npf�Rh;�"u�zK�_�"2M1U�l2�N�Z��H�ΏRc�`8{��aи'p;c+��p�
Y;h�B��=�����$���Ґm.����AW������O�%�=����;��+C�	������b��x���V��X;Pl���Ŧ5�nA����;��}CS�d�3v�}I�Ju�D.�A`MY܅�S��H�}5Q_3��X&�� %��6>�L��]�+����qOs4J�DFP��$���Cܡ�f��M��&�콼�K�_0�����|�E'+fХ�"�[�9`��m�SuŜ��o��XH�Gqq��G{�k�aD���K�e9�h��ٰi����uZ�UT��HN��M�\��yg[r��V��b��dA���aT3���wƌ�f�P��2��$��j���N��;���iON(�Z��k��@�ēVRb+�P@�gJH+q�]��׉��
kG�t���OЂ��:��W��)�*���J��'k��QR֔�]���7�w���]��S�1�υ�ꕍ�X�7��ݪ���P��^�_��0��[_3�⢿>�`R;^�)��wr�^�u�::���������|���	=��؃+�$�J�;eo9I0�5���Dnԧ(�q�����3����\�F�~�\��ꪎ��M��lԙ�h�l�D��U۞�-�� 7�� ��{�2���P2��]�� CɱmS��b��@�����Mr����V�G�N0�#�_/��q�4��_�Zyx�>�,�:а:a5��$�@N'�*����P�� ���<�6.��L�*NC�z75�����]�'WR4��m3���"��$��c�,T���O��$ր�1%)'�����}R�tYM�[�1���:(G֮kpCD�v\�X/uu��7��`lp��rf�(�:�6����b�|��@�0�s'�a~���x ��K1A�_�\��~�H ��x��/e�~kU�u�R{���t��i����9۪��w��J�����y�H�w�I[�h�˥]�8�$ ��=cv�*l۴=�7oea�7�(�d�Z$�~�Y��v�,幍ˮ���;/��yɒm�'�����y.�
�yp��r�O�鿙���O}��׀��xBv��QaϵG��{�ޝ��?R�	����$WӘ����	�B-És��\��Y�M��̡�Q�}���佉I|W���%�Ѵ��삒����y��k�sN��a�Ķdf	k�����oy���!�m��~R=�iۅ�W%J�𕍓�`�9���S~0�:,WX ���4������3NB���957������׀�Cˌ@��y<q�-�G��T����c8 "힢z�,���|.ϧ���� C�,m"WJ�S����o p���2�ë��]�s���Uw�,�G���79��Y{��E�W�A߄1�����s���^E��'���ЙGt_���$�� w�ᆫ#�*�G��5\���.��}\6�t8�S�������׊����#���ϊq����0����OJ��yC<b�%��&��`�|a��8V*^^�0$4�y�P�+E�f�,�(K�nI]����C*߆�hK4�r��5ޒ%_3���{,��*�YW���抧��bn��k'��!��||�9�h�Ad}j�7�3x�0���PyB�%-i�2��/�7�3|�_��jaڸ�& ��A��L�����\R�A�v#$r�vp������O�,6�;9'<.���1�RX=��/�bO��2��$y���{�_ J���J�v�b$�"O��#�:!J7"�����4>�ȡu�,-�^��A�`;%�x[���q�X�Z�@S�ҏZ�A�9ߺ ��c�N7c���a$X�?uB�H�C���%L�߄��~x�ݧO�`�`����uK�FNDE�>ѵ��lE�$A]@����2	�X��d�H����>�S*ɤ��v��	�9��R�"&;��-�|	xZ���h ���������c!�$���O���c�n@�N.yG��3p`���`��-'��,כ�hP�fUe$x�U(��s!U���T�$�Ǎ���f�?�bE5���F9�0��
�\�V� $�t<������(��口�ы^�Uh��N=���6�6ݙhô��w[Q�K��VQ����	��F�:J�!���nZ���`$�0���W3��%����~�����D Srh}���L�P(i��w}�_�H��5h�P�A囔�;.�����\빗�����ϵ�;#�(K�5o���4J�f [4�
z��{��燱I��S&�����\~� M��f��Q>~��,a.�n�GaMe/ɘ7��Y�D������Tq8uG5������'5�9���A���V �>�CX��(D�n�K�iI~��bH�p�	+���(����?�*C��ֲɇ"�N1W������G4o��j[`äTf%vL�U��H6����h*X�]���ǤI�(��% J�Ŋ���"&Єog�r'�o&N7=�Y��+�7QL��6�@�j;�6�͒��y��ۛ.�9�
R�U37�.�wH*���z�bQ�_rƟ�{��5�@�o�H!�ų�~�x	�<c���O[��@�����+Z�����y���V��ִ
?�lB���(Q�c��pN��֦�1�C��.L1��g��	��ׄ<���r.,�+���sƒ��L � ]}��g{*D|.if+�~�@+�S072l-�m��7�ĞR6Ps='K�1`=R�z��8�[�QD���Ru"�5P�7�i=�UT�O�Yń����<>�m�o�+}54ӌqy
�h~�X�����*����_���eN��E����[�m]Ձ^a$r!�Ҫ��b��(���j2.�z�~���{$��V�Y��k��SBϸ��m1u�>�#��C '�̸)��Z��� C�����1f&:��֩�a�v���~���-�����#H幰�ר�^���vpJٟ poܧ���������dAw�b���[s��r	&6�������gδt]����tlث�X�/��QnʤR��gv��x;�rL���
%�B[!��\�f��.��("f�����N���	W�I��:H�5�[��2�����<�b@�ww<��������0+�0%*
��`*t��0��R{�{�"2�A� �b����Cf�Wж}\�z��QR�d������zq<n�O(�@Ϳf���2VΟxY��87�A���\�q���j`f�U�c��ƹ��f�
i7;짍vW�[m�?z�hZAT:�MG� ��!�>�~���*5���ъ���8��k'V/S8�m��r�S<+FR��5��ފ)� ��8\w'<�������a�J���������^��L�iS�V��P#�a/�3+��<��?��-�H/%R%]�a�h����6RFY�{��Jd;tGܧcr ���5�6�c����h�|ɩB��$��sʈj���Z�M`��y1z��.�p�oM	<p� ~�46
�Y���N��j�D���ݺ傇���ܤ �`\]��66��@2�/�����x`�N���4A���n�y�"�i H3*I��4����#N��c ��7'ꁚ��k!fƀ�?�ŝ`?ۮ`�H�R�쪺�Y�v����T�S�и�q�X��\�x���x��gX��R�Y�!f�X�f ;(%����઱�a2�X:�9�k��F��1��j0���J�r�P`x��;]M�5�����,oq�4��.=>^�6��헺x��Co���?s���e��UQ��ʪ������b�wDyGY_Q�m��9r�0��k����.�ScQ/�J���I=��鍴�qȫ�^�H��F�U�{iz��Y�t��f�,cʨ�X���Lx(#S[�Հ�Q��t��)��i��/��j��Ӄ*G(`�dGK���?���V	
6�(��`K9
��M�i\ʫ��2���zBaU"P�Z��D��=��/���j����=x��G�CEQĔ���(�$���id]	�E�nM/S[�$�T���o��C�{m�?!a�I�S;jn%�n�I���h;.4�#o��6�#<�L(��fs��AC��9;��b�*����j/|@���ԇ�	~,7�D{
��|��3���X��­-U�oa�k-6I�
�l���"�+��[�p������)lB�{��d�f��w�����$��Rt���4�?d�Կ�T^e�0�X�kDi'd_����}��\��#
'����9�1��&�I�q��E����1�:��%%�#�6�E�̬�,��v�I}�zZ�C%��=F�ț����\J��<k���Om�UaW?zx����ͪ���:k�oL�toZA�]���/�c�����u4]e�N]{�Bz�"��r��ּ�E���[������ fJd�tLx�!=cP�N荦�[JH��]�Y}Gd�5l�� wS�x�dx� �f�c�H�l^�'Ne����j�46�Ŷ�M�%S�aȫ���3Xw�7���uՑc��a���!����+<&����������D�����V��.��C4����<�ǈυ���Gp�zp��Y$̈bu���'�����ͦ$�l>��k����F?X^���Y��l��3�&��C����΍�)���g��������4�p�5s�@N��)$_�sC��{�WV���E"i9%z"Z/ی�������:X���ѴV���ĩ�\�wu�>���J',Ι_}��h1��.I������Y��s�4�ܐ��r
��P�����a0D,s:�^e��U��
b��PBg���ip�������P���
@Gmg�ȯK�vv�ڝC��W�I$�Ց٩�����[���i>��|X{��x�2g�?�����k�L�P��f��Pt�U������Rh0~H	�\4n���TFkuzp�9/{Z�G5M��e"��;�mM"kʿ�G�v��c]a�����R7�v-iqy�U���_Z�l�u*]^�A%zN��0�۾:�B.�#ŀ8*�l Щ�f���L
L�~VO�Ƚ�������Bj-��X�B�!S���F���ځb�Ӛ ���:��*6�E�@����7��23C��D�c��x<�CN1Խ	�R��Q�
/M�&���?;�P ���_�HmS~�g=�k�l;"w�H ��O$�Wj�Ui��H��\��f�g�F񤜻�OͰ�nu��G��#��}���|q�j?^����ש�nB�K�# �����'��+B:�#1anɳ���>1B��H�M��~:QV�Qx;92/���ӊT�N{R�����WgA_��ɴ�}������}c=��C�u��[��)Gk�ל��S��?%'��/���g� iAvt�ˎ����"�`�.$�x�$�
(�gm�B���0��;#`�Q��لhQTMf�R.r��YfN�or��O��y3U٩B��U��	���'����$�p�܌��/�Ol%2�N�N73y��.C$���\Q�~ɰ	���/A��}mq���2�85>�ҥ7���e�r u��Xӄ�5��y��I�{��`�andqY��HHI��.�`�m�=��HH)��>��jD�ԷA�@�һd ��qLɨp�Ar�%:�R.�(������!9��ce2��[�u_*��>%=�� ��z���Q�[n���@�WVuyLF�P��%� ���� �c�,�	p�4Y#mT?�@O.{P.֐���%cb�H��9�gs)��pC��"M�{,�5���R�}����2�^[{&?�>2�G����v��4��c�Cޔ��!9��a��:�EӨҘ�;ҿ�.�+փ���]���?��%�;]�����6M����2(n�����������:�u��\j�CC�=L��I~���^����Ӷdf]�sF�V���R-���0Wt�t9Pė���7���=S�=s�bB�DeN�"?����:�j����W��me����"x�3"���c��� �#�o|'�s]�J�ʧ��n�bv�h������ͼGGm;�y�p9�Ԧ5�H)9u�ǿ��X������ʡ��T������s/�X�3��I��(�ϟ%�ÇĲ�,"���K-)��,��r�5:�_��nI�n�K�1�y�j��3<�ҕƅ���1�$�cղfou]2062 �����m`����soA!i`GC4���(	������&��Gj@-�HB`��"��i���,�G�6
_ fseR���ڄ�
�A������P'cN�a
n�C��z���@�:�P_��A���$�^x� 
�Ԅ��Q�"Tp-Ǔ���w�`�?�����J��ҝ���,���P��E�[_%�ⵐɵ.{�f,��!;��Y]J�`Z�f�&z��3�h�
�uҧ����H�Nڝ��mP�ZG�'� *�v����go��"He[qE)�~d�ښ��{l�NB �Nt���?Ԣ(�˄?��r'�0��7�NG��WT?Q�YQ� �\�c�Y{t8i�v�P�؟�2۬:�O
��q�ڷ�4��B��w��<x�����C?�9J�3;���$;�و�M/{N�G�|��m������Z�W��������%�YP��V��u��3Ȟ(Yj��-ن�0	���W��ng����sϴ.N�&]�}�a%�0l�u��YLR��C��c3�W#��^���gvF�+	VPѷ�H�i��z� S0��J�F ������� �[�Ń
�t�q�­K]l9V�j����mN~>�j�:�C-Z�\���7�?.�f���G���0�V'��k=2:����$^��$��~� ٺ���_��S�S�,���ר��a��&�#�8-5R���V�a��a[^�P\JG�bO�ΠA�c�6�*�")Q�X9[�;�n&I'���U�e2г����h�3̍0N�J���LLd��VWO6X��i{�Ͻ5���z� D/|d�'Q򬔠�D矔d�;�'�Y����%@:��+���`x�-� �/�+���'�5;*b	ڼ5Qb��h��*j߭�N�9(,M<S1�o�q�� �@�pd]��X�|*̭ ���/.��U��qn6���8�4�v�xy,�I%,���H{P5�> י7K��Cʯ��Uh(ģ�bؕ:�Uk/n�#���L,�T}�t�{��`�:.|��g�
U���n�˗���@p�g���㱶w��֧��rSs���..����.'c�Ě��O��D��<|* ��%�R�)�°�g)��ճ6/�;�~Pv���?�ْ�����ﰸA��,9>��ZB�J�	@Zjp_��	���V�.���x]�18E� i�{�Oa0��\�E�Ɣ�d2�v&4܁d��'�7�6W8p�
����st��}�J�f�H��w��Jb�F����Xa�"VLb]?���(��P����vl='���u��_!C��:��������^>0���mT����]D`ށa
iE��~#���g&����z��L�'����t_��z�,�u�E��8/����5ɥ�'�����XD]4�G�	�ǖ��s���C�/j~|u7�L�Z�\���m�-1@�,6ĺߊ�l�Na5+��~�&`���Q�_�*��X������l.�Gh�@(��ϭ�iL�,�O�*�N��n{�r��-��-͊Tg���5y:�d�7��s���Z$���{�B�g$�B Mc�H�N����sIF��6�+��UN�-�9�L��C4W�kHU@�+OS��DGa�9��F�d����U�|g끆@��P�>�%{�:魩$���x$�05-���{{���ڴ�ߜ��vā߹{�W�hW�F�e��n�ua^%5�?6B� Sh%��^oc�F�k�x�Ԏσv��E���+�u/�YY�Mkc]��%�f�;>��TX?x�\�wrԄyLƈ(�wI��m�UA��/`Oq��;v�<�<ؘa��3-�	��E�X����b+�x�0W���c�%�߉����F@nA>��ES&'���/�%�Mc�Y?vt	�q���VK[vk��W��E�i����U�F��uk�mYX��n7G�
�:�!�Sz���<��v�e;2�,f�)H��b�7�����pO�<�\��*�� �D'�H�.t�"���WlJ��O��r�k�R*�k�����1�i?>ݹD��ܥ��&G������|�Nn[�0��J;��/-<  6��^�x r^вXV:s�4������9�����q8�=�l������oHxS��������$�A�O]gL�u�i�-V�	.��׹Ӣ���hI���6����>�M��fZ���-?�L7fZ�:)����|y᥯QR\W��zq��Õ�.	��|י��UWJ��!�����V�F:S
��᧠�<��Cs�Yj|ɜ�-����ط��ms��;�ƴ	/t��V�B�#\�-��"���H��AH����'�o)�vq3W��3`��9��TWL��)ۧ�2Z�a֡V��ʯ0����an�%���{CI�A{�F��h����L��u3�l�_�__ş!��J�������G��'�al�$��.��򇗣}�h]fv�BXU�Ϣnw��<�$t
�6��ɭ9m1Bp/8켱�
c]l%�y���Fʩ�p��{5� �Λ��h	������<�p��N){d�:��XH͈��D�d�k0����d>nnI�W�D+�-�>,Rz	n��+D|x� ��ps8��֣��c��zRJU��,�+���FSW\4��|#n��o����M�2�(cЮ���ܵ�;�c��`�H�{�M%SQT ��A�u�/TN/��q�z�gZ �/|���)R�;S��N��������tn	�/˫Ր�
Q22Y�4�R����@�Tc¨���=��c	��f=������I)�y�斣f��;�u���(�L��L0��Fi��g�܊��&$�/�b�z=�a�VK.�XqɃc���x��.ܯ�1
��c���e���	o�D����B��R��$y���Q��X+��Ӳ�� ��,Q���.+t"�����"�C�+*������ �;������8�|��u�t!cK��5���"��a��ԫt�,�$2�jX�˪�G��*�����;��	U��3�6L�&p'f;�,3Ö��!�����Q�S3�peM����C��섃 8[7d1�/���M�ܧC�k\���#��À�e7Qƻ������a��m9SE߅�7��PK���G3���S6�(Pm0ުu�F���`l�s�9��K�������D��b�X�/ï�d�th��	W����E���KT៤�F�%�>�������Ś��Wߕ"Qa˼� �.���T�h%��A��<2|�ΐ�tm9���J�w�G/6���[ܜh��O���{I\d�B��q{���)xA,-�!}����|)�vG)x����r�j�̯YN�@`��"}�qs{N��T��*x}gR!����{z"�"�{:&$h��Rqu���6�#(K?�~X>�H�S�c�m��2�H��)�N�`�# c2?����cbِ��b��5���� z��C�`d���Fdx���E�D�2�z��2�m@�?��?�5!�0��H��bKVif¤7O^�j6����O��
�ݲ_zb�kL04��R�vb��L��_���=8H�<�ך��7`�����p� =!���}�6��r�����D�����MY ��گ�x�N?�%��dS[dP{&���O}#�^}��՜�E�:[�A�{i0�R��f �1M��d� �蘍]d-,��挿\J���4�i�cCFd�Z�N�cg��ZOhɻ[��L"۫ݷk��IW�%�P��5�u$ r�;�w�n�y���R7��̿[�=i;F<Q֒����~��(���/�J=z�&�g�����	��N� ]�tlŔ��Oʕ�	�~�%~-�p&�\��o=H��u�C���n���T�FN&��F?l RV�W�޾Z�R���n��90 ȣ��&�z�xX����J|�}�#5Ņ�R���Bl�<���<g�HI�ߣ~�'A��@�|ęٺ`�\�d����<�"�Ȃr=E�79�e�IŬh��Ւ����D��E(�"������0)bAs�Г��8�u�`��2�KQ�<��}�#����69� 7�gW�7�~@��&P���	�Z�]��̩��uZ\%��f%hP��ן/��i俖�B�l��N�.�oȢ�����S���zs��*����ϯ�Ɵ�k*�?9`�qmh��0$�� �֛�u��}9�p;�()\i�$E�gI��\s�vf�O*˸֣�>���*�`��;9
)��M��o ��=BK���\#U
�m�{e�V�4�g�����zj�Y��� �e���3?�z�zK%�K"fX.�M����g8��\J_1�{d���b��x-��ܓ���-y�X�(9fP.ߖ�N�P�ʳKF`U����p�& X�j��������j�!��E���<տ����gg�������XW�-��ws�&D���+������-�h�3�k���ډ��:D}��v��4aEX�p���;<��L�L&V�,�g��՝��Y��Nz:B���BO�?�L����sGI�\�R�����[qэ������/��}Ba������A����g!9�������&���ۤ�ҋy�ܻ�|���������jq�c�kv����������,�m�6�Y�v敁<�zS���:�i5�fE������Y����+Q��H�_A��j�c���vZ��᩼�݆9����������n�5�ZSn��9�aq�y��B�S���7㯅��"�^<�X��||v����=#����M|��w�bi�����7,J�ٺ;�^�)���1[MH/}H��r\ʍo�����v�[�~��9�������%���*����QJ���É�Bc��{Q�_m��e4�5?['2K=f�7U7 A�c��V�h�Qb6:{�nwd���	ſ�b���sffXv5�	\\��\vhp�5�����x�\*B�t�7��	֜�z����qF�=�kTf-���>�h:"f�>�f��_���%���|������'�w��4��Tx6m
=:�X �O��7�a���4�Fd�i�C`�jN�=�6R?O����%���(���PK=�z������ �,��J��]֢D8/.��dKq�YeM�18W&{͜4�b��=Jb�������x~V��`֡�V�d���0��*oʌ���J`�k+�}��b<pk0ź_I/����1%1�D��H6^	�!Ts�ܯ�u�f��{������S��<������<~�Cz�K�~Vߋ~/�
���8]�/�	И?h� $�8A{�E���$����iܳ�8����$/k�=ל�s���?\�ů=��pR�3p$y�O9�U�Ym�6�'���t��zz�C��h�<�ԑꑌdm�y�n���"DlR3\g��F�c��H�qB5���C�A�Nu	�)3ׯ?O;.Շcz�^Q�M/�<=~Q�B�[�3bL�8��Mg��P���&�x7��y��:h;Z;�v5�m�x�ˋ� ɺ$�o�*Գ�#*����;RJr� U�F�sp���j�m���a���	�e��Og0Hr�7����橣�4uI���)[��(l�����C�;��:���k�A�;z��h�O����7�D�O��T��'���p���#�aZ����j�m�A�O�h�1/]�-�ͥ�����@6֥����t�����j�� §����/VVxd���fb���,H��+�>s�7�,�]��_?��wt��2�ě��G}L�ߠ.u,:��㲆�%*gY���!�B���:��Z�ޠ�x�rX\Ȯ6mJ�,����;2h
���+߈BƑ�?�8gq��[�/��Q�`���"���N]��h�:��Tb��oP.{��2e��D�_���|J�*Y���$:i���t�)�.�� �i\S�◂�y���.LJ{��}�O�So��� ��/@b�J���O����sa��	_w���;�'���i���&��B/R(λ�{��,�a>�VƎI2�ґ�0�Ɂ��e��I�M�-+#6�q�.�{���-���IO�$���h�C���#�����̪�s���7xw�$���{���Ӧ9+H�$��zD��'�?u�'�!"�qI H��M �m:vbuf���Yb*%�O?Ib��^�X9��jjL!�2�f��\��L{$�s$��]()�M�W�|�;��]������i�KX����e���7Y���d���1�fT�W�;.n���t���w�׍!v�@;:2_�,�����p���@K����e�#�>�_}��B5���.�u�܇����fͬ����<F�}vW����� |egs�4i��q��p&ȧF�$�U �U��31��#��h&|1Q�_?px�~��n�er`���<* �E�a���?��n4�X���(�\Nx��ҭ2����;l抵r�y�4kl��B@���Kz����F�&e,�@����diy���;���w���}�03�8�[%�J���C� �P����A�/LBăf80�+t�Ϊ�̓�������fq&nJ6R�XO�j��{�Ӆ�zBRǻ�wle84jn-�>4��]��u�0RM����C�2���5F{bl�M�=(j��W��buЭ�3���qm�U�Ɨ�����l�dY䗍���a���6�l?���/������7AH}��������T�Lg�\��xꛟ	^�C��.��x�q��(?7g�SqU��O�:za��Vd�\9G;�?Huy 
!ܣVNa�Τڠ���ޯ��(FtV����Y�1��Α%,�͔t҉��"����BL�ln���2u(gv4$S`d٭�t��:��姾>2j��!��1|پ1{���n`�#��vW^a��ێ��,�9�J����H\Z�h��N|�e�Q.������c���!Y�@t�����0t��ty4T��c��Ì��t�9�Ӿ�萈Y�`�lk�����h¦�	,��hl�B8�A`s\��C�< {��WcbH���p�|���̽&�H�=�JTр&�V�+(8뎜���U�#������,C�z�>�Ж�/7>�v&�r�K��9�5��x�͛-m�Ğk,�#��2˖I�k�J̬�&��=���:�:�ż��/|�|V���`�]�5VR���V��S����w `1te��Iϕ|�[����4e:l��0I�,C �|�������^��ԩ'ذ�K��=g���k,���sX���������Ί��Q�?�8AI�PZ����@���0�H6�.�J��1#�����,J����x�B#�[��r�8M��&��NU���A[L�PA��wM�$�p�-ئ�K-3���A�k��Wk>��p8��P
��)vl�y��PA�{����2��W�<1�n���A{��s� �ע���R3gW�i��ב�v2���
D��z�v��A��	$_=�e7`Br�q�8|�`xBs�η!���yc�/�nL6����ATe��6�-����iJ�
�Љ���=5�L[,*���t݅����"r��M�@����8���N&�5��@�y���^L?���uQ(�Ԅ���؆�s�[���Ncs��;�u�rA��Ȓl�sў�
;wb���>B-�b/��E��ͩ@�H�P�v	�����T��o�<t��9�?�j>#=��m�|v#�hX_�w�����K��1�]7�qc�.����9�?S9��G�%{�]H����9�n�S��l��E�٬�p�F3����YIA�f�g�F5���O�6?��h ���qdk$[�_Ɉ�����%��8��рt�Q+��ڍ١0X;��q�D7#���{9`/xw~��
(X�t��<�� �Q�51"O|*Ns��j�6���L��gx2Cn�ӽb�17*�1�'$���D���]�tʼ)3����8!���
,6$vL�4�ճ�q�F@t��\��q��ސ�r�	Dm�Ҁ��;��
�+���!� o'�����z 6����@�����^��ط��
�;a3��bN���m�[I��'>�:���g\�λ�td�/z昱h/��C�f��9_I��ӵ���/���n��R��X�Hi�ye�N��e�e�DS@8񵚾fq8$�E-͊}V�Q;��-qMi�B
i��mG-�?9T�'�ߗ`*��������Ŭ���z4x�$�{�&@,��`�;c�G���J��e)�O�ⵐR䗢�@� �J�}�ER�KV��ܙ<���U�2vJ��	B��n�,�=l�S\z��:�&G�����fCxL�����U;w��)�M=���=[���pN*��ѥ�)��`bBB�} �og���y�V���H�ȩk���s���a����F9�W���V�]���-͂_g��qv6p�Ì�2�&�,`� p���L�y��+��(��rR��B�5"���f��T%Tbu/���f)-L���	q�r`�ޮ���N���#�,
�����R�p}�'�knrg�P��Jꎯγ�&��pJ��lU��=N�F�I�o�sY����5��q�+�_[��Ϙ�hϬH��Ot>l��?D,x�{���/�(c��qa(ՙ]�6}G�Us����X�$���2�q�Ԃ����$HA�*�Qlӄ�u�gVQ&Y����8�H�
��92�7[Ѯ]�YP:�,-��ڈ����~F���eת�7�:�p�O�/��2�`rw]��LLS���\�^�Op(��ٌ��CKC�,���;���*���ȬY�ˢ��s�ȁy�i�8-@��k������u ʰ���pP=vl��)x�1�R���s��۽5��ѹ)!�l��I��j�8����fj���>�Q�kՑI0�������"���5-E��4z�����0�@c��m(D�չ=Jv3���#����4y��Π�Z���,���)�$	��h��ͯg����3�@�!-\����|��Fb��m��^*(�'d�m�x��p�
K�C����H���6"�Cְ��G��h�D]E�����sE�e��L촽d�rA@��9/q�V;ZfA_�og9	�C�Ac7�o
�F�_�" @�}�ſ֠���A=���ld=��R�_L�������o�X�Zyyīu�/��L-� ��c���n�<z��g)j�_��g,r) �7olF��F�ظ����HA=v�3����pِq�=����W/����`S��A]qfx����Y�O�ey�ى=���B��d��"�����g�R�PRa~���0�5/�,�I�w9��AZV�l�t�n�^p:��C��� �i�G�N�ɳ+v�I�~֭'T`�������3�����BZcj�Ds���dv[�q����q�uT�%���Z
,
����S@�^�
���g+%v�?R�f?���m�g�_�V@�����.��~?�q�:5/�,(��z�w/]�	�Zg��J��*u� ��
�&���ƃ����C��Y���-����Y�#p%*r�S�N��3�υn�W�`n�%9��2����&��9q�El���������T�>��^]�9��z�l����K,�E�lP���_&/:�}�xpq������;��-~�ﱿi��
2܏��q�)�>�|�0��e���<̯*���Lh.ZE)I����+��8�S$�����2�y����$iӛ�.~R+#����t$8~�3�(&$�p�=$�6{~[' ��� �{�8��Ae�M����2�$�6=�J�q���=v)>4��I ��p��1�jHS�ҙ�E2=�p��Q<�%���W�>/%v!怜N����rxz��]��O\I��9�'����A�&�V@|�b=f0� 6 w��OۼK�� ��l�g�.�����e �a�0�Ϥ ^��O���.�۹�{��=��W��g<���=bd�rWA�h��t�QyX>y��T�񔄰�A4{}j_�]��O~������G�����9�L�!0�O$����x�+���O_�S��-��̶n�:�����U��A����5s���5*���z������{ʙ>�K���j�O����
7�1,J&���к�����4+�k�3#��4L�Mm���˪ur���W�q� ��#�*�\��e��ާI���|
lzOj�7\��j�2���d��Qfȭ��F��ftն|�峼b��"d���z}H-'�T�AҘ �����z��"B��r�c/�,)gn�����fdlrc\x�=8�.������n2��ݲB���PE�uZ�pL��gxg�Hy���н�����yn�0栘}I4N�h���R ����l~ \�|T	��~�Û�-�d�e�Z�(b�1	U�Q��D,��{-�X��M���ױr��C��IA׎�9s�%�nu��/��Ah���$&6�e`���	��هvI��E�_��ͦ��%��D?P��/�>���
��4�e����r )�3�	��X���_�M�RM�g^�+?�z��R�C�{p���.i�Ս-�ӗ���m����ͥZGm
e�`�����6�=s���o�7EϊVyw6���V}EO�T	�ګk��WӢ�(��:����]��/���Fo'�o�#c�eӬ���8?$ڸ�n��N�7�����-ނ�#P;���d��Ĥ��_ӯ6O1�\&`+�8��U��C���|0 Y�a5�.�3_/YF���-����oI@*�`��8��yi��V�)���Q�7ZP��54K�D��4�qF�r��@�ZѤ�rB \u{I��}i�S�9���0�ח����:���.jN��#�r���Oq��=kHx��_0�"�@�-�~VbL�O����F���YN�&�&1
�=Fdycэ+E8�&�;�A$)KZ.`���/�Y-�︊�]�H�І���صK3�-M23˹U��Q���Jɱ������*���C�с=�p��w�DԘ���ޙ�Ͽ�-��.Y�_��`Lޜ����ݼ���������r��c�\#ЊM�Ș�/����i�`~K���}8iV��1������ܡ�17}�Q�-C����,`��T����wa�z�#Y��X�'�x��4��.m�Q�Ğ�E�a/L#���$��Qט����@�Y@�!߉��@�ĝ)��4��0�~ߎT����ݛ���NZ[i�!iM��dmG���'{�G�l�E6�U w�;Ώ�L�����$��jL�+!��i��>�:Qx�i3��Ysy5V=��$_����#b��B?h �ε�,� 9�A�Xؚ�zѫ[U<3�}#K���7�Nx´�	b��r+�C����}0�7��N��]!/�E4����u#I���s�W͊���3��J��.�p�\��d3!��f�R���W� U��8!Ě~�(��;�|�
ems;�Z�c<�p���d�_:ߥ3��6(#����"�2�Sr����4Akώ �6~���>�M��٤!�0v�Y���,Wf��Br�q�A��.+���򮮉���4�a���	l��*A����� �V5�����i���,���?��bq�� ��b�kn�
ׅ�y��+\D[��(_%WS��vC�p(_�lZA�M���$�r��Pr8��W�k�	�;<'`Lz�ڥ�4ȕʝ4�<=e)//�ƞ@l�5���\�/�Ւ׏H�>��#��V�����o��h���>Dat������u��G�tW/4�f��'0��	�	ǅ�$��ɝʛ�u�3�b��u�{O��o�P�W�@P��u����@�
*7����I2%����`H�����Jo�����Y���t�&|cFE.7|��1��`���FbcZ�{��Z�J��]e�~����']���p�5��?��CuLv�^LA��r$�d0(�1�f�}���$i��52怪~'4����O�gwM�Oi�$�� �!qؤN�J2�5ݢ�Y=�cV�!4��@L��A��E�
G(��l��k�����x��n'���W�4�%Ql�##��s'���ڬ�k&�AC�5΁���i�]Y�-�d�T�xxmٹ`~���L����v�~r��Zʧ,���1��or~Q��k<�?�ܵ�8'u��R#/���%=;*�S`L�l��"��G���@!+�ʺa}6{�*��6��#C'4AG�N�Zf��k�xv8��_ȇ���m
*lkT%�"ԑ��`Y���a�c�����ړ=�ހ�~>H���0�G��7e,t���w�6��ʫT���� p%�>]C\�ӈ�d���5~��j7���fSC�Y� ��	���0�g�[ٖ�Z3��q�,f
�����������R�W:ʩ#G��{���G.Y�����'��[������)#�f8R�	EgC҈="�F^|~4�
(}'h���B��QO�r�ֻ��`�-�$����� 4V`�LQ����Ѹ*g�-1��0�*����3Wʚp�m����v�~�w+��E����1P{=�_W@2"�'�j&��3Ll��4�{m�/e���/U�zal!�ST�_W]a*P��ϳ$q.�Un���f/x���&���@&���U��ݹD��jw��,�H���"Ȼ����)���revJK��*��dw����?h��VU��e3U�w�E(�S��|p5��6^\�q�I|�#�p�XߑO�%U��_9�j��W�����YUW�܄n���^����82�����gI�^o�����-r��;0Q�q��l �&�;�%!)��������%�5����Y�t��.ٯv_�C���T�P:�|����UTe��74��&3wH�M�8S�L�ۉ�6�Ӷ@�����vp�xvy�����	������6ZP�*s%8�d�䉨ON���S\kFr�*�L{�W<���
�<&�=5 _\��%�����U�)��? c�t:�U��Xt�����B,��8�C;��wT�S��l;�\j�k�R�R�eT�����T;Xl+C/�l(Zܲ7��?�9�}�)o��(�a=�n�~��F�V_^◦��ê`���9�����g�.�+�� ��ƕ捑���|3����bJ�bI��o� �yVlf}J{�x5B��A�l%l�����vo^xi為|�<��6Q3_"�r������P�L�n3��z�,�z. r��o�2�0��oS�H�{M<`�M(�xWf���!�Ui%�
h0x�� �#��u�5hѢ]�o���j6T�Z�y	{����	M��1�cP��%����¶�Q��׎fc]M�g�S�?V&����(P~�I���k�5���IA����x|�:�[��9�O&���T����g���n+��~��myf�O��~����C댫�鶻����Y"Ûy"� �<Dc{��!�)��z]XrR0��[��е`ú81T��Z~�QnA~G]�e� �z���8�!I�����t.X���_�A��壁^Q�q7� h��T�*"���b!��o�7�����)��8$+ȧ����}�v"����Ƨ�9U�|rH�q3AaJ3������Cǰ6D�"R��*�6^:N�yj���'�x��\���U�v�8�i7^����������B�m����~T��{?�b�jg����92��l3I*d�P0��H!7T��TBOKg�����Z�Tr���ڕ��Ai�$D�)�t���i	X`a�Z'��-���(��x���"-�i�"LZ�N!l��=0^�'�8_l#��{ħw>�ᨒR�Wu�m")x� 0@J��O��i�6=���O���`��"�s�	�H�d5xz���v���J�.�J	~Cy5L�X�l\������S�\���2u�ƃ�U�@^�/��Ll���A���p��%\��6�����Әv[�q-�豹�2$e���N^θ�pH�EL�׏��G�0qe��P��5�VUQ:�m���� �تiv&w���XGQ�ͳ�3/ ~�b!Ŷ���*�rO1n����k��F��3lO߁�D��'�0�,�|�>�2�\֞~sW/dJ]�}�.y�.��hV`l�]i
մ����y���z��n�o
�n���u�Uw����n0:@?��e� b�~��2Z�G��}i� �T�w�U-c�Um�����;;�x�s\�(�T� \�E�J�T�V�K���oE��um5��=��６J]>#��3�\ޢ��V+�Ɍ^l|l}K$����6�k�����|���q�T��M,�08��|��{~s�C iR�Hb�9�_�:i�������N�/ԇ7��Ɉlp�C5����R1Ҳ@;Mg=�$np;�]]l���}H��� "�R�/�~�[�(��?�H�˸̽S���a(8 �Z�˽��p��,�M ���R�f��m��٫�d&�x[��|���������g�?��_J-`��ωD
u8G�9��%']ګp#^.�����D��I�	��~�d�d�35G����]{�E�a�vTpz��F�
nY��/�5�oP�ר�w	��+�&�k�z �O�=�3@5��q^���;8>��S_0�*~��gA�@� Uy�OS�bս�����$'<��4��Cכs�!��D��%6�p�?����[_Y�@^��'�}B=�&�mH����[�p8��G޸�� �ݖ����{D�b��M;YV�F0l�b�����l�YtpbI3�2�I�;�	Y���o��32��>C+ى'����灎xEX��F���@�~"(�%RA(E�~:�� ݝ��~%�N��oV}�l�C�0�1ﳯ��D$��Kެ��Wr��m�A��<���"�<�7.��#�]�_�\KAri�2)��6�TN����@�ⴎT�{+�s���z `����FS����v�4>�EwJ����.y�F��u �Y3P��Z�]d�Ԧ��e������#+�b���K_�}�0�F���JH�tJZV�K��.��+=�r9���a����;��%��ϰG.­D��?]�Y�B�hY�x��,7�)я�UV�KK6IE���)���m���v��y��N��{��?���pԛ��gSl_�\�]Rǰ��h�tq/�����y�������_����yfC-����K�X��p� x���}_ ���L�;-��`��V�~٘ݞ,����d +t��:��a����YA�:F�6�y�o��e7����g�s��U�i!���%>79���o�<�7v�r'�Kr����S��z,�"�_1 ����ִ�p�����0۾��P1�B���=U�;����hT�[5qASɚD⩼|��P�4S��.�y�x{��M)#�ֺ[3�j[��r��/��k�{�U!�3�>p�(�;���C�wW������bG�
�p����3����YD<�e:OW�����퇠��	{�Z�q�E��>������W1eK����[Ǟ@��z�H��pOL���˂rR<a�9�QǘQ��G���]��©:�D����V����JzT�5�`LP�.�mL����;ޮ$�axn~����?�DD�X%�����{��{����dTl@����b���c�Nadpu0�ðW,d�57�![��j�����Gg����XvKy�gƋ8"��d5Um�
��\[�
6�pC�3�.��?}+k��%U ���6�C�ηȶ1��n���)"��s~ �g��gQ�^��0Z-�/uv>�1�+����I0�N�+�"��;Nj��pEE�G�Դ1 ��ck��dJ��AY��V�\�6���¶&��z�Ì�r�
�CO8~Cv}A�R!����z�O��ϙ�G~�pu�� ��SE�8a����Gh�e8��PN�"�/C�T��;L$�V����?�}�!��,o�ݰ�_�iO�J����mQ��C8u�c�P�j�"ҦDdE&D�0��}�,�u��.�/�8G��wG��/���55�g�����?�t�g�;&���� H�:/����@AA�e���R�P踫V�]� �L��8W�ym��T�P�PM|��:�5���r�ˊw��Tǂ�ԍ. ��q���n��X�?�^bQ��5����B���Z�E��x�'Pf�$��<&Y-���hg�LH*�M�^���,��6ܑ�?�����#`:��p�+���ʔ���X�Ҟ�	�]!h8�u�9�J��t.��eqL����&�B��z&�>aǒ5cr��}0C�8���ϸ���S�H4��w���o풋�	�7��4 T����
!�Ч������%-ꑅe�|u�WD3o<��E�v7�����£ں.Ƚ��/���]d����vzAzN��J�C��?Z� |���<f#���Eb�Y?�|������ơ����Dt�ܐ	�Xpav��+�4X��f��[W�A>����F�i��4�[FoT�t��0<Plp.n�^���f�R�c�ضve���uce ���Q��n*(w��B�¤��mW��8��F�TP�>�O?�n��zcA�V�R�"�^�Ѭ���.�Nm��4r�A@����\e]�W���;�7�o��s\�4�O躵��~�G������X�G$��c��'���2Ғ��/m]���K�����/���E��/Հv�y`UY�эP5]�.o�@���ŧ2���
�hzb����	r�����!��q�ٗ͗�L����8U6�ؖ��T�{zv@���	:p�K����g&^���Ju������>��'�6WG~�&w�S}_�z���j5�p�X�
�mE:N�A@؊}��F��:OK��/7�k3IQ�s���p+W5q���Ȅ<�G��H���8��Is�.���Υ*Q.DT��P�j}���r�K� �)��Q�w+�r:J�j��r}�d�q��*|���f����M�t��Ì�#!���@}���B����jI�0���u���C�ubei�)��s3F���Q���Z��'YՓ��I������E�JxYgEH�L��+տ5X�����%���|	�ؓ��tܴ�N=�
KCe�c*�z���D�Fn~�]��Ra�M����e���Ck��g3����h��{�!��v=�> �CX+�?0�Ϲ�x��`w� qܹ�H2y���hϦzW)�`�ۻSՓ ����̉R7�g>��LS���H{=f~Մa[�Q����g��@ 2g_�i�j�d��A0mY�g(�l�1rM��4Q�u�'�i�8:�A��+�9L5%�����9��K��^�Ș�$�=|��c"�a����$������`�DLj��F�	 k+P��9o�Čw�PI���j�9���-�`�}�f$�8�x�q�0��>�s�͸�p�q4G�4��T��XHya�x��?�'&|�~�vDV?C���F/�Nf� j� �L�QB|-P@�b�w�{	�J��3���\Y�܀|퉉E���;/&;�la���e����^�/���m�ظ��҅a�n6T주3����Jh�	������χ/i�~��#�x�������3��
�y�&k��{�_pn��{|����)�*v��n���Y{�s�;��&
��:.�Os�f8�?�W�P�n����u}W.�N��`Wl���wnq�XL�-vL�Ʀz��z���5�D�H;��1Y�ss|�$��(N�Ga靜ۨ�6��ƨ2��(��u�ˎ����I�=l� ���.�Eh�+z����7��Al�;vn�<����R����)s�1=�
s����j� ��Bi���;&`B�B'9��=]�/������B����I2nH��I,O
�F/�����K2e���s1�DX)�ȶ,���v)N�<��@�O�6�s�zV�|�sV�vA��iH����꛵f����_�p����\VUգF]ZH��j��}�y(m�
��n �f��k�g@�
�Ic6�"���Z����L1�c��ǂH����-��cJO�h�9��wF��ᜑO����e+�+>���3U.�����C�,�5&�A��U�-��0�Pэ?�_��I��3K�t��@�(9��y���"q�>>]Q�|��5���T~I��q[%hP���?�f-���M*��ZvD��#��M�X����P��k���p�i���X���V�5�X�b�7��
YV�p�Y%t��Ik�L��_G�5�d�!�#'2Ϭ��C�����hա���2
q��B�Hc\��mΌ�8	��mOK��Je'��7�i7�݋S��*�o;S<�g��u)��o��;�Z����?Q�Ŧ:cⲶ-	�u�6��W��l���J|�j$1�(:$N�m��&>��郕t�-ΣR&zs�a�� ���e��km��^TG��@��q��$���	�)�$��M�}b�(]��5}X���S���q�GAc�N��3:ZyR�z/?��T�~�ik�}P�`�N��=�����8��a�'���Y�Iy��R�pQ�����b���@7+�ԁ�ٕ�\��f��YP�ց!�aQ�v9.���hv+�fZt�2Ǌ�mg�Y��G *l�O�l8LC<�ė�A��-�5a��W`�D�~��^�c�oM����6ʀ�$��mT�y�!�v�>�-�w[���^�
hY>{�����^��(���6	'����W"E3�F����է����W`�����D�n �**�uk����S�"3�_�~��&�l��bL��M��ڣ��#/�Hד�d�}P�j���h|kh��t����pC�c#FXa${�@����Th��ĥ�F���4qH�۽�.�v7�Z�S�$r��O�"ɦ-�����q���J�8�C���%����]k.�mݳIrx�{��!�l�יSz��_H���`��(}�S����# ��v,t�rPr�)��Lr���;I۰k�|�qyh(�J
�Q5�w�H�J���B�/w�T[����vΠ����f
$�	�5��|v�Ɉ�t�2�t���>�S�:;��`'�Vi5��~�0�~�^^������=��b�1�%��d�f�l�#�<Я2�<(�m���D��2�?�����W��C�6�f�f���b�,�E��t`�[R���� ���Ϟ<�ҽ��{.��������:�R%c5tG���tN��{8�q5�94�D��]Ȩ��������v�G"h��u�C���/mv����-e��� �Z��v31[�%�:��/\tP��v�_ʄ�Н���Kq�ְ4��N�z�ĭ���O7pc>�Rx@sh����ގ�W�х��ÑS9�w��Kq2Q!0���!D�h+F��^nl�B)U��"��'5�+a=��4�yC�nRԝ��"�y-T\ȯ�f5��@���&n>Y�sGL�;�	��i��^:>�z���\p��s��$�2�uǬ�j�o+ǣ/vNH:��k�R��)��U��sK2������,A� E��4�TqP�3$�\}�t�0�K���H��^'"Ye����t��y����AlΡ��� �ћ2����%i�z���� 1p�� tĴ$}-�x��Fo����aK�0y[�]R 0b��Y�ҌDc�0���x��W����a�=	@��,=Q�4�*j����c�r&<
������R��-k�| �C��VB��"�Fn�d[�o�����7����G���V����P�a��ѫ�� h�����&��ƀ^� +H�;�W�}��٪L2^H��Seg��#�=�3��6s
yE�D5:��Pf�Lv�{���G�ȱ�>��q�a*)�g�n���{����H�q�%���1d��S@���a-Ӊk9DOS�� ]�V�y���]A@D���T!�o�_yG�8fZ��L��e@B��B��e���h����t��~
t9�(��������}YF>�&����}�M̧I��&$-�IA���+������޺�3��m�Ԣ/���ϛ���#����R$2�.ّt�LLg��*8 ������:�F�����uD�q��`�Dח䣦˟(�Ș|����bw�Ǚ��6���8�e�$���[��gd���yid�`zlr<#7��,l(R�b���6,�a"�y_@�WW;� �
X���X�I(Vq�/��2L�>�^EݽQ~��\S*ϔS��U�j�m$?�@��@I �OGIF��C��:!]nC�3J���+�Q�t T\ ����̖�<9�?��u.���T}nT8�����Vr��1���(ٜb0G���.���N�̴)�i����W�(εF����a�,`5[k�P��qÓM�j��$�=��~���?J3V�Ӿy��2lk��;��+��'牻uzP�:C>X���.C���-Y���(����Ò)ʕ���ti\N+���kIU�E�����G9D��/&�n��`xz���"���Ut�M�Y}����S���G91�qo=���a��U��9�m��@�Lj~voP�S�W����F�,�E�����÷&2x�)|f�-�X�Ȗr�_㇩�{��[���秹��^N�sE�|�M��]�%\�v�)W*ޯ�r�{�*,�C̣ܦ��`ɐ����D�SvO�Рz��.K��o�}6A髤���A��C�^49{�h/S��5��)W� �f�Ԍ�Ǧ8�)�gj��L�1�N8y�.���Y@._A���Ѳ�J�>܂�=�P�������%Q�<�n�����&6ҋ6���u_�`����俪��b=�i��n��`N
쵻�T�0>}���i�t�zt�%��5D����3LG�-!]bbm���o�q�sE�+!�Mao@���wj��b��'7(}@�"�H9Ӓw����Դ�ko$�����}d{p����Qυ����!ס+���r�;?�D�7��P.�o�q�u���^ޤ�aٛ��Cs��a{�F��V��.,���~��V�_������Ĉ����,��K!���]+Έj��b#�E�V;�����/ӥ�$iȷH"QF�ê�>RLi{��V�� ��df�B�C���s#3�gJa�ݘ=�BI��LK�v�gI�c���i�ߒ�η,�ʍr�Z�l�ж)=��T'<i~K@F�M��;�=�k�ʁXl��Z֛�=��b֊�Y#�M ���b�Z�#�W��?�9����	h��G@	GD�x��.���I喿������qJv��#��4S���\���p��fZ�6:�a�S�q�Ω	i�(�f����}���RM&éZ�j�?��j���E����@^SJ��F�UsO�(�+D��j!��XV�FB�	�+�w�ǝ��^{-H�����z�R$)_�`�W�Z��)ef��.ux[��F�r�tX�.�:�"���	�R�x*��ScrI���9��o!K�&�5���ERK*�tO�A���$����Cx|��J��B�� �v���,\08�|6��T�L�UP(��8�-g�03l�n���i,@X%RF[���Ii�If̰�?e2oC�^�9�����%�m�d�1;��D��x��蟊��3�I��X���y����O-��dF��x��B}��Ҵ��%d`/�����6줹��Y�F^r�r���}5s(�܎�
�
��p�ssR`e�ķ��8�Qć��>s����b�H��Xmm��%ٟ 'X���U����:�ľʅT[c&�C��v�;�'��vWL�[]���)�0��Y�ӗie��|?2��N��Xo{���f��8���0��� ��&�gK��t4�;P�L���3��4	���^nWn���B6�/Bi�i�A4��rk������N}@~k%Z{O[��|^0 j�S�^��ʨ[���vXzJm��6�r���󚤃1��UU{���eb�MJ.kX�@q���cb��d�]�~E�+_�1t���� ��ͩ�5��'�'S����]��3�}�^�S���Z���)m�	���?�	�w�yQTV�����v�������M�}�I�ir�I�|�+�ZK��D̈�����<- �I�C ���{m"'*էv���J�����t1��N�Q}�ܽH,E2��l�a4���9��������i;M3�.F��z���W_��.GZ�ip{� �
ѽ������g�l��Y���F�B��+d��U��u���-��|¨�}���h#�TH+js,a��dkm�繨{ؕ���B��g��״�EW�C�o[��@�>�
�)���<����χ�GCAkZ�)S�o���D�;� 5_@C���o�Q�-�IK`�U'��Sk�ߧ��ĉ����v0 b[�З+�r�ЗpR��\c��zƃmn� 's}���������f\��P�wTV5A�q��a�P�k�Y��;'t1��?���9�imjV�C���ņE�j�5C֯zX��݌��#��%�C*5�q�L���g��	=Yh��|�s�V��g��Z�KW��+L��H��-5R)Q��^dnh��]O�'C��y�>��*,��%�%rF�2m?�χ
�MԽs�I�B�'IH-�t��"��~�x;��i���sjG�6s�u��L�;�)�0Ig)�9��K|�M���A°,8���,q�l�e4�#R{gD�j S!MA�F!YX��.�%��h=�4qBSS[q��Χ�?�����_�!��U�`��Dk�I����c���y�0'6R���$҆iG? �{sBZ6v m���o�t�Ui���x�#+_Z`L�%�� ��;��_� ���I���%w�F��AZ���Y?�F�%��� X&�͑�/O쐱��=����ɀ�?XS�\��u쮅?��X<�8I|���'[6>�N���>���������q�~j���1�%;aO����f�����:��ӥvX�##$ݱ��fk�4�xpl���b��v���j�#�-�&H��#%HFH%�ޱ�tc�a@`�Y;��!'IS}fi�v�� L�641%8/�*=J�ltX
�A�,6o\��XZ���fxT@�����*������%:�J_�$���Ԏ��3�/�G�KNbi)s�O
���Bm���M
z9熓�A-Y]��aH�WP��P�M"�䷼�g�����Ƴ��
�ӻ<��pO�����O��{���7���V�<;�v��5e"�R�΄&	�G���_�:6��iǦ;��K?�C�ik|�NsG#.�8|{���7�9+G1=ı��"�����Ծ������Ǆ�r�[�� gpbLC�\��p/��$.	�R�'��2��bv��V݃J�ʨM���ñG�5I$�b	������fz��̟��È}����1#0���%i�Yk���o\?>_��b�N�L;r{�i��P��_8]5�I���2Q����*6|;�M��0����cOLf�G��G�����M�{ԃ��y�aE6�%�/[��١dA�N��h�ޫ���x�"ɧp��J)U��Ｒ��8?��L~N�[1��[�n�X���X�Y����!ʥP42���px ݽ����C>�%-E�ؕ[����L^�\`��� h�R��o&ݣ6K�����I���<K����K�������1"z��]�1򻑂�K���@��5�&�Q���ډ�8�E0-�1��쐙rwQ����\r����v<�9̥� ���,r��Q��>�_�l[1]Y�s�|-�����p��A�����lB�P("U�1ni{y�?���fz��:I.Wу�O.Q!���JH�B(�?d���f) +<��	]���I*���64�G�W����0��C���?`�^3��� �EJ��~Mbw���,�����[��b3��W]ߡ�� 
��Q$25��ѹN֌�)��ʸ�/���*�f�nד
���������n����.��K�D�m�0��qH�hJ�L:zc�oY�3r9��B�e�g���-k��b>�~ZmkBm�h��ԧB�ALT�0��줌
=[�T�j���W��*V��c���s/�ʠ�̿W��c*M�� ;��]q6�혭�=Q����f>¥24\�B�3�ć�h��g�V�|���C�yj�K�Cp���~�(���F���l��GYX�p����f�r�^m�;߼���!	�bZaU��X��}����|r�{��V��xa'M��}[j*2(��m�U�]y$��B�?�8�-�N�7m�㥸q�d}��b�ӴU¤=��<�/�"&�� i�ب�T+�#4����C�����GY=v�[������Ss����ÇjV�b%�U_fJ.�VkQ�+̙��Mn����&�(�|v0�&�t�y�>W����ܛ"��I�qU�B��(��3���j~�«M�z)[�����d�~N��! ���gVbF9Z�o�ox'.d��3�����oӆ�@��� �_U>ms�P��O����ݓ8�d�)VQ�,`���v0-�fN!������j�WN܋�ͯ�Q�N$.�rѭ��3�1��w��j`�G�Uvv�!�`�]���s��=�1��E=BC~dj�,hz�����Ļs5Ig�E�(\�n��_޺���%KS��������9`�HϪ��h�B`:�;�n	�D�
�z����}hݻFM)Ff��v�i��w��%9!WmV��8&Tځ͛�RQ�8��;/��)����Y�>��Q���l�QS�ӎ��Y6�0��b���$~:nY��9dk����9�D2zp0N}�ȸR�Y��P_e������#ex��qy�ӡd���#�X��ž��(�_z:mY���f�b8�w@��y��LbM��U���-H��4OC#q��yÿ� �M����&�eQ�N/ ���Rt�'���i0y�}#6��Bhq'�vt��jF�{�?�)�� �%Pbɣ��}�yI$k	ZP sMt���?B�ee\5s�q&$B�wD�NqX�]fh�Aқ�k=�d ��i!��0�$�l�+�F9�2W8�L�%��1���r�"��jjs�Ƀ�
@�]:vfЀԆ��[F���i���P�����)]�x*��T,K6`�hg*{Z�T��#'?�X �3��:(R6A�:�	���{� �^��@�޹K���B�΍W����V���Xhtv��Ǹ>x  7����p��s7Pβc���c����O�CO�X����f
�q�:Z?Ot?ouNQǒdN�͎�BS9"�'�B����x����r�eg��@��N%<Rj�[��׈��|4<��b�[�菈)���4�Js$2;U�
'�_;Qvg����Z��n /f�d����A[���p�N�����Vn�'�!ŋ+o;����U��|��E�C���=F��K� �:�"'!�MϚ	"�$��Y�B���ɮ2+���=̣b����>�2�	\��i�%����瀑NW��n�VG���"��XJH*=�܄�?�-�)XM���bw����Z�]a@4:^�(oI^����Kьo�t���ف�YrΊ�Ta��@����tO	����tn�z�����87l��׎r��� ˇ�B��M����/g&��W��-vS{(xоM\ғ������~RtĤd�[���2j���ZN��c�6�*S܎���hG�q�B���g�3I;��]�̓RXb�u�r'��!�d?��")_@�BQd<�*P��K��w��Oq���>c�����o��;�9�#T�h�ѣ��L���*/�� �Dq�Mͷ2��,G���D������c9Ub�>��Fj����s�L�����c��j��_5�;�g�U@�ZQ�5y����/x�)>��~m��ifS;0�
�g�/���h1���*1W�R�Up�Mp��1�k��ȡ�GI}�tQ�{�C�N��t�c�/dlĔB���q�Ij�H���d��GQo3Y#�},�c�\�H��HY�ڙy����zK4Y?���L ���?RĔ�e6ȑ�vG�L��_�"�2�)~*Χo�yh���?���w�q.�	�����'��/� =�4"A�G2����[�[W��4��������R9�of�t?;���o��3�A�YRb��4My�)mHO9���l���ck��"�e�l9	v,O��]|�҆V��>h��n��%`�u@w�n|)q~���Ǿ�{u�ѲH���>��P�ڙ�<��efڧi�����ݘD��w�n�3r�~�N�iZye�����3����:�{���z�%�@U'�'&��u�B���Gn��N��34��l[s- �몓���B�-�?����&	h� )�P�g��1���c�G����W-Ð�u��h<�֠qL����d�R�Kc�*�CTb�g��I��n��B���ܱ	LJ(�d<� ��^<��$�������YU��  ���ܩ�Q+g�c
ꌖw� (sQ��`�%�z��&"o<蛇)D�?�\����()��Z5�o�X���"w�!>l�����������v>N����;9��)�[��w^��i*����[�l���'�Bhh{�$$��m���{2�1SD��0�\m�_�0�<s{�R���9�?�+�OD�p+B6aE
���Z�٭i�z�������hh���������Q�(�(��#��s���SU:�0?0�k������H�{�ax!7�	JD����gV�b�q��� `�=���4ނ�*�1I�f�����FNG*��f5lճ�[7��� �����D�M�.Y�aMp+�(��,�QF)�m�U\h稐P�ʲ:� \ӧ��÷��U�erQ��txǐ�V�?!���+�����oq�����
�^�_7-&�����a�'z�򶮰&�)��8֧������N�І:����S�z�$uZMG�׆��eQhP�s�*w}���Iu����o¿���9Pl������=����nj�ߓ��u��b];!AZrA�Nl穵F6a��,���	]m�������K�?�p��n<�b�X�,�c��n���T.�*��\mT�i`�xG�J�
4���ٲ_���4���k��� ��=��ù�.g�Vg+���w;�ܿ���K���Y����n�up�J�ƷJ��'��o\& h�`��' oO}�Q�t
�. �o����8��_]oC"�p�3�q�	=�Ǻ�V|A�?��K��B
���@J�f�Uh�8gς��z�M�o�n0@p�����.��svݎk�AxFL[� �p�5�3�,�?���hv[��yi���Y�#�o���H�w�#R�?Z;y�)�:Q"�E��#��	:X��`T���#"�I�_J'Br=�ޒ�Re\O�����v�׏�]�K���ԙA#/�I�Z��A�\��j�am�C��;A(l�1��?24ӇnGzc�E����2��3�?�Fr�4�贘�(�(l��3N�e�ߖ$�A(ev�NU6���(�m��G���������(�C�2ǒ튥d�\�tR���W��W���]u���Bq!kwiW�6��ہhW��y#�J��]���T܆��\���_� H��Z+����1�_SH��{Uz	��tґo�׃�*����x��쳶���0p\h�$}���� ��~"���N}x.�֊�n5��ۦ�~L�1gm��U�ב/]J�;{�������ݻ�0���7UX/�"Jŝ]�g������� ?�8]Bb��X�dƫGL5{Db�aU��r�ఫ����K��B�l5�c�6�+�?�l��y�
�+pƨg���_�~΀�0�SX��`�ͮ��b�ͯ�0�����̙ܲ��0���=��:$'��Y�=��n,F���0$g���g�������v��������6	4UY+��}.���x����<X�6�d���<���� ���A)����(�( d�C��X$R��0uix��q�JC��@j �Mwx���o��d)p��Il�c��ڴO�Ŋ�t
�������	M�/������I�mߡ���ֿ:6M�ss�c�bm9w���6!B���iqM�ĮT�3,��ĲNי�/i�F%�`����5iێ��� կ)�ڊ?}(8����TN���c-�8<�D4!�3H/�#L>��貭�,�pIi��ټ;Y�Leb��,�>ƞ.�-69�q�+a�(�4��%=�x]|���6����S1��%���<����2X�e۶�5M�t��׽,W�w�:.R`�rJ�ޕ&fG�㵧�KR��8�-(��V�YP{�pR 	��G�sUf���~��.x�`!	�x@|.�����O�j��.�^������	TQm�]\��l�h�r�u�c>H�}�fU?�QSe5��=Z���	Z�L���P!aA��4��Yj����2Ooy���;mrcl1����%��<���_��y�	�f@����)���y��(?��Y�G�?�*�k̒x{�_�Ɂ`*�#����
�L�5R�Qsg�_�0!���`�/
Q6EJ>|�Lr"���� Y%��F0��g����i1��#a�[՘��J�B��SY��-��o+H��<�3{�#��XNO�:|.�:��cX�LR�ڮx?��Q>{�R~fW��h�P�Oپ�@�����7��N�R�u��މ���o����'uԮh@�%�{��h3���뀱?A���H"Դ�F��W�<�TJ����j$(:���?�I�n�G�%T��auj*�!T�퇆r!�.#7�=Xe�Eҹ�b��=H�~j���Sߒ�b�����z�i�GzYX_��%��%��@�C�Mc*��<��]��w玟`BrA��F��"첿�5�%Zu�x/������_��a��W����V?iG��J�Ґ�ZU����=��^L�ST "ς�r�h�F	J����yӵ՗Y�Ϭ��(�����#!y��g��]+-��ҍؠS��O�]^r��U������Z�h�ϣ�U,���z�-�ऎ}ka�����+���9�Y�vrb�ҳ)Y��a�0J���`[٦δ�Si��CH+��{���=Ę�+��T��?\�*�|��қ�+J�z��WTa�� C�t�ٟP����X?R�գz7�܄�>{ez��T��G�W�����������Y�;O�uq�Y�偔����𿠗���|1�n1��{�]���l��ʄ�"?K��YQ#�f��{�3" �%�tc�6 ��g��]�enٺ�f3�L΢��O���d��m
];k��, �D�́?�]�wz1��G%,�<=��B{e��T����J���=���G7�eK_<���n��)��q�l��;Jm�Jb��L~4?�w�'蘦� i�\a����_�Fڝ��^5�[Nj� �vk�I��(��9�7�J�4�&c��Ia�#'���2��_�.w҇��G��3��*�f��`�	gأB�-�l��u��aCw����Y��H��C|�xGY&�q�k��U�]'��rP~�
�{�9�Yg��c杮�6��2�]����iz+��f�o4 `�z�+<�b�Ui�N����=�7hՇE��L�0E~J)��X�ܢ5��f��RY�1��!�����DR��<@y�غ��gi�?t��ٿo��^y��[V�W��WS��QC*���91�g���oFf�TAj�gk�V���L�(ꃯW���T����h��f���
������bFTV����z���"�K��n�Do�k�Pr���bEPE)�Lz�p9��rZa/3��q��"*8(����%-p����=�4�
��a/�a�/O��|��k�rm'#��4��B5Ґ~���mᬹf&�95Z��G0#�|$r��X0�w��M�p�QQ�*� ��f�]>?�3�¬g�Ƶ�CG^xM�UR5�eB��r����O����;�Tg��~ްzi��w*�:6Ʈ�7L�$"�����:����"N�7G\�g�(��s7bU�>j��W��0��B�G@7����α�t�\"팾6�c��~bk��p����7�ﯹ�a���\�"%�J�a��5՝���M(q�}����)�\�\�J�7�0��I��5Q ��N+�:�t��G�2B9f�C��z[vr��ka��!SV�k�̈,`�^ÿA�������8L��\q ��L�vR�"��$5Y�}j��İ`礩'�O�_�5X^��z�e��~2k��8TRj�EC�j;@�j���_��ܨ�2��S����>��_+adi�6o3�H�$<����wv�#����jg*�>�~��z�z`�n�~��МxZ?�O��y+�D�������>�;�����PU��}� ���H*��R,Ap�a��('�w\׼�p�ȇ��w��(-��k'L�������֦�2]Uk�����S'C+���̒��'���^#R������nq��g0z�!dV9b尷]���x�m�f�s?.����u�\J�}������Eb|����܁�xZ��A�Ad���y���P�"#�D����Ci�$�n:�XV�}��F-@g�	��X�碦���"��9�IId[�*3�1�l��+6�0�2��Bl�o�<cM�a���:Q ����λ���k�Ch���%�~�"6�'U����и��ࣹ��y.�.B�N(}yLgOME�~\������a�H�9�����c.p����T��?:�ð��V�>�ؽ�:$�|bN���4�&�-��&�._�_t܆jGY,D�N��Rl'S��QB�Ƌ��M8ruO}0|�}ǩ�[��wUxQĜ�h�:��֔�lD��e�ӱ�o����}*�̛�d=ߣ/�r�pj}��^�0��@�,����+��	��w��3c���}��e-'@��n�
'�nh��ӧUq����-��0����.Z$ї����}�S&oT^���8̈#z`'��cD;z�+}5F�[I���o�T���e��E��o3��{h�U=��b���z��g���U���v���G��eu��O�9��N�MQ�-�J�<7�Yx#��� ���Bj�!�o�+*Zif1#��C��Qo�F�le�N#"�n>'�4X�P:xsNs�>���~��}�Ӹ�4(�X�je{"��P����k����S5��K��Q�8�UjR���r� d�0����i���;V|ļT\>W�E
��}���9�Wѫ��r_+yB���̛ �/�&|"���?��1��m��b(����er����\=�`��\�#W��A󎉲� iuӑ�A���cs7֓5\�1�裪}�x�w��c䯓�W����3,�/�o�(D��j�	�wd��$���v�;!�ڄV�+R'&�d�1�9L#4`�ee���i��Z�2H�n��*/ra�ߪ��NsN�����C�y��-Չ�_{�ShL�}y�^bGơ�-�R>���8^hԐ�Cb%�{-�ooAali�yg�
�S�9ʬ&%��<.��c�i��te�l����y���`�i��ܨf�a���RY�����n��mB.���!�ƖaZ�{}���C�P��bP|�f5a[h�V���tݖ�d�4�I��=��|��D��B�`��b{h��Fӑd�F�����.������Cdƍ�6w+�i��;��kآf����&��<�K��I��H�?B/΀�w#<;۾����v��U �y��JE�)}��q�
�P.�"HM�����m ~!���__z��l;���/��|-u6c��%@ܖ�+sl��k�q��K���r�s-�Ր�	����������I"pΤznCsp�׼;-
[�@��Q3�п�dg�� M��u��a� �I����5Cut3���?DǦ���j�n��\������x��2Y���Ժ���e��S�_����;��|��umo��Q��Z�q�Z���aVi�a~���2���s�Wĭa7�a��Ƶ+�ɋ�)��V&I���.�^��&�3}��.��g$�̴ڟc�<Ge<��(���a�q�?%�s�m����"���w�������Q�����m��}���k�S&#b�;���$��*B�D��\B����C��C���ؼy��k; Q/�͐����u��6�������H�P9���a�P6�*���_PG�M��^��<h��s�����彼��)�l�G����S٨���gζ0����4���{��v�a��O�g,�VO�������`�T�N�.���^&�ztt�=U�!iC!\�7��nN8���pI/n��Q�_�I��d2Y���L��Ɏ��ā��]^�(vq;��"i~�Fz}�<A�;/{�,������6���3)����j���@p��\G�"W�H��W����e�����@��NqQR��S�(l�S<�ȢԈw0�V��Z��{�\O;Ʊ������aݑ��>R#9��+�t�y�a�p����#0OH�F���ǚ	���AB&&��c�j�PNy�$��Q��:�ޗ��`[�0#.��Gg�MSiҜ��M�y[�j�b0z3�z����-�b2�O�n؀��u+�����/:m)��[g�8�cG�Wz���@�mn���|	����UCs��p ��۹ >�:�.�j��ӥY������5N-�Y��+���h�(�q���O!ɚ���P�{��VNVW��K=�.�HF��L�ߝ��&;�X�#��I�M߈ў��T���� 9���j��ʺ��z��d�3Ay��[z�RbƄ��-E�t��1�K��D� �o}YLk R$� ���e�gq[ o���e;����Q-v�S��u8�L���_J5��5��g�M�lC͡�����	8��L��_�N���{�'<6�-SˋU�-ȏߏ��u����b�%0^��!T���ʅ�sV��(����J�FpB��66����a�]U�p8��G����>k��QΫ�RhSŲ�rQ��Ъ����Q,&�a͙�%��L>�&��K�U�l�h]ލ6yk׻��tZ��׿[����#:�F�ޚg������ȸ�(CcK��"�#�a�F1�����S캛 ����ϟ�*��K]<�Ml`�����ª��S���ȭ2r'a�fw^Stu�$_������.c�k��Q�6��{e[��w�R�7���D�� ���U���B����g�s�5S��,�j2a��*j�{3h7����`P�a��Z�D���M���W�����X��Ӹ�yh�L*%�f(Œ��+��3ܰhO��?uI_}���[��9�� ����f�YJ֤�f&��O�4�~�^���<\����ں��6��&v��K�����3���S�rgi�jE�ʽy�s٤vg���ʘ-��Щ�7���l�;	и�&��<�?@�+� ��ۼ�f�y@���m�	U��0x>+����JE��k|o�4�@�Y��~�ɂY�0��)(fY��u��gJ���=g]�����)��X�'�K�p��5��*�j�Q�Y��_c��;��[,�!���l}���u��������4צ�B��q�)����v�?�y8��V�㩁D����EJ�6�"C�H���)G��|��h;�c���V�CX�����.��rْ�b���ň�?���i��C37��N����,*��33X���,�=X�/��̳��a�Q�P�vw���OY׏ir�&G� �X�X��1�˵��q��F^��I`-��coLw!l񜍭\4�����/Ò����E �S�� K��K�����N>��HE��֧H}[��.�m�xW�I����T���@3�O�}���3�SP�ʸ��M���[m��hKK`W+2��yΈߞێ�H�o�9��G�
��Bx��ܩN����2
��H?�|�+��:�B	��z<��]�>�(m0�����m�x�Ί��,E���2dk��m�u3�[��� �Z_���k;Z8;�v ��
�^F�3��7כ�� ��W�02-1��l��=��m{%Q3��
�	Hц� ��N�$x��V|	��bU2�I�]LhCS }�
� _��	��[)��4��m�+U+��3'�ldϭ�d�>�9��q��@{ -���X0�lRTA�u���%��Z_�mo�!�il� 6����Є�$�K�=�S'�(.�J���Q7�6�K:���;������g��-,a�����e�{�e�sGB���8d5��<�?�}c�����u�9Ii�i}��:ν����h2?qQ���߂%W�ހ�a������q��c���9�!`�8�^�w��rB�Zq8�
�E�@[�D(��M`G�3XkuZ1b�u�=���x��g�_����^L��-Ȱ5|�#�f��~�ͤн��~b)�-\���cƉ�Χ��������q�K��-�a?G����2��fX��0��[��NH����+�t��t��N��e��>׫�yt��0��P�p/�������g��������̦"֓�����iζ=�
�{V�D<~��M�-rY"�/<`7�3�y��)?2Ň�����c��cK��b�Bܳ�ȡ[U�<�Z��8�=�w�Ο����=8C~+�r��fB~��)3_��e��#����;��U��'&ع��SK;���KA(��7�gl�ECjq�����U!���w��z�.�K9^�R`]����&l�G��s��x{�r� ���Ul0�����ɇ�*��V3���I���N.��U��0��Ene'A��L�|���"�D�*�a<?6��:����v�r�eXǯ��"<�ʨ~��}1j�jɓZ���q���!�:���	���9 o��,z�e1�C��D鲔vU�r���=Gkf��EB�Ƨ�w��ڱ�n�j�e��Q̻rX������E(����r�\$�#Ԭ�Rs+���al��%��r�ؿ ��A؂��g^x9&�k��|!D��;���O4�B�P���q�й�՟Zw���ۑ�ȯvc� [�t޼�+/��R�����,���/T�D�����5�Р[F�3�ȻI�TcCQ�_&� A�)�{kYJ�#���^&�?�#4��Ǿ��y�Ѡ����`���@(�Cީa��݀U�U@��$7CYk��l$���$����՜�ҺUS�ȕ1��6�󧄞�V��'q�;�8�2�����|�P&Ϙ\�l�!���0�N��Ĥ�$�$�PE�އ�Tq"Y���Z����'ixE�$�+qgh�E�>��)7��l�4�{�g�+�o��>BY3]FL�j���c���&w }+y����m":��Z��;A(�cCB�n$Tǻ7�`ny%�M�K��� a��r��oz���<=H�S�`Y�Պ�G�yR@,��v[$W�kGf����A��_�Q�
�,P�W�p�h���Yx�/�Z�J�fh���(踆y#c��4w!��o��I�����#�H��8�'z9��w-�!㜅^"SΈ^��0`:Nm/��(f�?�7�y��biN˝u�iP�9�t5k�9SXXAjE"�ކ�:��>�	�����)
I�� Y=�8Ӝ,L�7M�a7��S�I���O� kD����s�eU�}��k��+�#�.��=e:m�G��vm�WLf
?�"��{C�;/�)�j.LE��%��r���b�!�a��	g������I��������]�u�$����
����U���Ӏ͋m����Q�et��l��~f=�F2K��j��N29yNu���e����60�EB �L�k}�?����~م��C�S�Y��^��~��~)�rAF�;�D9@
`�\P,�(��Z0ZA�]z�����b�bS�|�!�&��]<,ƍ�~�t/^�Q���Ө;�\s���P��m�I��T�B��z~r�5�� �����Jx �0�-9��ae���/�����d�d+�9$*lW�8'DG�,M솺/o j+�����!1^ɦ[ūy(Ƃs�9���䥀{��)�q�k6��k�h/���/J-�Z'�R�Vg~!!%:��yBDR2�C��#i]�) �	��R2<�*�\�����?��l���Ng��U�����q�b���m3��y��q�^C!����EY��v�v"\�X���p��S5b�����ð�謁�.?)��8P^W]5���qq@`�]�t�)O&�� ���gP��~�%B�/����,j� $���ث���.�X��[����'�ڇN���ۤg��}�`�K�9����Y����
w%�N�,K�;^����J
�qW�J�@����a�W�a��?;W�8�b+
�hZ�W �fa(p��Ё��1��-R�!
B�gv��#�}g���:Wd�����v�3ai�6�KAw�{6ŋ8��zq�C�5	���uu���b�Gs��ʪ��S�$فh��c�E'��9�0簮����g�-+`?qQJ߼��VP��.�"��@���a��p���mQ���t0�,��~��bd>��}F������`��ֆ{-eS�F�6�H6��,T�	��4:�Q�B����ط����]��WD���m_�����X*x��6����Ttgw�u��D��Jʖ����)'t�a�pu������efƛͅ�����T�2�M�w��F���RI��emSG]���Sc_x4u�5�>|}��ݍ	����`�2m�ȷ��@c��L+_���L0S�պ!�.�N���y�!�2-L7G��5�S�P��u�<\�c ٹ�\_viګ�~Ts����H_�B����r�'{�9��T���E����N��0D�T�:P%���R@�Z�%��g� �ِ�j��NH�����9���8ƥM�xZR��sh>�8;�
���R�U�H��"樈�8���:?�Ϭ�jJ`��hG�N�ͩ���k ���. t�*}%Si�;έ��㊾��*�(*�Ȁ+�Ϟɩ��b;���H/I� \rj�㟱��=I|AgQBs����}�C���	�	DZGĒ����
@���DbC�3��i[�4���0'Ӻ�\1�)W$���}�+��	vh�R�.-�}rse�W��gY�n��5�l�w; ��2�?�ur���A"�b���k��ܻG�kPw�Ϡ� ���ŧ�?��0N�D���%ߨ�R��K��?��V��d�A.�Tm9|a�躩f�6Q�`�kB�ҭ��v�]<oM�1�c~}˒%rQ����T�
���ud����� ����ښ=#GT�nA�BS;��>�ٺ�T�H�	�=�:qJUԝ�^Su�ey�5 �Ö
�d��+��9�ߋ�0�{���Q�m\T�9�<���J�M<�;q@�h}<fp�E�<;2��?�y]#S�!MF����xʳ��|��
�M�,��}����Wy`�S(�+���z�%zV"����%�����+.��a�c��Yըf;+�|�;��MN8�Ȍ	{L�Ϛ ��a�����i��F�G�n��#��v08%V<��1��j�4�שa��e~�7Č���1̇&�$!��}N�^ �1�Q[xdğF�� �k�ڀĕv��@sh�Mx�nd��a�qI&��b6�3F�e�_�.Urh��n�.�&U��5��y�Z�V_��&wXi�LDa��I�nD@��O���X:"8�e�b�c�"n�	��S16���m�E�uYn���^�Av)"� 87K�<����7�nuS1���e*��\âU'�b�Ư�tP �N��Qn�I�JZtթ�z_���d	�����\0�b����JzC�;6ۯ x'�`�z�� ��~5Va��1��m�=��-|���fͩ��Y7�Ӎ��&ն�X�<�y����:@�0���W'Iۙ W�>lS6�E2�2^��f��2R-^U�=6"�L�?�ĽZ�Π����w:�ױ��zRVHq)j�����7�/B96S������P�h�{�G}�\9�,]emJ�H1Ġ^���v�Z2@1�G4Z+�̕	b��*K��G���#��*�yV� ,Xf_�5����g+�Qڎ0���i�c�w�[��T��|:���Y��]��gWA;ݽ�L���
�SȌ��]a��t�� �>s���j�s��w�W����Ok�[�P�+X-j8j-�R�o��n��KƜv��)�����-�ڥ��������A�ެ9��C�$?�Օ]-�;E��e7!��j�
;�$�l.2s��%�[�y��A%�?�_<p+-��09�Û.�#�kզH��v)��O���œ�{�M\�^�ei0�A�s2T�JcU2��?�����I�+'��ۙC��Ȍ!o!Vլ�����rW�:�l'ef��0�Z��r�-W�E4�!S�Q)�/��!��^�w)Wq����ǡ?�?'�vA�\�����$c�ǉ�1ɮg���H^�0r�Jg�o�����[/�o�ؚ��Ӽ�s��Üc�F���P#�������L���o��D�ƥ�,R�iw+A�)1�
�?�2ݹ��������݌"����41�K�6t���x��u6���ʚ����Ǻ9mi��:{�<��A�>�I�9!EKey�2��I���\�c���@��Y�r#&������G��.B�i�Kڟ@�$�y�d��Z�k�	FDb@u�	�{��KF G��/--9��,)���Cn�7e��8��b��*�� ���"S��gZ��e@g���0Dv�٦G`�d�un��t���4b��S�����Z���1�Jti�7�)����.[&}Q�D���)�j'�Ä;&�:c�D:����gf�(�j�ʉ��JI�+44�DFq�%]L��)�l4�u)~C��K����h-������s��@��bv©�(X��Sj�) �fr��_��O��£
��c���O����y�5ȫ��f�ס�NO�� 3<�Z4��T#�wh(+x-���d~�d�zO�*�"�7��Wi Z���R�޼��H&�%Dm߱3�������G���� �-	�1@��\ڑ��5�����f��;�Rjrn)!ʮ���l����}�4!9��ݏ\)��#f��P�Ť՜�M��p� �� 
�p�5)<��X�Š�џځ飇C;�^�TI����XH�]ӽg��<Y������ٍ�E{�k.�Ӓ��ur�k�*e�(!�U�ODíE���i�,��k:��
�8�JT9�j��<:M׆f�jd�gUW[����N/�x��a��B7��Ab)_7��'?���Q�4���ka"O�2T�$��u�)ݐ`d��?D:���S}}�,��u$lb2	�2nNU�~E�{�����0]v2N��QM�̵�Wg�3�C#��׀\�[!/#�DF'o�;"�K�,}|�(��/��E�D라�#ZX�t�O�ll�s�<�5 �ݭ�ᐃ�`�)	����xE� }�M���3�BC:qΈd3��դ`�k`��N�6��d�ڱ�f-����x�����h`�r֊�'�ڱtZ�8#�5�$'T��nl�]pp�o���I�l�h02���.�ϝ� �ap��O��iO�����M.s'lJ�J���Y,�'��3�/����~"yn8��>!6��3��B����ŋV�Ob��߄)<��Cl����M�3�t����4a�w���k�0m�7F�~BW�'^T	������1�v�n��4�lz�	�#�ke���.��*�����J�~ɏ5n��.dT$�ſG�~nb�X'=4&�����[ZW�ZWsZA�;Ŵ�djξq�!ۀ�6��r-�3�s��*����~u�B�>���28
�|����]����R
�0oyD�]�}.K�+���Fi`�㔁��6f9�={��6Z�:c]bN|�?$[�EGAR���>ih�e�g����aK<�۱�t��V��ү�pc�Ex��q�G�[qP����B�'0�{G7ν��n"À��mK�l�{͝wl����E�nah�`Qd�ro�8@�<���1�v԰J�ЪAb�����WٳYx������%W�bl��Q�cL��)���T} ��G����L���"=b��oy&�$����+i�#��ژ�C�:����;9���1�Ə�\L`�6%}��c�ܚ�q��$�Je��J������A�;�a�8�.W�H' a32�Ź'���kT-�ꁀ����_�}
MT�bJω֏����N�ȹ�p=�(��(�3���j]�\S�P�4�Q��n��.D3��Y�?��"� A��: "ծ��^�_i�{�)�jf�4����=b�ci�c�k:/Fy���!�	V�Ӱ���4���Ԑ�,�v�
�޳�#�	֒��Q�5?7��~J�?l!.3��&*�������-{��a���0A���`;ׁ����P�T���>n�R�Z��2���$<d�d�����T.����7��.���e�졋�% �a��jbǌ{���ʂ��j� ��L�V�my~5�	^��I�M:K�&jяH.��=Ŭ�.3Z��%��
ŻX-��P�<?�g|c�i
���q��p[�!���QIg�˔@[�����Ҡ���#����90O�#~i_1�TE�*���V�XA[��!�؁�K8��p��1�Q
R"�+7�\��Ÿ�M&�X�O��۳5{*��)r�r@x�4�`��H�6D�ڨ�z2x�	��u�f6>.��$���� ���;ޖڸ��컄�pXv��S�PC��k��E�+��Ļár��cG��!�Fb�餢8�k#��&��u�m�[#��6CI��x#�������/tu�����8�2<���������� � 
T2�7���%G����sG�5�Ϥ�X^D����(e��4aGWX��I�k~=����]�z-k=��2]w�i17����;�T��n��]��F������8����1��˱��ZR�v����.k|V��¹C����<�m^@v��O����Q����\��A�R�X:�s�SI3��u�(�
1oY���2ɯ�'Ǟ6QrS+����H��H�J�	P�]��k�]��9�:U�6<�?��Q�{�5�������e�ܚ{ŕ�̬�W�t�u�@���Ɯ+ �2ݣfTLJd6��#�	���Ú�c�k��mdQ�N�����W���;!Q'�I����^�8
��b�$RM�*A8b8'������_����ΐk�����@��GO�l��;�J��y��|9b��m�F���)ʸj!B�%���w�c��)�>��3�;_3���?�N�F��5�$���o^s<��ςzȧs���$����B�Y�l8l�)�AK'[�����j���J�W.?u'ă̫'�gq�)2!	}%����ܧBc �9{�N�m,���)�p.#�%��g�|]���P*]mNX���˶+٭�&�p�I�4tOWzt����bm:5�q��NQ��ڟ�3�dPsiU204G�v�7�������R�M4�x���C�͡����*H�|��^�g	�P�DUq^�q�@����G��I��Q�/��C��:�P��x�wt�����?�"�/X&�#D�}���-�4��ת����|���E˓���/�%��(�E�SΣN<��ˀ��1H9�V�3Sұ'^	�m�I��`��=`�7���f϶ߒi<v��F��F`k�����u͜����9��v�����ZSY�ʕĹZ��2}ZL2�=�7H�d�^X�7IC��^#��;Q!u0�Ѝ�� � ���E3w���(m��r �h�`�*�Z��Q���>��T�ke1Ufz��/�I�W���L�=�~�eT/B؛�-��02�b���Y����tغ�!���\�+��7�V���1A\^���3�"�v����JkA9�!d7�Z��+"�q�<��'�����W{������kV���hG	Ck�O�p;���'�W�
^@'���\\��H��tB+o]+���3��bٵ��à�6���x��k �,�۶�G���!�$���2ʇ�=G#O�D�9)��7�t�|���Cm�wx=��Y��hHQ`��jk���5� ���j��M�1Fx�R��V�a�U v#T���E�T0k�-ͅ��hC�����coԜ������j�>h����f(�u4�MU��A�����1�hZ);E�d�]��S9���>? ���ι��!��Ň?RP�8�l/�YX�׽�i�������	^f��k�/� %F�r9����ҟ��ה��@ '����u��>fw\p���j�V�x�����ť����������)`.�q��O�S!� ��2I�]����<��qq�jG�=ݖE�@��������a{��A��u�f�O�1��S}Ғ��%rP���y�������A�z��>ߵ�ɒ���<�eA�Ͼ�,!�6���T�v�� �M�ћ����S��/�L�zA����Fo���n�Ԓ��_Pmnl�C��Q���M8 O�M�Sk23ڰ�>��p���bY��W]�sT��i#X�ea|�\�C�\��~��^�)>����V��oʳc6��:�a���1چ��yDyɛ=�YB��N��!O�ƀ�����p��i �z���ইSf{D1�4z5�р��6��X��*t�B�kz���U�:�!粊/O�������� F+d��)+��@� ���~�2�m���/�JZ@��&�PE��KcM����,�pt��C�3�[�bv�c<�z���=�ܽ�˖j{�S2@*�� ̋a��)�1������!�4����`�����s���?1�sgGS�!ٷW!�A,�����y�Q��!V� �`���hXY�\Ԍ���c�W	2�pA�ĕjx��]���;�c=�b#ײ�ӟ��Q�N���z�g���k�ؒ������*�Cp׎H_�q�R���r.�Y NM�pY�g@Ȣ�w�m@/��S"�kY�ջa�5v_�ද*��G�M8�Z�Ѵ�.��p�� ��ÇۦfEK�Dh\�GJv� �X'���^�"�+�����eڪO��3�w#�xv�8z�FM���C��A�p� �3��N��
�}��=	fp;e��y3�����B>vIЅ�+q�he�y�"�E":�B���ϝ.�J� ���@3�́щd���'��_u����:C���2��$Y�Ɂ>��� ��v���?��>���!���P��6yt��EYNEL�|À��Wl'%|~��2{u]R�n���Jɹ�����l
'Cz�����4� E`����mfd���q���4W8�Wc�	��s�_^~h��Jh)ʠ�b�MO��%g�����-���	�(�H\��y>M� D,����ݿkAW#���Ж6�����!��Xw������68�Ĝ��[#/�?SSf ���?�΍T��Mw_6��2ƃ�9�h9�����8�Kc��!|���mF�'�y�TQ]F���^�{E�aD�;#�7F���UJH�h�,,:@�&��砖��6{ծ�1J��.��c�e�+^ة"@c�����.�7a�
/���P�G=��`4�FCm���\�f�%`�㛷��*���@��0���8nO٩������sc�x�{$�QT���?bj�}�;�S+�7%]��bH��������x6�=��O/jI��d�uz�pOd�q|�O�ݼ�i�=���d駏m�,��/V���͢�[��ع���^���^�2�d���Ȩk&�+��|A���3×�=>��ޠ��`��$���C("6�(�P���,0�1���S���b-�\�s�Q}�=��ъ�<��}uN��j$�����N89��]-�	
w� ���8�^���z��"���Ӡ�Ű��jw�+�V���QXBf�qih���m1�	Uy����Ж��eIO�e-�<"/�=th�,�rG�n:8"W�!��+�̵���/��$��<sW�>���=B#�p�ɔ�L�6�����Zt�`K2F6�_��u�5#n�[���+�*��8�0s��sEdۯ����e>�an�J<4@$-��{N]연���	�b:8Բ���y�!��1ߡ~҈a-x]����Q[�!��%	��:��c�Բ�#E��>�WT��mf��M�Ϝ����c�?o�����I:��0d�wɅ�x���d�N�x��6��������𼠇�/�0h��Z�.��"����l��s�I��g�3<v�dw����Ud��~�����W��zĔ_��<������+�L�"������ܿ][�AL�:���k�Z�+PY��j�+1�֍����Ĩ:i'a��ϙ5{�
�K�6x���ÔQR̶�J��R{_B�;�&b�T~�Z��<���+Q���b�R	�O�9fW����p�Zl�ߕ�N��a��!�;'Iǘ��iCo�!����WBr�t�� G�I�%yG�9}�~9vڵ�SHm0qb�h n��:Q��?���.3�Ä^i(I �[6t'S�̒���ط #���E�:��>�Z��/�5��FW���T�1v犐�}�W�4���{�ש��n���xH�(���o�  ���L�q�Ľ��l]ReJ�YijE�jb{�����;���ԑ��"���H;��p��O@$ �2���j�y����O��C5�����N<���f⹚����;G���
 &��ʺ"��8����z���JyL%i��
� �]y0(�cL�pw�/C��[�g���?���k
�w��ܵc��s����p�ٿb��
�=ba��V�1�"�t:q0�ʇ��R��`b�hҰe����i\?��G��X� �]�Q��7)^��ߡ��T����"�z���Ff����F�Pu�K�2�	��R �"�����.������*�6y�Oe9��L~��lDM�0X�u���<x�u�����[�\/���U�au�c-A�q�� �
%�gFy�	� �Tm����U���.ʤ�ck��b�,�u���^ҵ���G�N[�R�:��nr	���*�<�nY�Oz����x�<"�����������O���" �E#~��yF�D��8.RX-,`�F��X��<�71�6�+�'�p�Hm��rc��4'@sq�2�QP]�����F��6{L��&/���?م8�/h�ȗ�+ê8���ʹ�%���P�,7����$�+݈�9��08|1��mA/m5��������?Zf0�!���%��R!��mٹB%n��6�����sT�S{��UX�ărYe�u�5_A�B�S��y<�_�Օ"������U�'��);�7V����f{�a�C�:J4���#S�e�f?�����`�Տn��V��u���_���L�!��i�$P�x����}�3L�l�������f��|�9$��@�	�S�O�����;B�^2�z�^Q=���5�:��X��,߫˿B��\�l���{���J	f7�i8jX���kh$)IU5�$?�n�����7�'[��-��$��y�R�	�_�_ݳ2�ah�	q��ѫi� �o�B� X5�po��w���Oz���1��v�q
V0�c��G�y�C��:8�U^q�~���P����^�|RK��~�C�_��r�jbRסb{���� ����
(���V��Pj���;�7(���w7����� �!VΞ*x�몏ƅ^��Q�����2m�!���<�%0.�f��i�b�&��Ǜ�o��+sҞ����\c��b�DI�����:CߤF>��.q���q1$�1���j�C��g��&Ew�f����O��G��촘�&��n$�U׿J�������%�w3p�0E���vˣ�=�+d�N��8���S�Ǵ;b��)ZE��+�ϫ�$�	S�´�0-�Oz��7�*��։�=e������Z*�^f��F(k��? 8Z��Q�z�6�O�R^�q���H��?K��m�~�0-��x�B��k0��bw�ri�*�ZzO%�=~��O�B�M�&gz���%|9��,𿾡�3�kanj1��tz���X[.�Zs{A��J����ഏf�&xW���1�i�6_;Rw�,d���s��/'pZgJx>��`;y�b�g�����^��w`�0mWh�@-���l$��ʗN
x�e�t$���YUWX?��S	�!)���� �;�j��8͓�n8�1��-��.�����W�H> �d�(b|�q�G͸s�psXt���YNu�{3��́��L���0P>���=3.=R�#MFQ�/�Y���/H��ƪ��T$��g���X��\���0 ���w~��-  ����5�vZ��4�.P������5�ϼ�n�Ӱݑ���C�`>8�$���H��Ճ�ק����zzs�&�c�z�XnS1$���1;��SU	B$6�hgB���� 1B��E}����z"���i_�A&���C=��X�,`�{�"8,ؠU�/k!f����u��D�!�ݫ'�FU�ɓ��s������-U,y��k�4��2]�H��Ď�dOkք�*NT��e��s����ţ2e9K=D�5��y���?���� ��>� ���o[��5.tB�cQ�&lec�k��~"��BL�bw�E�x�d��J�,���!��l��"tc�rq�1ε�F;ܑ������b��u�XD�{�q����Hb��45cl��=[��o���g�ȶ��A�Ê�yzV�3�,�����C@��E�O�95��R�������ڛ�@�ɟ�y�X���K�% M�$rH�*�;Z���z�$Kp�7ݡ'��?m� �Nϒ�v#�ߓ��	P=�*��R��?VĲ������K���ɰՄ�:_���??�U0H��M��
"�gA�5���VwD��UD�~\���[8p�π���d��ͪg{��Ur���VR��@�c����H�{�C��%&�P�(�/��r���
*m6}�F��У�i?��x#�.�]	��a����n�6z�Dҧf�@�m��{�~�}���^|KŎ�l���?��3*B�*�s�2A�|p&�2�+�w�s�g���XǦ���$�Ԣϥfv�v-T��(sق�����ގ�GS��K�"���ZG`�z�l�$�?a�Ϫ�%Ůk�
�WH�J�^�bq��3�s#)+p��6�A���`�-�<�B��|����/Sc�HO24�;�NOr��i�U��Щ)�P��o�����G�Ѣ?�G��L�b�¿6[ZKA��CC��F �0�.y�Y���n�ۢA�jTm�_��+�[���,�[	Wu�I��u?G10s�voȓ�V~V-��a �_Z�j�*�PZb��Z4g�sw&�6C0gl���+��
�.l/��B�(\⿒C�|B	Ɂ�y=I�!������|A���0�O�2d7B>�S�����)!��Id���z��©�W�1P�e�MeLGU�j6���e>���@��qƖt�V�ڗo�:�5O�Q(?�[��:�L�fD%'��Mϧ���J*�6Q�
�a���AO�c��f�R��
f��F-�iK/�/-�͜1_,R��\�S$J�&��@Q>j��􋃩z�L�P��N�<%���O�}��ya�h���~���͘%�+���_۞)^P�a�<$�2�dKf����.4¸�����1 �v@dhx|W���Pt>?Rܵ%:	(oBm�4�9>'�@� ��E(��xA8��\��,�_-ɭ��LG�rm�4�bf����,v�(�NV��8Y�k�vU��;��j|լ�a�h��rnd�)��,N*��%�̤�����Q6���nlad���0:�3�'B�l!{�.������ �%��=7��z�M�M^r���P{iv�(�cSA�ͬ�R	0�)��O�e#H�!;���0���E��T�­>T��"��]N�gY��44�6���ޡ��{�zi��s�w��"$�kư~��1�~�K�lOK�q��[}�[T^>e�xB�UET�S�,��D�ޟE�KR V&y�~�^�I�BGQ��ì�v>*r��eI�g���E
4��p��m�\'��.�.w͚N(3��v�4l�D�i=�w2m0����J��h����G�؉��gE���fg�m�6G@��w(f���I�/�K���K P�g����=��"�||�ɧ��?	�MA�e2�r�pe��^���̏�͜:.e����EIm' �LY�����)r3曫��N�N��x�K��/.��b��O��5���ᾼ;�z=1�G���'�#ĵ`ဈ�������V%l�0��][�ҜH�Өo��9�6
�D��U� /5	ov'TiArA+��n�S�(d�N����!O-�d���31��K��S����&��G���e�5��g�{5�S��~��2	�iQ��E��:&>��t�]d���s9p5�T����!<�}h�w�>���h�y��!:H��jn����%M�|�0�w�o��U
� |1���+�Y ����=Q�F�Y�.=�-���;�;c����?�n�ܴ�* �79�*��7:d�H�Hγߍ�A�(�a�i��;�۰G<ޢ��	�N����w�c3"�8�X��󬈝d�R:���ܼ�ʺ�`��W�ls%t٧xF"~�(���}��Q�5�5�<��ڛQ�A�p>�dz���������:�f��*a����3*Y*el�Q�C>N^֪b-sn<JNb�}�v�.�39�&`IYh������7������ɫ_S��z�k�c9
Î7�E�X�q{^�Vc8P���~�wV]wa��0��4�۷MB�!&׿d���,nu���� 	���o��vp�-»*�W�k�6��sB��Ȃ2/ޅS* �0ƾ�X�'�x��2��?lD-T�Ц��ќp�K�> /��3�Lg��M����q�B�>��1�3E�y,;ɺ����X����"X�����i=�����新�����ϸU�����8���[�_�H���	Lu�G�qC�f��Ev!�l]�}�c�ͤI0�p��OH#��[C�GH���6�|�p�:�կH�R`����[Z����VW��(&��=�t��v�:����-)
�q �����ҝ&Е&R��ύ>>��cQNh}���p� �s
��۽u�����Y�M��,�Q?�8�S�🀾 �*YKU:3��ќ�?J��Lelޮ�w�ɣɣX$~�<g&��q�.����n��p���ƣ�Gם�Z��� i��_��ݪ���/T1�;���*<�1e�B�h�OCQXΥ��QH}nr#��E:@ѯ�05J�e�߳�::u,�$K��ZՃ�S�z�K�T5����u�0�{��0��vZ7P�RV�\����#�ZQ_M�(�g�	���'Esw�w�tl��E�����"�c��I� u�R#�ӱ*[)�4z��Po��+�5I�(�l�oȿ{�m���ٮ��ĉ�Q����m�T'�爠Y/13hڌ�U#�M�j܋TˍB����Zy!�С��4�n˧y�mx��2��@!#c�)�g�?��,D��;��7-ĎS�򚜋��4�� �R��x�Q�q~��_��r���A�-�r��;_ο}���F�zS� �I����7Q�u�bfv���V�A��s4'v{L�Jm�Lr��!��󮾐6u�B�P����%c��-f������F��p{�q�P��c��-<%��/4��O��Tp�NP�-�c㐴���8�}T,�)(As��L�&pA�M?!�N�z����!�)�G�6���l ʹ�~�O�%>�׬a���~)�s�]�E|�π{ׯm)��0�����i+f�]�����I@PǛ�-�)�A��bZ��j��T6s���+'��uK�h����YH��,<�N�h���Nr���_�CpiQI���\Xt�tN��UsDbTB
Ǉ�%fUc�^y�v��π ������[g:��������"$�p2���^0v��k75#s-b�JU'c\�9���U���|�$����v�m��E��v{F>e����7U�E��^�Rl��1<J��oߡ��wE�J�N�7����!�O>g��Q��V%�i`��e�N���(`�k��9� }2_�,;;�0UO���X�7�o���� �mT��j6��TB�x�s��ُl8	���������ЍC1i�~N���-��ˠpjP~:R�Õzu0�cR#N�h.�)��Y3�=?�!���h��c�"�D:�;�	ڹ�kBq�-�ڭ*����Cdx,l��{RCLy�������v�Ϋ�N~ 뤌#^i����I־(�1�����
��~�cDJ�S���޻X��#�?�$�Z�x]n�`m�9a��ǞT��g=�n,�Z�2n�u8(ʿA��iA}��?*����8'GYl�t]5��q��+uSw�D[ t#��PY�t4�Ѕ.��o�JW��nK�D��yTb��'���6���NV�c�ؤ��^d3t�^�+�qg�qpu����6��H�3)�����I��B�{�E���W��Xa�<&�U���7E�Z+Y���D_w�+��5�G�M��O]���u�9nl�&iPG�t� �p
��h�`�3dy���[���6g�u��8����:����ԢN&0v��5yd׼i҈�]Bԫ�<'�:��NGJ6��f��~4�~x2��f��Tg-���3�y�G�������nذ�HV��U^E�յ��N-�����6�֦�E�u����{�K�\���ޭM���ޣgz6"�u/(oS�<]$H�C2����x��~���FJ�%$�����gZ�3�>j&�*32D�r,���vL�/����A�}� �}��v�.�FQLv��JB��xt3�p+�p\g��>]�5�Fv6w�S��gF�x���IT���KX2aa@���Mw�V�L�%q)���m��:15:���pC�d����'�:F��8��(��bGi��5l�Q:t�0��Ġ�t�3��s-d�V�I=�, �uZ�_�qWRs^�s��)����q�%�rJ�]�o5�8g�R����02G�Şv�;��nGYPv�eٿ_uR�`���m���v�=���7�f���J�g}�ޒ�4��[��|1m��ț��(Y�Νj�ꓮw������K�#T�e嬅�x��/7��)���Z�jǃ��Ѩ��0�����~C�qV�DٍN�����	,����m�E,)M��f�:'�pB��'���n��?�t��@+0k4�Vr�i�:�í�ů�.��jG�d �]�1(�y�F��>��욎=Z�}s�Ӄ@���0H��#u��d�L&TZ�Ի��Tn��|2x3a7�c���*����U!�| 1��e��P����;�~�Z��L�L�q[Zn�~�I�e�R��լx��-���.������6��O��d�y�i�����/��?��I�~|l㘲2W�8�F�F�p���4�^|/Zr$҆���5̜>��9�u��JY�9����f�D)^xZ�C,�+�)�g�W�s�*��R����m<��v
̫� ;�d�b�槫 ��O�Ê�9���"�E�f�'�	��ݯM��Jpp���äB�b>�5;t�п��� ,���\�jGԞ3�s���a����H�`(	ѡ��_��@f��5��o�2���x"Z؎�h��tn�=u<�a�Y���+��Ue�XpJ���0�	�6�/�k����s���)�	='��=�\����ҍ�Dr�%��3K��U���i���!�kj��K��� R�8��x(,�ٲ��"_r�����r�;�W�_�M���@�ă>E�ȟw�~֊��ܼVj,ju�N|0�$=��>̽�J�;�Rl�`�^3nZ�H�an5�jԤo|��1~bB7d#Ư��0I�&)��"KG���3
`��(�]�����~}��U����c=�5����I��ޅ������m�-�D���=�ʦَg�d�<N{+Uv�
����`W�i��ȹ%X�#([�d��*;H�/^Z a֚�|'a������sP��}�y+�BX7� �"o����*��=Iݻ@<"��� ����d9�S%�^`E�W�i�����dJ��;|�WP|��P
�,���1ky%�	JƤ�0�;1;/���1�	�υ����1��b�A���M��^�Եn+��"?��n`�>,GmhYr!f�~�a�)�Ȧ���6�_�eR�y;��IX/B� ��w�Fi��iK'�A��@s�N��%Xw���,.�O��v�� o��J�b��1���=t}}x���Y9K�f��J%�7}�ŮJR����g���\�E��'3��ʃ��%���W��tin+��,�N����4�lzmMZ5�ut��T��#�n!_M� rf�#�ߨy�:�ab�1P�H!��@E��3Yd"v9ǚ(gM+��y�JK`cU�Tӆ<�1"�h�a��Px ">���B/��~W������)*ԟ,�VdCx5`�sw�ys���������$٠�a�B��SRv�Ս��P���qչ���<��}"5g��M�p��ʎݩ�M�b��Toϭ� 5i��N]c�@���:P9��|��c|�@�	�:�����H�^�5Z����#�DkGg7��������` `�#s"���<�z�5(�E�8M��787���K��F	��N�P��� !�m��zy�,��������V��4�!�,)
�������������廑�U�o��`7X��F/o�<����8R��9�Y���c�ad�����k�7���= ���鄴q�<%��$j2>e7�f%����͓��8\m�x�0�e�co@"�9E� mF�"9Kv�9�Qv����#J8(T���!��`��}4Q~�Q�ԗ��G��AB,4<�=����n��G�1��ڕ#��"h�HҶs���F�Z$���K���(:I�~��S�H���ė���l}��(bcv� �?1;��_�5��ܝW����yL���!�j?o�� ��(n⤊�gN���r
�h����ƤY�*��p�<"��PSJ�Q�l������U)2%U1Z� |��<c���m1�*��� �:K6�-�M��!�L��Ib��'	:O����D�4
]!��H]�����aOX&�=�S�Q�nI3��ᑅ+Q��&�fK�y-sզ�l�����M٢�(,k�vrě�d0,'����R>y�����4�왒���H:ȩV4_�Z��_�*G>t4�CXJ�2>C8	����R�f���g/IV���3��\_��CE���z��m6z��Cߩ��ùm���'h�r %Ne��m��/w�+��u'å~*k{2͇](�8x@kl�����X<Up	���>�����_�
;�~��e�sG�4'Z*}u����%?(� m���'�*&�(ς��p�̠M����4��w!Ө�,>��"V�to&@�Z�B����)i���Pn-���������OD��Ff���g���+�j��׾�)C�	�p6�i�˘{�L�GA�gV�:�Y�g�97!��s��ɱ��W:��z���&���W!����|����R>���)1+ (�~5&�|{<TC)P:��Y�3� y�C[���0虹��9w�L���Hy�|?s��ن:L"l@o���F�}vEԼ�RT�h�ءN�8�m������f���6؝�+N��%�R/a�%�_!Jtu�y  ���l�KP勤�E��qFk���c(c.y2^��5of�ʆ�ː��]�i|��b붟sQ�X�ebLr�$c~�`�>R�2�q�����6(��+��vQ�u�eC���rǴ����t����G�՜��U�X�	ʵ�6���c��h��m�k�>��H�9�X���?������Jr6��~	X&x9^1���q��2��E���,����+�";+���3/)O�J�
Kx���G#�i_t��55W�hI_ְz�W0�h��c���u�s���tT���~��
��dOŗC;��)�@�\����O�6r�F@TdS�9��9ĭ 6b��%�9M�H�۹r슷c^�E����+�S�p�׉~��N$ϼ_/� ��ضL�\��wb�e'�C�]�c����C��ytF��v|������SO�Ns�W
,7���l$=.�ɟ���Lк��2��)����M�}Nu㋁oV�9���H���[i��E��h��"��9�Қt���I�p�T�P��r��Q�u�hm�td��;Ā�@��O	�e�l��J�����V�����bj��}��j�huT��W���{ɽ��=˾���s���MH^e���YU< �g�W�(;�%� :�v�Fg�f����$X�E�3߱h�ėA��|����u�1����e�c�|p�\�9�4�h���ȝ��n��4/��(��\�A#�-a䜶�� ]����ÿ0OS���?6�Os�����L9ex-6h����W��d�dfO&�tb���[z.-��A�TP�Y�N(O��������. ����+/:�<jG��/�=!H�$5�����F"0FW������#W�x�f�~�䢮�VP���M�L����Y�ո^���ً���/���y�X�����=h8vy�˓Ɓ���LȲhA�v����p���#SER�_� _u\�s5iiq�.�L9i��*���-��[�2jR�] ^^��&\" ):C ������~Y�V�-{�_��[s+0qZIudQ�
��XV���U�����=)d��,��68�1�3Y.SmY�)N��~��ͪ��}��皴+[A�(���S��/6��2<�އ�d�Cnt��!����oW�n����S���b��4�vڿ@��"�tH%�F�CC�w�Z���r����4f2,�{N�?��8�)K��f��/B�}�ļ��{k/ӝ��.�H��Wh��ω;�8Yi��f i�m(U�z_��h�2mH �o�Ҷ��½�<�^���g��7-��JM�����M���@�Ǉ�}���۱{
���<[���n�? d*�GVz���>��-tY��J~���~�=��@o�����v�����Ib�B��9t�-���>y��mѧ�`�q�skÄ���Ƶ׷D� 1�y>�����dg��Z~��b{�
ñ$�:?~���T��A�y{$����.dhh*�۝�^:=�v��	a�<����pS#�Q�)���v(�{b��(�H.�����b����_�D�g�(�e�r��ٓ�y5�!�s��<�����b>��#�����t��`�Z���WeY^��p���'(��/f��@t�3����e��U�X=�|˿ㄾ`�g����ret�#HW|�PјG��e}Z�T�
x|�z�����JX���;1������m�a��b�HCMN�{�O"�������)�><��-A z�*�`�m�5 �Om�34%�NF��{`�DmPlg�d���T���#�O���׏J���<Cn6Nb>��t��BA0M�f�b4S��a��x�,��qL!��x���P�����]O\�*L�A��<���x�A�ʍe�G�%,�iVW-[@�e��7�
��������{��M��D2dj�o�A8����kpK^MY@:XP�i���k�\w�f�ʣ�2�rF٧(��!vh�ش�]��v�b`28���xv�P�)�Lj�N�_����ڈo/[Q'���,��]��`*^ ������uE���䑫%�\_�[�5��PPP�����31��Y��K0[+�<���X9/KI�L2��|��_�%JH�S�n��ʭN��_�������%,�˞V�`	a00�Ƕg���Lr�i��y� u����g<�s��O� �-��'A�c�#ꔇfZ��.;k�J)v�Eg�b<c���Bl�x��<�
�i���-u[pn�� ޱ�B.=��܉%l�pu���xs.2�n��⪸T�A���dZ��O����8��]
�,0�z�ͤ�U���h����X�}��	t�sSƨX-��8�)w��/v��~�7�p� #�Nt���4;=g�I/Hz�gv Jw縁�2$L_�K08Ȭv�f��6�YL1��5��'�=ݤ�Vw_���+��U��o�I,<W|��v� ��3��
����a��=��2>5p,�#��H�B�ƈ�k�T��?7�k�!D;5���1q.�Q��C+-��*��V�;) �o�9����y��1Z���2���
Y�II���]u�l�U����@���o�"�LJД�rM`#̐�X<��,����r�������%���g(ٵIr�g6� zTK��y�<������$�2�!yN�嗕|�r��ڋAP��9���Jx�LC�7/y�b&7���W�ҝ�á
_B�>���0@z���ͷ^�
��gժ� ��)Ppfѹ��q��U��Ք���:i{^	�� ��_�b�ߤ�7/C~��u�ۼ0	wIt�լ����0�7��6��]/~��cb�$>���av�i�E�����5P�7�	vܫp��4����gq����д �:2�SȬ�|�^.W�R4���%/Q��t��z�q��7;h�P�Y_&�P0d{���_<r5��ҎՅ������oE�Ō5)����8Z��"�}ԧ�Y��"�tK �M4���[z�}>�۬b����zZv���|�����E�d:_�ބ����'H�Ֆ�C}��ө�9b���=z_��&�m�h��_c&9���<p�)�����֋mE|"������P&�4�-�"�5����/����b������q�����.w�H����F�?��0v�h	���]�/_����K��Qx�
-�IK ຸfkgp�8��Y��sM4����Ĝ���wZF��UHw�<�n�� �3��{5a�dĬ� ȐeL�@����O͚`06u]����{� �̏�@���*L9��9�Z9�%�����+u���$�r�9���{X<z�it�aϝ�S�UKCbXYJ5J�1q(�hZYIe?1K�X�$=+����_��Dc�bT��~~$��=|���7�@��J��o �'�=�b�_����,���í�>+'}����������*!��"�p��ݹ�O�X0=MR;Y�<7:�9�e���;�a�۱ɨ@z��1;��mr�j�9�v�̍s|N�A*#���%�����mh����E#�#)U�s#�Ѓ����8��|�}]F��-��G�`j��s|C��B驧�ٻ��)I�C�IO�8g�d�](5��3<���&��V2�l86���g�טF�l�1I��������1�Vs���_p�Ա	lӊn�[0��˷�|k=��g���	�@&H�s=U<����*p93���U<6�b'?zY҉�L���`�|����u�L�3�8��g�
rO�ZB�j�$�IT6#�b,�+��?�TrDt�S�ڸPA�}��� T��.�C���?��1v$�WC���G�=�i���Den� �i[�/)aV���Z�Fһ�'�r��nٕEK���GkTW��yO�gB��ST�oH��[�rs�c��2��>k�J�o��_A�Z�aP��˙#T�DXF%�/�B���f�\�I�1fv���h�B�M,��&���Q}pž9k����w$�}������joVM�>y���-�0N���M�<�jQ%��-�tP�`R�tP���l�;����:1ؾ�#Z$>~�o���:�ěA��y۰Nk�bﱖ �jc�b1cG^}}�A8��p=��;{�=��X+�mW��A��OApx����u��O��a��q��J��`� wxQBk�*�d.�A�ɲ(�օ��1dQ��1�Z���?&&�Y�K�k)|�UR�� w(��x�:��Yg��4�	ܽJ���DYlZS�#isR��|0 d�P���^$�M,@���T䆹X8lٙ+�	brD�m�+{�qG��&?Ga<�v��2t��ݸ�u�O;�8UI�!�F*�����q��ل:|�:����+��mH��-qx�+����+@��}�~}�S�Ă��PS��:a�{Yb?�tA"�h�Aq�2�i��0����'�Z�	���Yk��Ѷi6u�C�a�n�/���u:���Bk����q�9(�u�������+�a5���8e{���kb\�Y���v>��qwm7�Ԝ�x�=�n�,��lZcI�}-D#~QiFP��U-���m��4���p�b�u�y��
cy����޺AwQ�����ր��7��N�pGN�Лm�l?��|n��mMB��ï�L�#!��dQ�!jB�l`��� .�֯��~[Q�l&�K��O$����rF��S�q��fM��Ӕ�5�X�&:@����,x'C��P�"ـ�k8	���o�)W,���
�����'7wD/�\X�>�i��2�bY��A�Ζ<�u<�}
��"^2&��u�j��r�q��Y�1�=.)=