��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
���ۇ��������)��T�'�L�3*�51?+"�W������7���׷� Y�[�}nP=�PyW'���J14��qKxW�୽�V����+)Ό���-�o(��Q��`�`߱��H=%]�ȗj�u)9P��?L\�Y��rq�+W�||ꅡ]����Ҿje' �3��V�K��4���M
j�t�҆Pd�{�u�{d?������կA9�O��[�&�o��ʯ��j����Ǽ��Y;`�=���7B� M Ry��X��[�/�����f�E\
�`#��qK �T�PM_�?����w�/����S��Q}'�dS��&tZ�l�ϵ 5g���q�}�-ft���]�..pх)2}��d����[sH��;��D����џ ���AWBP�PJY؛U����6�?U	�	�0 ���_K"����_��m��T
wy������AAG��ӯ��`�t��"�r͢u/�4��wj�l|�>�h��㉏��c��#�8�g�{ۇi:��?
�P:
�ك��f$�F����@��P/�DH��;�f#@�LjaFO�`E��{ �]��N}o!��M�m[�~s�"��s�p��o��*#�q@��(��_r�����h�R�҄hb�U��+�7��p��ɚ���xWs�O$�r��G�$Mϩ�P1N���	k��Lb��V��y��Y@�

���͌��sa"��`&�X]!�'a������0Zepr��3���U$QJ��{�Ѯ��Z��a\F'l�;��?2��Y���l��c�.�2|�>�o [\��*#2WSe�W,��_��7l��u� �'z�<� "��.��sn��{��O�����^�2>( ����3�#�Sp����5�q��JpgQKi!�F/��̠��lл�-� ��]���6�օř*2kS��h�o��$�����p���Y,��>D�S��mJ�5�d��탮��ë�n" �M����]�j�Lk,�=�ȏ
��?Q��У���3��I��K���7��c���c�%,C��(L���yɶx�$P&���Y��k+�3_!k@��	�LK�Ӏ7��إ7�f�N��w|�!�T��9w�[�`g���e-j���⚡R&<pF V7tZ����w�c�ei��T>�D�U�I].�0��6�%�4���y?��(^ލlu�[����� #O�+H��{+�-aL�d[,>Y���:��S�-c9϶`�J�rjYoL�8�5q
;�G��bўf����7���Y��I�Y��7�ɰ��V]�I96BlZ2��E�]tQ�풉���� 
UAL)���G��Y�U%-b�4>O�d0+��Ta�-�3M��(�m\@�lco�TV�E;m~����'Q�������+
���P�W�������s�*;܇q���i��U���4�=z+��f���o �YO�^�\�g|�_Bi��(�� .�9Jy�S�=h cU�����Mw�7D��������A(�N��h��l_W�X4jm�ǔ&S(-7G�&�Z��tg���q��*�οR���q���a�jv~7e)�R�q	�\s��o�|=���@�Y��jЩ���hS��6�pG�N�*8v������<Ɩ�U�:|=I�g*%�1��X1��b���{�7L�aX}�z@��<�t��&�r痧h}��E9�<3�ۆ���?��`sn2��M8���qqNm�l��������&��mŐ'O���}��ĬCfd��uOhX�-
 ����;yJ{1�6�Z���	�?Bm�o
���Xx�&�<��yl����Ghb��Q�R�z߿�	�ҢßyV�ʰ����Bg�l���a���rڿ;��(����l+Z�q%1���'�WY��5��n����+��B��Uy��㒖�Y��H�՞eK�̔�U���/ B��
���}:%*��l��0�
�+m.L��Q�;-�zJ��em%�;�]��HC3		���U�@C��J{ޕ캋�@�k�ߤ��[�uߪ.tG�~�Io>!�t}�O��� 9I��c^�F��b���-�哏�,����p!C(T�\y�A��l0�������@p��/C�-��(�i�_4PW��c|�����	�|.�a| � ~�o��U	I]1��k�����J����p��I�P�{+G)(�)7k=��Mht��y��f��w
��yL@�o��1���ͳ0n�b��n	J�%:�3��U? '�ө�;O��bF�}�����V�.K�T�����S��RRߊO�]�R�C�Q�	��`�K JH�*���@o�U�gV����sUi�9A���&��,��9�]�)g���~�A�D��!�7W�����J&�@W&��L~����&?��H�z&�Qέd���D>�<�?�'��_�;����k��(�8���I$���3Ͷ�a'��0�u���W�|�g#*���a�m�N�맡�|�DMmR��<��K�=D�Sג/�s�	�KO_Do�_Ց�N�(�-ś��"&&X���F�k���l���An�?��3h<	��WZ@�WUm�3~r!���!_�T0�d,t:E�
Oi�µ%R��O<j~�����BЗ�ήNW	���D'��1[3K���R$��5�~�	�rY��&גG9��~��Y�4�{I{��`��3N2^ ��_�%z���Q*̃���h��g�5j,]|h��`a�sg�����W;�p�X[v�}$�����xoj:������+�3�8^�-�/��D��� _/T��i,�.����0ˆb����G8_π��"�N >�g����G�<��M,y���z�g�]^P��k�)�%���j?����%�%��aBOR# ���?>�pT̕ ��G����8�ʈI휄�����(j]��d~;y+�y��m<��_���� %�� L_��<^^.i��S�xS�Vwz�5{���t�eR�Qw��C���H;�����w^�c0"�� �Ȇ��c��7�zG��"���ү��^�9[{J��J�׈�V�3��W���j���u�"⟕�����"|{�AGW��EOL����#
fup��I�*+3�����E��W��T�ƮkK`z0=Ӷɫ�xM��h����>�ATAH2�q���o|�n��J|�'�G�v����4�����_��Gy�>�@�q�����"�j@�u�*�%�ҹ-Tuo"^��X���[�c�ۦI{,ڪ�Q�0 �Ĳ�}ey|~�5WW�q���x'�[�!8S`ˎLA�A�p$=�K�E.ya��r�'��R]ߎ���M�$0�rt�(�=���r���J��oD�@Xt�
2:��W���}NC�e��u��+[��*��7�yR�Yq���c�XT˭��
E�{jാV��/
�NZ&�&�{'q��L�Ó�3�ͭ�ŋY�41���{Ȕ��"�j:�����}�����_f
�5h�{�=�$JU՜ٔ�G� �k֩ضU���agT���MW�� �l�֏ى����½K޾~�πKe3_����eL�d�mR��wA�wM���C`���m@m�6F<@>��oD�Mj��yJK����7X��h���h��ւ�xC��Ϗ~x�)����;�
RQ��Ѭ���͏N,���s�E�����7+bW"{)c����+�z5�i� 6QJ�]�p��~��h�k1��?�rea��Z
���(1�9�N�)″1W���@�]`���oH�:��N�bY��}�ĸ��*�7�Y=9ۉE���j^�U���0����sݔcA�I�X���/E0�E�|���LY���������F^_����c��p�<����n��v�TC�T`A��t�	������4}|�$����>��֦���+tPam�,��m~���ރ�� ��geH��<L�?r�&dXa�DL�{aa��Hd=G�׊�5^���k��+�!�/iB����֥�U`#Rʊ�6l񂢰i�oηtPr���@��[.�c��/|��!��N} 1�}hŔף�Nݞ��_�.eԨ�Pb=��k��U�oJ^��ڕ$ͧ��r��V�:~� �hpð�j(բ#0�����:�c��ft�ȝq��oܬ�, ���0���3<�O;�塌������+��f@�<�yw���rC̧.5-�ɖ�)I*.O�mj\�A�Z<��O��Ǘ�%Ǚ�ڬ��|p?b -- �{�&�2ѽ,�X����)�^�nTb}Dv��ļ���I9��BAng��Q��Z�7Tl�8��ķ=��i��;���t_غ1*����y��N����#b�䓒���W�%+�`�J:=m���m��L/HbCx��V��Z~����+;1��@�+�x��L��?���G��{\�j�kK�+.d��P��|7U��.����q`n���ϲx��A^jx�.����8C-z�ǯ5�{�CS����}e<���ms�ϒ@�o�o1ۤ����L��������)�w���3�#��0_���"}ߠ@���u����R�y@�k9;��y�,�K��7^�-!���c%X�����m� .�RYs���$`8�Pp����Sѧ&-�� �L�4LC5�һ�yA�O��Y|υY�&�����,&$�vk4�4[[�jԗE5�H`�;�G���
'(�T�J���HPiM�=���\���7�M�+X��B���6�IP\��/7�F�� 8����l@�fB`
5�rO�"9k�2��$��D���6���D��?��lyQ"	6U��Rsw�����s�5��/t2���odE���ˌw]	GS���9^
�����
x��L2r�,���g�L<@���Oԉ�NT�l��'
�ј�U��L��_#��HgL̯�^��z�2�������¡�L��K"��hB�^��U�(uɳ�lO���aѦ����'�^��uqVf��x��xS���y�*�{�v.�!�%	~��m��� �CY���h��<�������gJ5t�֝�J��N�t�����Վ�es�'�}J��ſz��U��A;�;G�ļҫ�5�k5=��oC� �;��a��HJ7��d�0U)s��o�'��Cx�����{ѧ�l���$Y�����b�����f5GX�tG�*��ด�b��it�1dO�N��I_��Y�EUʒk2��u1:�{����RN5T����9���Qe>$ZO�
�P o�1şx�t�1��������\!�I�b�x��@gF8t:�*��1�Y��Z�Yz�%b�D�/`�J�/~�o(vx��b�X����+ae�@�e;zȭ����F���%Dv^a/�ȸ���#kV�p���������d@Ga<o��!jm�t�n����>���F43�a=�G�������}�3�eP�*L�I-���*}����Å)�ko%*��
8�ϒ��=��6����>L6�s�͉cN-@O��EW�'R���#��Ϋ ���YY!q;�s�#ڰpq��cK.J'p��IG%���NqUG'��)m�У¹܇�`�X��nm���\�y� ��V\KJl]|���qp��jR1��p�-֌h`�#T��~.���iPw��e5ِ���(!J.�:@h��"�q�x'��_�}x5Õ̍縅��(C�QX�dx	��zY���3Ӗ�'��w� �����yY���|��ۜ瘿�3�\(�VGO Xd{�k
F�~�)�a����WeT$��p󽪳4�U��t| �K�'�V�U%Z��O�����+��HW��I�u�3 [Ê(�q�쵍���a�4MK�4�h�,��LbEc�ζ&�Y^E���'u}�(
���Nk,�C�Yvr7Y{�/e��[�o�sF�(W�x��l�l)�Q`7FVF��{�7��V�Yҽ�[	�4� �〗���uSHi<���7���hb��Lx7��ǻ�8�#�%�����J�%�_!�����#�(-$�E'��0�uy�=I5�*����3���J����Cў&3�z=ط^c�J]�t����L'�ѧ�Ѩ��h�䯿_U���Z+�_X���F�4%U�J����� ���9���H�꼶������H�����s>R�
��8�$#�5�6E,�\�"�����"��-�z5�\W��n�ϗZ'Ÿ(�t����b;C�N[TSe��"�kU?G
��G�vXAa���j`H������w��5
���F�"��M�?2pJ�S����b�ξ�S<�%�q���S䶁���|*��vQ���-�͞���(i¶�o��*]����h��ձ/��I�ˋ �`�ԥ]�'xU�dJ���]!/�>�B�awfz����V�A������5�8�v,p�Ml/�em�1�ڤ��K�/A�ݖ��#�r�J2����.)֐�Qlx�i��i恵rD�%�$pGS���/�C��6ZT�&�Ķ�O$)����^(��q����]���Q���tۮ��uXa��?u��������
q�C��ښ��̕��ba�V �2#�)|c[��ſ(7%B��'��=r�(�P����gR"j*�����k*K	/\��q����sI�z�!�i��3D��Q[��p�@Q��;��A"h�I+/�S��u����>����PV��YOh��Y��'a�Zi�^�����۵�=��/�8 �(��r4�jp-���F�yyn��EƐ���Xy��nP��?���)y�I��W26ȱ�i��^3��qj���pk���'QㇴBr�u�~��m� ��0K��
5��������0R�D��ix�~nH�{�J��?�T�^�J��w�+�S��en��|Ė�[/��i�cC4J�
�Y�j����W� ����e�.���@5�����1�ݯ��xt,Q3��ܤ�1u��� �0���p����s*�_"uE�	Еr�K#��p��I!��#Ɇ"�L�=ۭ��'�����sW#`Ȁ��ysYc�փJ �"�yk�A��.�����]-�K��QMg��������S��D�@&)]�EcA� �#��0B�����'_�v���}����ڥ���!B���"�2���S��	�w#�]AԝE�zOx��[�rlɠ|�q�����4�{���}@㛞����27oȋ)�{u�#u��V��g�v������T�XR7C5���~�24¤���귃��>|���;�ʪ@�mv�h*�J���j`���mt>T,H0����ϭ���pǠv��B%&?����'���B��K�8�P���R��f�Z�m�����!ߖ�;�&�l�$����D7�n���d��!�>SEeΤ�/R�WmLb�-��|Z���=�yA�R��UW��Q��#�So�� �l���ߧ��S��:���U�͢�h��⼣��l��
��j|N�X`����mz�j<jV����W����*xy�����DM5��������߃U&@I[|���"'���PЯ�f!���q��3�n�o{������9 �_h%e9�	r��a�|  �82>����<�$z�q|��v�VZ����'M���P?��g�܊�Ġi�%7cD�c�����?Ġ�,�y��,|������ʁV�Nա���G Py���psf�_eɍ����h�T�D����`��o��q���Rc��{��`e/�a�hQ�h���SfS�u�bC^n��]�BU�'|{�z+sE �n�$J�(�ns�r}z�ܰ�u���@���N�MtINt���M-�ȫ�B�j%�oAa��w����>_ jGw4���
�z��5��J��v1(��/N��JD�ִ���)$�~�����0��Q�+��r�|+A��$N�9�����r�.����t�n��B�CM2�'�n/|����l;-^���l��5\���cw�bq4*�x%f���h�ǾjX���N͗��/����e�<O��6m?��%1ϖΝ	���~!Ӝ퓍h�J��37�/�����]2�U���ۀ7��@S��Gʁ�~Y�m�X4$�R=Ç{��4����8z+u��oM �ڻ�&��-
9�q��Wp��5�n�㚰i�4P�5��+l"���of4T��Fe��_�o�����/qx&\U҃/���S�e8C�Z9è�����P�(aL4טĚ��
�	J3��FFV�S�p�}W�m�e�;ݸ�gA�S��1��A=�$
(�0�t���ѐ��ċ�֮��>43��Pҵ�ηr�Ԥ��Q��v3�k��Tt٥2��ڷ���otS臃HC哢��*����XlǤ쉭c�k9�����7��t��	��0�|�.��Q����
��:���iD3;��_�;W�{�0Ǉ?o���PKf�y�*}j_�>��	e�(r�#m��Vs���qa�Z7���|6���ϵ1;�҄_$N2^�WX��T5E!<-MG�9�R��0%j��Ư�=����p�d��H_.�Y��.xPS���b�,h�g���r�;C�3��U�emElTX�&v3 4pdN�S�K���A� Z�^��KLU�qL�{��������VP���O����M�f��P��w�K$�_���)�勞�����ʁ>7�Jֽ�m�Ӆk����6l��蠭Pc�/T���t�=�/X��R��!���5�i8.Ţ�}(�YƇ�F�!\��Eh]� U� =�\�"ȅ�3��� ��>��!�l�㼫a�is!ׄ�������o�Lץ�H�;�tAm�1�s�f��wI����Q�_$,uoڜ�	��{snPm�@2azQR��UW'Gފ�������+px��Ch�=��]����9?R��x��r�|0���wK��5�)�G}ҖSg	�d��\��Gr�2�1��lӾܾ�P��~����k�^zj�œ[�Sy�L�'
LHdc$諠>���z-����l��Y~�V�5w:hA�i1s��/��~�/,����4��@��v9��/��e/X���`�� >��7�d]4��.�ǧ�CV�5ޗ���o�O���*rD��
�ִ%D���Zd�MѬ����\ճ�����.;yڨ`f�<(u����{�S��q[�I;��>;��vC\�͟�#i�p�N�(�`�����gR��h���9�d>%ر���^W�ȼ�c�J%��擎OEAq�����*�f�צ9d�]�B�ΏcX۝*��p��h��������'w)mo�Ht�}M�h�n�M���y���9�0v�^6+:YvjHk�Z����/6�􌏊.���á��*[�8ڷK��64,���p#{H�~	�S��$�U�v�u���.��V����&`f�<@h���"����y�����>��'!���D��lU���P��y����mvڿ�
W�0�dˡ��i�q^@s6���Nߡ����DU��9} ���Z������X�F�mhy��-�V�H��&|[����(�fy���y��`Y��&{�ɰn3���� \���]��$�")eL�!��r��؝Rt�d{A��R�]~�@�X���3���
��4H�I���F����1�]��\��KS��ǫ����6n�/���%Y{B���כw{r��A����-}�<���TJ��/l�9��5�UI��u�7-���>�����cMh�����bt�/�#8�;.�M*��&�{px�#KO���.���m��*��S������p���'1B�S�d�$f�=���t�����Ĝ��NS�I�Y�w�P�����R�]n��ai40u��Ĥ-��*�v��>+�)���w@�J��Ú��굩��H�M����)\ �.ȴ�hWV�.v��)Cڜ�Q]o%�����y�w;@xd��n���?V
9MT�B���Dq��	�D��`�h�	��/5��������0. �H�a$/������0q�SDi��r?�&9h������a�D�by�l�9D�
���0�����调��8!rg����lMA�W�?1�#�
�bo�*f��u��n�q�5�J���<������h�{�L,�dZWe2��X�t?&�1|�")o�A���S��:�����s��ޡ�6d
�
T��] r����g��a3J��K�c�A���Ԭ$��5�q����<��$�YꠤTalM+�Hw$���/�mS5��d�5�]�H��{�7�D��4�M���h��=�|TɥG:Y�"���~�40�h2@��:3!�n��g<KS�#��xZJa�[�m�dK躐K��S�|Ń?�k<i(�����jAt�z��Ҍx
���"����P7�c�"�Ss�dAɝ�XZ�$�ȭ
d�r�xR�lB�Ĵd���$c`V_'D]�[ΞCk���q^@G�!*�`�'�/�e'�>��jk(�RP��`NF�%��]�;c���bXE�C0��߳���<�ן�ǐ3�HD�`X�_�ٮ:{�*\��yd�����H~�7Y�n�����ھ�O��2�sP{�I���}��G����tU���2K$,m�x!��x ��s��P�[r]�*�<�.�M�����O!���f^�Xͫ���L�L�%n��++nr��