��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�L��58b�Y��u���ۭ�E �i�s�D�9#3]w	�B��(�Fͤ`a'z����1��n��n��oD�DHU?K�N�<�].�K�3��d}�a`F ����.5aE�?jR�(��_�;�4�`P�VG$溒���UK��1;�+)��w'I�Ҩm�THO0��|h@#��P��!�*<'I�i� 	{JZ:��Aw���]WLж���ͽy�d.&���&��-B\��Ni2A׹I�������z�`�I݀��xu��<x����q�tC����6�"�e����\��I�/�g��8�n�r�,�Vog�0���������9Ld�/<�V�Z'�uX��r���M7���i�@���6�ݑ�׸�5T,���.:��#� ���):Qc�c�w&*��/P���샞��U	��U:/�.��gx���d���*̭�U���w7��.O��]"����ˣ�;��֯���ٿx�Dݴ4%�_ZtS	�O�8�%�v�_���iɫˌ9f���15A�G��BS����.���pA��i���LYM��u���з�?���*�J�;*���7���8b���j8|��D	��~<�i),��3��r��Sz�e��N��W\�I��&�=����ۀ����?Ҕx�:��څ�76Ԃ����p�䣘9[�Z��"k�;q�ք]H�������Y
?�y�HҧW9�u"��k�pN�ƨ��DB�ˑ���f
Tm\Ǘ5a��(#>�-i���٠�� �- �r��ϱ�=kT��u5*T�΍�I=(���i�����5PO�2p �R��e�#�1�TYʄ;��j�7?��D�} �O�|�}�;*XF�������5O�e��_X���Ǯm�'���W�ra�6&z't���2I���$6cw�@�pc|׸7@"{�Ժr������#�n :�o���|�V^���Uq�|�ዄb�/~�FX`Q�N���\��1�"㴅��K�~q�7��K��ͬ�j��Rf�'�>HǮ���-��e��䋃�o�zd�;�A�qW\�r0��xƬE����qn��J4k>�u�஌�\r��O�w�n�1�r����*���%��g����G�l���#�Nl+|[u���s����it|���v��y�r6��]�>�;��V��]������_���U0/h�� �1t�k_�S�rfђ}38yx	��9VI��s��}���o�!����5����7�t�n���3+�8I#��kC $?���y��H]r�8���2��]�������P<O�3!�R���_,Jk+�?x;9XN�i"�,�o$����<!oߑ�`��g�B�}4�F�|.rul��0����ӃR���z
A�~WH��s���SR+�ų9�*5�e���u���T����sN�JR>~D�o�6�_[���U�/�ѢO)Č���z��ݱ�	cn��7X���a����J�/���V'dZ��vE>���*��M���-�p�03���HN;Ϧ� �$��,�����-�+0)uX�����:n||Z8�E��3�zdo��rgQe�ξOk�<�`�W2�����K�C'dF�����f��u��Vg~�yx�@w~�1X���]�����`��?�:��*�
P`8���\A���E�^�`]�8���6�cM��UZz�����a��c5�$i�DL`;�	6��:@X�$`-���hw��70�/\ޙ��^�̚���rb���6��;�rK
(��"i�B�/՞�:��
5��d�괤Շo�U��S��.[��7?κб�*�ev��=�m���o�4�n����}3U��}#l�\O��"���6R�ӽ�!�?s*�٤<ChM���0ڏ �B`BY��Q58FU^�6sl!5i�^�)u�v�"�*b r4R����Z�!q*��?�k���H2�?����G*����iَrv�0��L���I����W�(UTǇ�Ue|�襞�Zk�C\�}27�?e6	�dJ��!�������<]ؗۀ;�TQ{�E��)���$5�kW��c3b0��f��R�Q���솓����޼c��ڊ0si%�h�d%c
é4l`8����@#�%
�L��|3\�a^��*����@n��j�����8=��	k�]��KY5y��H�p�Ol�og� ��10��X7�M[�f ��L�&R	�Fsq/��r�a�z#\��j���g��oϴ }p����z���S�K��j(� }��r�"���ƽl��
����ʰ��ؿ7{��I;N���& �h]p,X���+Ҷ(^,��PiΘųHS�!8qՀH�Ģ�.@�ۨ����>�^m���9Z�)��N�X��X�[@�P�1��Pb��a����ҷm�p��#����Eԙ !�#r�l_L�(�M�p�F�7����<O�ܦ̴��U贐{�*��j��H_�Xh���i���2��	y�4����(�x��rX>�/>p�#{��Ϧ*i	�~�soJЛ���{=�B!�"���б����`�'����#1���cy�p����=��|�Z
��~C�-����^Q��d7U�(�z>um�n�+ibi�7y�V��ix�N`XE��>��fLhPqAabbG������R�IH,�0Z	��p���=��cqD-�NC[=ӡ�Q�-s� ��s?۞�� 'N�=��DD-(��..�wLe|XRQ7��?\+y'���.�Ɍ�~�'��6~|]���xYU�tR�K(�U�z�S��䲿�TV���Uի���dW�#�KLnۚ��-������Ч�n���	��d$T�iZ��K ��&J��=ciu��QId����3�������SjЪS���2!+A�3�C�=7���m,C%����q]!퍼��Lf����(h;�0ok��x��;�3`���m,��p.�3z�zLD���X��3���ī:��F;�W鲒��.�&qP(�]r�y��ۖ��o{WB*3�F���v��[Y�6��;H#�m�\f��Kg�t�Ĝ
I�GJ�HP7֕��"���8��*Z�����T���*�\�7��PXm-����mr�#Ž}$89���ϧ����{�߰.i̤����nH��4�<�Q0g� �ޯ���|�j>`�Z����oC��
���0�d�ZU�K�`�V����s�b��� |�`�T�P]z��*�:�5��C5��3�#}G�F;�\@��ۙI�չxI��tK_.�0q��]E���-�.�;�5	f�A���򣑤�5������F ��&*�@X�Xx�Dnd�V�yA|oݳ@��W~6��kp�	[0]��S%�E5�g��'���l>	�A$�02�SESǉ�*��!^$Y?]��U���O���3