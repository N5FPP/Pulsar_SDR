��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*���D#����=�6�c�p�GCE�N��+�xh�Eaa�Ƭ�z�5>��>s(�oƤx]C��F�i�TϚo�2���E���W�۠N	Rw��#fa�E����ǁ'�iM�$r����?�W���aݒ�3��L��'�ފ�q��p��FU����vJ�k�~���l���wFpe [�29��Zq���)Rq�� �CPu�)�;��/�V�2��'cu�*�Q��펊(�Ľ�|�3ڟk}wX��r\�� ,��E��:�Wг��P��t��4��o�=9h2إC���W(jſ�ns�\�K,���~������}�7�p�T|@���v�����f�P��R�ތ�t���� �ܥ����i�e���Nm�LZo�?\P(��?�Fg�V�%�.��d��NۗຢyˇLG����>�l�.���/�#��
T>�&�0�N7�m�&%X���:�G���¥P����A�z^�O)r��X�B%Kƺ�/�2�oK�6�W=��^�9��e\%�
��,Þ��#�a����mt5��۫����/���I��J93ض+��3�� �|WV������,���:�޲S���m(i)QV`S���o-����@�es_%.��Čɤ���Dǥ[I<^%�ya�%�2�^����[X�vJ
tJ�l��H��+e8�lB_ڨ_��طΨ��Q�(L6�]~�y��B��a�y��苈4B���Xl3W8���|_�|Fg�"���h`����w��P���fk�+�s!��0��FlDq��9�#�T�KK�vs��/zc�A��\*����+�E�����w������w���ω�XO�ٿ�c��h�e�6���J�$9`R	�ѓy=�a҄���9�["���v潕�Z����~�,�0X; jT��C3!�>:���$�Э�f(��.��1��X������L2̎Ȟ�S�k�I\܀�b>�u˸���Ds�E�[~3�Eu�0 &����_�20�3h֦֗��O�똯(�����In�Wjϱ���od���럦Vv]��D
L�@�Ē�LfJ�
��|.=:l�m�9[��)�y��i�`[��Y��DY>�Pp�c޾�MC"���IPU��<!4œ��Dn��C�#Q�	Sa�%am�|@}
��Q�CS�8J�ʇ�-��p�F��+1[d��_��̄��NK�l9Ep|��ۋŐP�>BD@��&?��qm�(荵�`<�5h-����~ �O}"s��rӶw�4�f�cB�zRQ���u��6��2�X�n��o��C%�R�B�`���/�,<�)u$!럩��ލU�ɷP���6�7
� \��FQd�	��A,E	�G��y����9/:�:J�H�"�UeSI�,̋�k?�K'J��L«|k�_Z�����9k�vY�3��:��/��X���*<�bQ���q*�x<	�Aˎ������ư)��o{Vv?��L܂�ˆiiP���BI�I�߱>
ԩ�i�����*����_Kݢn�i�6^:�5d��2b>�`����.:de�W��$>,����l-3~�Yݦ����*��;�z`± $6a��W�
%2����i�{V�[����h^��V��&�L+�ѓ{=hX���`·�t��K7�[�3�J]-�Ǡ'J�·0Qy
�&���Y����&�J0)�>U�H�T�wa�YҞc�U��������&X/��6:�����8�Yɯ�:����������{�t1 ]n��-i
�]�ݮG�i&b�xbW
Uj����7(�W����>$$[��[�m�nT��%�5�Dd�������@<���̈O��kb޺j~ߦ�O<>H5��f��8�Y�j��V̚��)�ZP�xj����8�d�
n�����r�K�{_8��v��}y]����4M)�m-��"�����HP�.��+��Y%���|���k���]-���[��U۴.R����?����`�p���G�|/�d)Ȯ�ݜ��0�\=���e�}\ު���BC�N�u�t�nU;���c0L�˒�)T,��yǉ?��P��g(�>E��II����Mˆ{���c�S0�/��P��;@��,b�1��3?�(���?�d:�v$��������cU��è4߾������E�@R��3_���%�#]@�i�L7V4�+x.�7Ќp�A&��%��]d�-$wov�P\�%���2��K��#(V
R4�H�I��0�k�G�!hknU	�5ꉜ�h�du���M����$$
$�2�0h��: jF?��������n*X�)�;b��s!��%a�[ePi�I��S^{�?;
�%^KkY6p�ʢ������eFfEӈ�θ�!ʁ�8j�Ѹ�Ƈ��[}���K	�#mR�zh�Fwz.�^�I�L>+�����X����7؎�������;���E�f�<���W[���$��[��|=�2�v!�c������8	
J�<�d���x�G��趶��,�=~z��}�K@�d-45�R�E�rӻ����V�|�Z�)䏎����s�α�$�v��d�� �(s���7�B��d��;�P1`��q��W�l8�z���\&3#r�3,�'�h�H�%	ߐ�;*U_��C��*�%�4!-ݳy� ���?H�B��V��.��	f���;`���3�b r`G��>�X�hך��2@�K&��j"7Q���t��xP�߂��L��F�$�!<���I��[����7�nrwTRo�D�k��:�r9fJc�W�5�<�[ǣ�03J|%J|L�\T�u�fe�*G��N�<�������A����$e����>�|�*fg��b�J?���*:�m��ym'&)?0jӥzͯ��a$(��ˋ�w�lqa뜜3�����L�b3n���
U����sX�>�?�Oqa�Gy|�3�0���[��MQ�vpn��
�$6���3#�_}�|oW�]=q;��rݏ'4�'چ������>�FK�G�Z�п���!X����>����YYF�N���0�q�&��"�kE7&�"H��)�Uf����w�b��׬�,��Y��Yf܄���.D�ߔUM�~��A+��Q���wΑl�,��,;��>�̵`a�8�ʘ���>�;h,�9ǁko:�?"��e]�']���AQ1�#���g���[�)v�84�H��F�2uK��"����(�vg�^]�Bg��C�A������y�B:�Q�3���t
���&mAG�?�s�H]n^U��;�E<5��P6i��'J�dC�%�vх�v�s碬&�%
����m{�DSh�e4�8&P�I*_��+S��\�Fz��\�Wq���i�2t��q$�6�:��&��Oo��k��������Ҝ��c�3�0����j5L}F���Q���"CO�)6�nU��5�FW��	>�^1��ת��ht�x)x'���:�X�����1D��/|]+��^;�g���@���2����Q�4�ny`���ro��*��c:D�E2큋���v/E03���祺xl��TbI`H�I����?��j�.�V{v������m�<�����A�fJ��%��'�[�3&B#
u��\=�k`F���Ǖ��s��.TN��CP{��&�b�9 �G����Rk.�B~��ܛ�@Ƿ,�`#)qb󥶈�t�+�� ���9�_mv�u ���a���yf�.�9^�TIF�\�l>��2��[�ɥ��)�gnfm����*��0`���`��lݱjrs2��
I'Ri`G�@h���,����.�C�ɗ�U���]��:���Q&`Sya�Y��/�DGd�0ʡ@�1�5ﲢa���vb�8�$��:��%�5Ѧ(Ⱥ��#����d�Dh nsVqQ}a �L�����887��¼ʢ	����
@��L��?Y�j�ֺ6�٬�m��8�;�mޯH`0D�`�R眊<C�0p�����Jp�#ktC� ���"���=��7H-��+�Эfu�6�B9	�8/rG0S��)�j�{e���R;������Y��a�x���v�nC;�[a]&쟸���k|��\�:�xs�����2iTV ����*��Fڱ�+��$	�z�+P���P����y��/���p�uV@J#@d��G4�	3=X��K�����^�J���}GP�����_�O�Nf��O��V:Ob��r�Rf?!}��d�¹����� �O�y��/��!XD�[�{X�y����bK��e���57��
U�>V&�\ɹ�&��, ,z��5����S��ܐ�r�H�J`8�)Ë�650�b�
�lC��ɴ��O|��pѦZWH�`!����B������r̟�L�C�Ȋ#�8����͸G�J��D�{��GY@в�{d>�{8=-|J%3��J�d��/Fa�m	ݢ驅�M�G����~��� �tH~������݆Y��y���R�J0F@���uqe����$�cɖQ�@�Ł��w�	��k��7����n�3�)9"�T��#J�Ê�_�k��T��y0�A��e��@5��k�$���4�M���]$�	���8��ʶ�<4��)��|W��g%��']��]�m��1ɺ@��6����[�%�C�y��\ٿ��[�Vଉ�k�+2��#�"�Bya{e���(Y��[��"	�bu+��(͑ê�ϲ�+ �W�)8z���`2!�h��rZ�	���_�_}w6��؄�l �ы��B_��ѭ��_��81y����}\��&�H�i�}�Z,��:��%Op�t-�J�3 ������뮱��2ß���¬�j�ݵ��U"��O�����l?7��V6�l	�� ;����Q��r���A�s�'��Q��-fnШ��*���o�_�/?��8h�.E�1�7�� ��<�$9N����(슍�B
� a�Z�>���w�^j��D��~2?5\��t�|7֖1b{+�ћ��m@���|	�P�e�	�xS�hi����X9~�)q�S�A�8S2F	ݧڳ�-%��^����&B,`3�Z7n�H�����fl���V��wT�f�\��
+@�a�/��ˇv�aT���2����>u��v�Ș�HIV?\	53���od��ٿd]�˲����3�l�l5�><�h�W���7R֪���?J,�	kr=�"߃@	���\)z[N�%�y�8�^�	���
fS83���VK-��������P�f��	^#G�w�3��o�a�b����V9����+��R1~w��	��؜��:u[��Tc�!�.s��w6k��l�R��/��L(I�]4^�Q�JD߃��a��N��L��Q������������|%�8 Z��*�(y)V��<���؀���ԻM� ��Fj�Ic[_!)D�"U�<�Ó�-�;�}�s/0W�4&�]*��)�f�H�V�&G8J�o�U�������v,��ny���Ik��ѵFQ<tS���+)�IM�M{����s��fWXؼ�B��{aL[@��hԏ]Q$V`ͺ.��D�ُ����f-e�c��v>�ڽn�f��ݠ���kW�oEE'����BA"��(�0�v:q�d�N�4�5Qu�͊k��ś��=2�S�X�nTf��n/�%��5�߫�Y�h*=����qFQ;!y��h'j.��ʞ�4��Z;G���R
�����v��o<�#�k���Oa60�&��hv��*Ka�Gah8L��.K͔���m��V�u {x=�qsR6[�&�ioaRh��3���C,,���s�e�x�����6�8�������t`vT�9�S$�oі�	�';4��� �$�FJ���8�A������x�J``�I@�Nڿ�=��[�X���SCCf�^1����{�'���
M�� $�2��~t{8M��?�f��Be6������3� ���!��jU�<��XH���{�l�N1���*k�L,��]#*m�P�w:[�-
haE)#8��z*�ֲU�V�u!s�f����Mm)/� nB5 $?�ꡑ|3km4�Emd,�6t�99�";���hbs�>~�{�%���1��Ǵ�:�ŏT�{�0缈A�v#	�n�A0��9/\���I���'�(DA�|I%ɑ�6@׵lv��8q��]�(A7ޝb��S���\T���s` j.U����0�D��z�vw�jotW5��6��̉��(�lج�Cg���ϗ��O]V����?��կ�'����e\���Z�������㗪�F������X�&��H�&���f >i��{
`��`�<_���ۃ����q6��E%�&�T�\ͪ���$<��=S�����4�:Ջ<��P�aO���\��(T2��M�$߾Y�����Ҋ��''+��i�&Ɓʷ��D7f'�����	D��.L~#�rL���9|� �B��$�X�q��@e��8v!s�"m[�s�A<cӡy�]��Dė@B0�X7��,��Dn�y��O&$&�o3Zh���dIb��l�8��
�I�H-oVנsX3WWL�?�@�S[��]�n���Ӧ�cXqs$[�% �2f�*���[��aS�-}�Z�ܔ�ܰ\�K�p�'�mqTi3U�¢�y�.�ixyO?�LH����p-��h#���Zxf��/�I�:�2Vr����Cu8�|�����s�����r�~���e2�h��"}�JB�םh�����z���R�?�C���,ê[��K��q-�֣��-X�p�_��	���$Q����S"�8�闡��Z�P��Ö]��k�_�lF2 ��[Y�G ?� �Ǒ8u*#X�:���&��:�4i&!i�2�a;"3-c��Z��Ӗ�_xW� s�2��-�1W�,��u���!;�6�n<j�^"�S���
�����>=-��X��4ʍX��g�|��z7�����- ��#��uNt����[m��9YȞy��~����Q>?���;H�*ŪF�9E^j�+���ia>���5r���CvTA�0�=�W)�3[˼��KK�Ӯ�V��V�*�ǐ/pg��gH����Oe�E1⭻\&h�Y6:w�HX��p� �7��
��E|{\�}�H��[F��|���j��./|����k�� <ad��^��}��m��Y���|"A��W����(r
��=f���b6�Y�	5��4�0�w8P�'��Se	xҫ[)�?)���t%j����74e�29�FU�&��='��2S�����Q��������[��e�3k5���(��vڊ��e��Q�!��n��V9���w�_��b)��	͘@��aI;w%`�EQ�aU��D�_;s���Ӿ�QU
pZ1���&s��¡���vPlN���iH,���E{c���X�j�V�)X��I~,�����E���	�
AD�C�th���N�`�eX�Rd�/�i_��Rf	1;$��S�̓#����]�#�^W��g]U��9ϊ�7k��-�#����bרF�$6֕+���p���Ӌ�Rw��"����^�ד)̎��b������ω$.��w`3���O]��xɭC"�E;��܁�@��p�;�����Ƚ4�[�L�pbQw��C�����aPr�q�r/���k+��c�[�Y�C�;��Ҍ��5���A���U�����;�"�	|��bJ��"Y���l:t�bz_�镴��ȝ��5#�D���l�:���K[�p���ӽ3�����B�<�����+�Z^�S'd6�"�Gl;6!�ğ*9��ר������A��+�8������*��w�_�(�;&�A�f$�������^^7e�Z"8n��E��*�^�G9����:̻�]̆3۾�k�������4v�����b���v7gC��O����|AN�q��l�\���[���|�0R;�@k8F��w��PM�W�%��%O~��