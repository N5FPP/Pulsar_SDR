��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��e�ik3�������w$����g|��J^]ؑ��4�����[!�?�,X��E����|�r���N���u�g5�'@mn�s�S	�]65
��3�Pkd��5ϼ������˼*e��~��QZq��1�*[~|�y��pP�'�����6�r��J�\�s_i�c:fDSj+��H��5�2̛�C�����k�.K��fhn��)�$�C9s��Dq�ӵ����yU��?�[�s���9��ʋ�� 8~Z���#sÓ-$���$��ߙ'm|�z�,�ѕ,�}����v�p��-�Irc@��(�8^��X�F�x�l.Ӧ�K��$2�-Y�������t���|�;!�T��s���B�N� �RX���098�K���m#�c�C9*��u���h��U�6���;�v�m�*1=Y�p7�C�"6=���4
��"@��i�+#�4z��b>&HGsSߩ���E����UjaZ��ci���b^�F��M��y�Q��������N��<���#�f��r�5ĐG�"���Q��7������D�:+?���'tO��l����W?�j�/��14da�4U�\&�Fڕ���'����aT�x�� +G%r�����T��ۨI#Ox�Y��/��ǯ[Qi�zD�G��}��g�H1��Ɠ`��%�-
&�����<����砐)�S����*('�x��h�/��a���x���X9��L�v����Fg�rq�(�ڐ���?�1�g#�������������b4S}`�4ZD�禷'�X����)=����V`)������#����ͦ�T�ڹ�+�<�V_k�}�:�Ȍ^ �B�pR ��_}$�bӉ"@���
�8�$���UC,6��]�&(]�|���1)��6g�䯴@�0#��wy�G=�jl]��YobP,DB�>����hG��2�a�)#c�������g�*����g`��B��b���^�(��v�|�s��b��S# ɄMV�0o�{}�thI	�BcQG�7�m0�r�a$�O=L�U�/�ƴb�zPH���t=l��0���kO���:Y�d�>�<���-�{�L�Fx5�4����ͼ��G��$���=GU�ͧ�W���չw�ͯjk>��j�T�QP/wX1�z=����w_����Ra���4o�tuczZ���2գ$����|g�/�� b03)���	���8��-�+o��E�����t�"�~oʯ�cɥ����6�g��h��E��̑�η���\�^k��r�c�
]�ޝD&]��\��k����v�6�h��H��'L�ߺ^t+�:�(�j;� Dy�/p��V���nk�INH��m7�ߑ��Z�Ld����ZKx�|��>u�ߣ����{Í���!6<��ezS�A<���l����EX��*��	�lI,�|u|��I�5��	�]��pH�2����M:��c�[��f��-�MU����)}�D���pm�hYSPb�=��:���W�$�d���H_*��ا�)G�~��2s�;iU��:m��U�3����{%�A/���"��vQ�Uo��|WHԶ������
W�p��u�����'���X�t�'�<��J�8�N¨w �N-�>Z%��DԺ���J����P�ٵE0N�Xo�|k:6���4w�����x���������|6��:A�����ڧa_(I�so����м��4����%%��õ�]���"J�e!�2Zf�ܣ�p0^��A�����r��Ad�٭1�D�>��G��*������m�|��8خ�p���͒��c�0�~�<�n��f�)��Ao��`�J���~�3�Whv�v���SţZ����^��!S�:K�js�du�OC��$P���Y���[�G�����ewB��e�p*T����̺}�K���5�*G���}�$x �S�X�����W{e��Tm{���1����ƫ���3�B'NG^���5��Ԫ�<�,2��(�P�w'�����������˪������[�8u�Í{9�y����wT�lE�Q�$��-��B۹n~��1&�>�%�@ѧvJ'�C�FS���Γ����F�D���!BQ����,/sֻ�eЛ���JNq@5�?�j��I�J�*c�ĝ4�#v��?����_�x,�K#��p��,}���Y�;Ӱ%���V�Alc=��<��p���ڜ�AO���I�%�ɗ�h�|�� �儊v޳���<�AD�7�a>Hy��F�Hc�bmM���.4�Ǖ��X�e@���mxׯ� ��yÿ���ŘLf>)���+�yk�39{�pGeѼ�\�+Q���N��)c��9n"�;�L� 9��a��%.j7��-�+G5��u������C���񩡕�ϯ}t�̿zb�1���al�:D�ƝQL
�&������L�.c�6���#D��?�x��"$���`��|�fW"��/aT����>�g�����4�WBâz����
������ux���}������4�g��+����l���ȿ,���QDLg�E�a�E�i .^t���n��B����D�J*+ީ)�P�=Ğy~V�F??��|�D�0�yJ���F[���c< f\n�W��m�]���c,����t��N�i4H2���0;��9S�b�Qu��u\��� �j����#<����$��Ĝ���3jZ-�\O-�U�%^[$�4���ެ,��(_�
�������m4c�r������I�{]�>����^ ���
���Ed�������ɣ���'�aϐĜ�K�+��v���j�.A���"�^شH|�-f�H3>hN����	��:��Fm�[�²�}[�En8�,%�O�3JX�g�t4����g"�E�P�g���+�;�'.�<���[�Jp��$枍!+��`���� �+�| ��tfv��{g��� "�my���ʡ�f�Zaό�Y�[x2?�UK�#�s��������8h�Չ��]�SM"�1�`Ē��D�D_�y�����P�>�i�:#�G�r��AdPK��w|Eaؔp��z�ٚ2���ŧ��3�Q��QZȅ�׫T�P�R�t���09�*W�e����rb��
#�����8��;�-cJ��".85m�o:� ���s�]SHƘ`^��@,��L]��FJ��m�&'Wy�O�d'W���D1����ϵ� L�'�I�W3�Z �C"��.�5����y.��Izݝ�I�;.z��nG8GߌM�E��%�>�(��� ��ԣ�
���J�.75Jm����*!N�KL��:�������W�p椀)�C�z�g��}�(�b���X&p�6�U.2�hS��(�J: (0ֿ�d�`�ƣ-�\,5�}ޗL�Fgc����(��l��*1�� k�}rϊ����H\!�Ϧ��~���u�,�b���AXfH):5�Y�����o�&�Ib�o>��1Cro'V����z��!]��mWബxA{���������0@�XR���Ɍ�V���n�h��5ٞu���zQ�G�¦б��3��1�Ht�e�s��X��~�x�U�w�z�y� �C'�����v��&oَqrY�Чɩ��a��	���}"Y��o+�;�Ę����,���D�'uGЋ+
� �����OtS�['&`�ɬm��4աDg����3zȮu�@%m�c��@I%�>�\O��D�
���n�!�4�C���MA���KN�0�6�Шe��WU8�Ԇ���ŷe&�j2L�k��w�/�j�^�=���_���m��kPT�P�M�H;�6?��	��zq;�n�����]H�j�LF�.�����m��zc�A�������nf���	����W�z �N:�}큑�ض��D���� �ۈ<�F��^�s&��#�u��1^�	�6��` ս"S���"Sԫމ� n�߽�F�~�{��F�Zl���x����$ǫ�:�m`؏�����zTsظ��W(͘��VG�H��@E�k���Ǿ��[�r{{dU��"�s׭�:�G��rȈBE]��i���;�&�
ub��1Fe?,�7�7�h�΋A��K�:T�;j���4��Bÿ��jTp�=b$�	��+Ty�o�
W\��'~���J)P��w'�k���O;�ε���	��c����7�R	�6�cq.�	sihN�[��*�8�nqc�I��<��OH0`��ֽ[Pa0��w3�MK�!D�۟��=u�p��Xqr�s�,�L���{�+���c��EP�G����U{���+DmE�c����ƿB*�d��<�x�oU9:�Xo�gYq����%�LR��ڈr�9��Z�+!+<��X� �	�@Ɖ_�P����K�ı�m+����
�6@���O_5�ep,-��|����E2(�9�K10{���Pf]�K���U�Ln�r�������������pƍ�+x��-�e�A7�9��=���a�0]�1g��1�1;{�� �-�%a�}g��aC�u ����v&�����'ͱŇ�&Y6��6�=Zkf�����
���7S�^���l��P���~ǟ����kI�C�C��tڹa�i~���Ta8	��z��������qi:iMOO��XJ�u�n7Ŭs�8��]`�o�b1���gT��	�����f�Bе������|ce3q=���ul 9jo��rF�zA�M�&g����= 	�|��s��q�����:���!#,�T�{��\�Y��Y�l*���p,@0g ��$�t�m�fw���ƽx�9rp	d��~��"�mG.R�J��`����r�׈S9�,M�7,���[������YS��g�ulJe�^g�͹?:߈I��|��D�*�G|���	��h:���y�cİ�����C~M�P���/�s ��^�����襛���A E�Cw��� T�O�o?���$�>��5�S�:]��]������%�ѱF�#� ��p��\_�;Įǖu�^\])R�耤����o��dk����u@�7$ʖ-"��Ԫ��)+-����n�����p4�`j����j�U>Q6u�h
�%�v���.�
�:��ĉ�?��H��o�X�;�-)j��$��ƛЇS\I_�ݒ�\���'����y�I��6�1�����	�[�뫦�����8��I0QU
'��P���M�ՐdF�'�ң��|��D/���oM)jG._�w�_Y��O�U;��s%ʊ�g\K���$t�=�?��j�_SK&sÿsx`��f�$�� s�u�,�3�C�F�����!H������D����c�R]J V�`T� �P��,*�a��JO����{gs�I�0�W�+B���T��_^�q���m��8D&���OY<Azv0���<)��p�����l8b� �sP4:(��rΨ��I��%����J�K*kn��J���"-�v������-��%������|p�b(����?�3����<kxp��k��wa�_	N�Wu�.G#Bwe}����C��H�b��O�k[\�S��6V?x�"m��_�'����&�/!*O0� ���2p)��&AbFh	N��ew(��k]5%ZwBZ'��@l�R��ὒŊD�p(��R��ipSg�^��D�^#8�撵k�aA��=�eQ
�y;rOX)��>� F�^����7p���)L>+�Y����#����>�u��圫��jim��j�Mj�j�:.��'�h6�ȉ��n���kdj��պi����ȎEU��OѬ67w>�Q^�7���O���s����3,D q�"�p�J��#����.�U�������C��ǅ�����i,w�#� }΄��D���i5Jd����9A�X�����x��c���D��������0�Q�UA�F���@�-	 �=���A�dC�Zi_ ���Z�+��86���#T�5\tM��i�7���%^�0.h������0�JX�;�Î�l
j.���������J��<R$�[O�n+۳�ؖp�0)=k�+ma�~�Xd���c������ďwe2B�,7�.����	����|�#�25B�XbH^�\���Gm[�u�]m�e��E�E�m�a�o~Ҩ��͋�B5i�pv�g�T�ot� �$��,�Ƨ��mIstW�	�x���yt �Ӑ	0>��%W���L�PvOn��A����վ�M���2}�_8a�;���N���*i{����,�: �+�߇����U�Y6��z\�VR���P�^$tF�֤<�7!127�-�lPɠ���������qDp�&�T�V��"BD��^wJ����ͧ*�&v��U��3��8a���	��?.�U�4��3N�7��UߣX)����+%a��p�~K��Qt^�U�/��e��Rt%�^e�w4٫A��#��L+e'U�C�x|��l��5�	w�Y���"���r����j�ZQ��~�4��Wߤ�՟"��{��U�r!U�j�OS�2�	��r_ihT���@��	~��&�;���X����B�V�@�\�l/I�>��!`*�F"�Z�@d\�Ig���p��\�ꂇ����0�m߅�:�5���5��D����@C޳�.C��)q$n��K�n�������i�狱y�-�7�v"�M*f\����3�h�1��4siU��P�)f���טDu���9������d��L��$&B��V����?�=D�'m�6+I��}���� �#�g.ߺ����B�E����bˁ��� K �hg�&���M"�2�����d_� e}[4�af�/u8�f�%'EI��Y�?+n[H���*�Q9�N�:��_��ץe1�[�����7|��zA�3�^����I2p�F�}��qp��/�^Z"#����	��D1?�`|��~���/��r�,٢�!:`f�*�f�t.� ���:�E���U�IW��`j�������
����������ӑ	�鴌U�ܠ�8�trs@�8�ʏ�b^|����i��+�b������360(?�N��ʮ���9�u5u�߮ݦq�R'a{�_#�(_@ȷ�I�B��>o#��Pϩ�
+`�[B7g��AT7�X_òg�l\0,�:�z��^�T'2VD������8oS����W|�@ѥ#��%)5��O9D� �%(��[�hD,}��H�%��{$�%���6JS0��Z��(�z���a�S���u�����	O�~�+،
���V� ��Kq1�,���D����b�CE�Ζ�6h��荲Q�ތ�(7�Z�]仉v���zg�1O�n�=Z�;�>$��g�J�W��ɂF8���]� �2B$�s4�煰����2���՜��Ǡ� �ҳ���p[TPȝ~T�r�p��G�M-J�B� mr�a2�>��	�b�������Z�]�D�WgW�Rl��FF6��$�5e���x�A�JN1@�Ի�����v���n,�jz ߇����¥.��>��&C�����@�*��>�o[�>ƃ�}>2��P��!�`��w%��ρ�J�X",�C�0ed=�X�Z���GUd�����a+�r��'�9!
���e��*D�?�N�j�b�/�eD��9�X��.�a&��g���[:��)�61Ϡpp�}xj�Ib��za������yyl�d(�L^�`�����/�Ess:�Xh��'M��`c�LB���*$�5��BC����f��.��Z�w�^�=]��]!F�udW��)}�m�SS:�8 ��&^YB�@���<�	1(�LI��i�3�/�|���%�K��gr�⊟kx�d/ɾ�{���=P���lm�R�¬�⋾�a����=r�l4��%��u>\�W\a}ܔ)v_��vf����i|O{6;��)��|8����|�Ո#m���3\l�F��UPYJ����/���]�ݢ8��[7R��dM>�8�x*ҩ��5�ګu&�l����u'�k�$��~]\��A�=��]1h�oac������!h�&����-�f�,c\p+݋�v���$� <�̯iI� ����:�B�8แ��q<f¯HD~Z/�Q�}G�n{�5i�C�j	��a�Xc�l+��)���}{t� ��QΜV{j����]B� �=�q%R�	��"=�(v�WQ�Q��r:l��u�i|)C����.�LD��N��\���%�O��+e�g�-�\E{��i8w}e#�Y�:�������iM/��j�b�-(����v�,B�}$u��b�2��>oh�S�m�3��`���K��7�u8ע�w�X�*^aW���P:��߶�>���绚�\��y�������y��o����o�����Q&�C_��Z��2h蒊�5y	�a�˿5M��64�>nNͭ�bS2��	���+�'�F�4�7&H@���l�q[e>������E���=
��I��ՇK���.�o��ܺ~E]���|� [���o�8�S�����	]/�¥v���1�����=��} �r����;"J4Wjvx��e!�>R��ǌ:o�X{K��&4�v+\�����v��|��WG�bR�m ��f�,
&�/Y,�#��6�i�y�s���R���w>�p!֜�ű��"ȱ��Uh�յok���S�Ș�9	��b ��T����`�L�ȫkE_�V�d�z�(���C�!va[@J�!��g�U����@�\K�[���ѝ�8�E?s=1~yD���w�k	j����̪fA?�i�&8�6.���=�%,�^��
f��bE�>RXB���2_�d��G��p��/���M��w�y	\ !)>i��imm��k���di.c3�>�.	�s�7dsT��ŕ��XM{��������� :�0����U��׶�a���P�����
������������X�Nڟ#�N�q�{�p9������^�Pw ym�o��0A,�����V�� �B|�C�ߡ0��H�&oT2�O梞�5����B; �������p����]�L�����?ی�%	�@������ m��<ILkw��>�I���5%��8��K�3 1Cت�d��&����Ȓ��gI;ڈ�*5��L�i�@��&_��W��$���F6�����AH!��������	���)�-Rǅn�+���J-0���;��究e�nr��OI��7�|��a$�kZ�ae'�W4˅Ra���h�F'o�*�
 �j��x�kT!?o�b8?�lsa��[6��v]�ڃ���L<y���cӐ/j�ړ7�6[Zn����ǇN��9ȃ@/9�i�pV���i�H�4"K�sP���_9�碭L�ɒ�/�� ��w�����������j���l�{g��jF��{���p�����}KK�
R�~,���Ƣ��B�%[&A�k� ֱ�i���LNd�O7�Hk-j~0!���[��W�3��w�
 7b��[���y�9z��3rst��w���+Ȥ�эɯf�6"�oJ&醬����1���';�]�Ƀ����i^�zԄ��%��!`I=O�t��U��t���_`�`�q�!K��1�q�
��CsѲ�KM��M4��D���R�ni�p��\��G� β�}����V��:\�{ڶH���Z��C���A�e`\��:Q�i��/�:j��
h�_ꦔ�*]�B��A��X|_-*�Ȓ3hbD��S�B+�6���0@�a���H�Z���)�-�Y/&?��D���[R�\q�2��x�H��=,�k��n��w*��� ���h� ��@G�/�����UH��B!]�jKsm��d���tu��[�=��*��̙u����ފ�("�y/�,����@c�Y��~�s��Pi���2�z�8D��|-������3�(.�0F��,������^�����։t�I��ʦ� #��6b����j�^!��������B�i�B��'D�R|m����@�l��1I��M�N�S��&��I�=�9��u�����?�%"-X^�S��7W���fb3�,�H#Zւ^�F֌2y3|����*������ʔg�����k��XyĐve"�������ā��Q�����p.ëJO!gX�@c\fE�����<:x,<�\̝+�䔬H���<�>�Xb�S�W�80~�R.*ћ���8"�?/�L���?lR��:��$���Q�}8U�_�����੤�(s'v���\"���U]{���(\$b m��4��䂁I�?��k|r&V�VT��Ci�QI��Feiʷ*�(�BR�*���75=2����QY曦ӊ�<}JO�������b��*5D/�L�O(���i�}tܡ���`�׬��a{�}g,���ȔI�uf��#W~֊Pg�ָa�n�B�k�2[5]x�!}.�b�W��N(�N�ڑq�����4XRwdGy\�eP��I��@�mx��-���Z�}���L�����O�� _6�g���7'�8o+Z�y#ثMS/�62[.kb1ga�x�^`�Y��~�w��������������=��a�4�&���8��<�q�л��ٓ[6+e̮����ν)Iiۧ�'���$5�Va;��F�ԐGg�f�n�)G�z�&͚��_�H��Vza,t�C�e��ʔ&��q��=��cI��e�V����a�u#	xމ�+�6�	���9ģ���^��T߽��}��D���P�_��*�#

eiac��.�]��#��d ϤlYx�	{��h��.��5>��>��o
�kW�s}�#����a.��~o/�#��5eіr kS�x,�s�ZԾ�A�$�<��W^r�����ړi�x ("��H>�%�'��-��'h��jD{���w�B(�<�d����/Πg������oVQ#Ǝ��,�?��([$.�5��qP��7�@Bz3��tw�^ޮb>���m����=-�B�C�δ�k��R"���+^f�Nd<7Pz/=[���u+����E#�6�t�ц>���rM枉W���I�<�m��Ʌ�W�ro&{��P]	��� ������fϋlaCwk` {�\A0ՙEA���  o�A�a�'�ו3l��3�jOK��8*��y�QTVb�C�i�����&�F6�A���}��Z�{��a����Բj�A�mn vɼ�����C�7�b5R�[UX��W�����g��.���sY9���G��.@�>A���\��o����鿐,ޮU�σw��o}��8%��;�bJԱ�,0= �X�S��c�-�f�H�i1f�~nI��܂�چ�!����xэ���>���RЋ��y�U���	 $	�+�Ɛ+"��P��<��
�3ݓ��̀�w��#����<s'3Lm��>(����ڧ�-�(�� j;J��tC2�X@�	�)U����x�XtC�h����ބ#Jut�:ӛ����Z��,"0"� +���?,��������,�x�f�A��� ����]קګh��XP�h�<�q���F����*A����iY��D<�2�U�Ȏ�����B�����s����4cߝ<��s6e��$:�eRu��ѽ��j�!}�^�(���xP���yo+��,'d	�ݭ;Ǳ�z�� pN����~�&����q ��b����0_��ג�[�a�3��C�3�]<�99r�w3��H��t��l�-�
 >se��y�^O��陮����υ�>g����n�1/�+�G <��d��3�tĿE׻-_N�"k}�^��_j~�"_��@���r��M4��z���ף�X�4�D�/��f��ԗ�7v[1��d�HBs���Q;; ���j�xJ4�UϦ�>�2���U8��nკPP��8�uy��$��� ��n��]�m|�b�p��G�I_��&�M�c��U&��	zOᥩ5�/r[����E�>�3��l*����]��QSܧa�����0��e�y$��r�:>4b�Ԍ����-�p_��2�
����cz�̱���uX�짚��A�Pg�04��uo��<|�mg-�	N��F!��� ��#�l����n���M�����&abO�5�<p�%�q,˕��TR�▝5�?���6�`��tJ�ݰntE;�l�G0��B�@�|�w��x�`��V;ȃ�`�f����9Nv(��Q��'K,�>�p���&��b���h���#�1e���qW,�i���MZ�y�!d�+�����
bB_I��S�l ��xu= g���K�8�h�C;�)�����sL}_�Zv@8CTM�ꔻ;v������������u����w�Ʊ������M�3!�:0�k�P `�/d�K�W=M��bi�z��91�Vׯ��zN���� �w� )v�+�G8=Yb�Sv�S|�ٻU�-�G(Zc�ڮ�ߜ*3���i��@�P��\��_���?�yg�x/�1>�7ԑ�[�(8 �c\�i@6�.�7\���^ Q��.ŷO��2䰼f�+�b��{���樸�i�0�L�F n�7��t�8�t������og��Tc�<O%k"i�?6M��exO�h�>�`-A�s\�)S�;T�n�[IE7���>l��/���]�:5��TV`�����7��������Ԑ�R7�o�*�s�����&eg�D��7�7f(����FH�B$D���F�좎��#K?_]p0�~$gPGO$��0�I�N㷐Yq��k�w*r���^�	ʆ��C�:)�@cl��*��Yp�f�*�4�����!����=�/E���Y]xs���<��r��&;���-Ƹ�GV-8n���^�I cMBf�R�ʧ�I�3b���X��O+7'�����	*0V.f�41k���������$x&>jTí�^����)��k�q����?��ܜ�B�����3;�dqNBj�|dS�_�"�\�1���D�9�L'F��(PL�U �Q��O�=Hǩ=P��YαXnAU�Z���C�g,g3ng��F
+eg�8�h�������hz�1VHJC n��<����t~|F2�sPX�����:���X@����)�歨)�C��Ƕ^�z�@8݆��v�O��=s��)��O9PK��bn��?#�ع-������}�K4���I�����E��it�g�GhtB)2�1�����Qʃڶ+��w:J1��?���mW�uC�¥�w�Ĭ��o���Ŝ�`�vt�~�#+��(��!WI��	��@�>@,�S��-Tmh�hJ�2)�����������'��n	�kXy�L�q���dt�x3Br/u_F�ڬ޻�N���Fu�6��>4�M��_M�X��c )P�����٨����R�ȿ {T^�Մ#���!�P/���C��?�'6<�+�I��$k�WxoC�??v�����"R6�%�&/l���%�tkN�+�M�q��޽���U�嘑�V�`�v ْ��:���l��62��%&M�rp�7�t�4��y�؁)�|���%o����1=@��n�;��G9h���"���F����g���ϯ$\.7�bg$>D�ܖ�u�y��b�[�ZY�4,��;4Ჩ0MӢ�j����B�룿������l%�ӻSJIj�Ě((�E z	ޑU�[~���:M��o��MNA�ޢ=�_q�`S\>=��:�K��ez4�;\	5zUˣz�����ܡ������{=#ޯ��y[�2���̃n/p\ۨ<H��w� U��������F2Q�4b���e��IwN�Q���:�	��У��-��yp8��R��92���̍�GW�X� aA�y_a�m��i�e�������&Idw����J5�mm�%��Ns���9��?'i�(��|,O�h��6�����x����d���]0'�����V(a���@�Ң����G�ib���]B�G�m�@x��{h�������@�=�lF J�.����cu̿�3	����i�Lߘ*H��*�F���z
2 &ql��eɗ��U�$����tXdܓ���wb��A �^z�9�n�2C�'�̌��ߔ5v�d�#-�/ΆQSʽR5���Aw�?x�ܲ]Z7��a�-�Q��V��z��e���T6'Q�\����:�Hc����3N~�(�!U�wy���:���#��\OLB��Xv�J%����=�)l�0�)9Q�͉W�8�C[�<�I0m��Ja5��0�R�;��_ۀ��j��/�6�(p�S˝�ݪٜ9�=}J�h�x�C8�>G� �A�^����DՁox��+x�Y���s¤���8x�Q�*�2�ה�ٲd�%�`�d˷%��"��?���酨e��<��%ۆ�6�{�X��8H3M��=5�R���%6����(��.h����<m�����a���n�3���d�<r	�8d�H�g(a]�ov������Q��˓V^06��w;�����盓$O����AXw�IE��^2W�K4�[�����ӇI���y�︈�Qz�5��1ϺY���@:Ė�qY�B�@?�T�&P�!\	�j���G�
Pg���8��"l�\��CW�ˎ�2��*��ԫ�eR�ė��F)���F���P6R�;pj�fr1����H�͌�?=�K`ZG���di�]I8�b:��gߥ�8��@�_1�7�>�x~�j�|�A�T�cp�ց�(s�`�z�o�Q�S�K�i�����[�t���L&��m�tQ{����f��'O�g�ݞ��p�Σ�*,Z��Z~[��/j���θk̸"A�zJ���Q���W�"3l�M+�C��r#q/��K5���R%%�݊]�|n8�dt�mW5�<�!d�^g���� �,�k7.�����B��Ϯwa�Ho(�i��D���U�t	��=so�Ð0�!��[�~��=[��*�d�)�/
�>n��SM.�7�|�HivsXk��j5��#�I�i�n�!�vV4����n��W�+|�0��i򖝘/k}]�:!�T]���m�f�K:���}�Z���dS���O��i�{~��G�Ze��V��[7e�4֊�F��
oH�e�~��&����3�U���_�x�슎��Π�?�W���gp_�-�Un��ڐ���m�쩐�xT9�j��D��-z(�\�93(.8�+G�8>�&�A#5
���ƪ1�Eh��L�L�(�j���UH��-Ӊ�]�!Q��H��yOW��Č+'[b���Hk?���w!L}?��m�nX�({�'�饭���<v%��5�U��`7/!����&\a����qI�ª�k�����C���Ȗ���-�88�5��ڄ�jJG1؈ �����I��>d�}g Hù��z�ʤ��T����
;��!���Ö��&K��]��[Y�$��=�i@vL�V��:���D�Yn����S%Ս��<i8�5���·*t�S�3�˱��W�l��z�|7��ٮ}��Ȓ�Ĥ�Q?wH�ω�f�8�FvO�+c��q����O��S`�Q'��3�a��f����\��E��'��������R5B3J���=��8O�@�/伥�B�P�Ɩ�����-G�8�3�<K��?�,�s��ݏyy.ES� ./�(���N`(�W�b�#c�WS;�i��/�.��
�2�G !i����F>Ӻ�ߥ���D'+����?	�;�(m-8�����]��W+�$�R#�G1���v`tQzK���� ��J�0�O����m_������� ��?x�Z7Tu@_�b�Q`*��VFR����k��)��]\Q ��p=��4_�掟�Xd��W)��<�D��������-��9���C��]����3�����s�|��y-ԟ�r���T�*�s׸�ay�g��)�Y2�et:�}UY�+����%��#�AѨa��
d[Ҡ���T.Y1�5��r�3� 9�Mf���e�p�G#Z	!������̩�#���K�b���fdXuv��2Jl^�S�6�͒uG|!D|fP������$���s���_��I����\�6SOM�2+�"���B�③���JLL"��n!ֹ��忲S��4
�����Rma~��n&N-jF�+�8(3!*�q���_�!Y��)����]
�F,�W�#�K��
l(dGi�~Ê����ʺ/�hX�,�>�W]��)���+�@��R����]�8�,����~	=(�������A�j�]p��FW��ʘ�0]^�>���:��8�$�ղ��R}�԰���-pd��	����OS9����H��V�e�j���8�-&x�W�W.=A(���"�՝�2��萪�#�?�K%Ʋ �G ݤ�a�A�m�^?z���n"}~r>4ݙ[���9�:�s΀�L}�cdrc<��6��X�Sr&�1`0@�kv��.ca���_튍�0r
��-\�|���Hfy!ҟ*=1�H�Q;m��t�5
��n��H1��+S����Sv39D��~\{��`���|l`�)ٰY��[lL)s��1"�՚@�b.S���ߒV�7H>����A��$q~!Tw#H
R AM�����}6�b�/{�	Y���jH��~j�4��v�s���;=v��ߥ��(dվ�_X�A7����h�H�
jObWz� �Pzįg�t����ߓ���o5��鋚��2�ПW,]��D�$��
2�T9�VO�~hG��n�_�<�i8�3�Uˀr%'�bv�X�.u�׺�m�,uk��5J�zw*!�P���68��	���I�/G��G�����7�e�g��ɦ�(��~���?���c���P���5�Ke���n=7��b��8x?6��P���T�		!Y�$�NE#�y����ٮ�fg�`�%	Dh�ES�����odC�U����k�y��d9�Ϯj��CqXbxԏ�6C]wA<���c+������	��
���8ݧ�9�C&�ou�z��s*�]����O��\��(C�U�1ק��y;����7��.�M�Ŭ�P3����ǡ��#��^��Āh� J�Y+��k��|5�tR���6���.��ˈ�t��/�A �6�7m`�!XZ����}�����'c���X��H�I�"N�j`�r�ȬrH�.��ꬊA�w���AA}SH�v�R6aE���+m9;�V���T�俶����=�	>Gz4������ ��������*�hM:6���+��c�K�=��V�f�B��7��І����4��y�R����(&Kp@�p�X�����aL���/��F'����.��<�A`E=�����l�l?y���]I�Y���*�o6˾|�0߫�*	��kv����l	r�2��Zz9e}-�;/��`)��}��쬓�fn����JV9���b#��D�eA"2K��Ma�L����x�|����g�ǒg�ʄwW=Q��N�/�̿/W`��M�p�V?�����$��_Z��A�/o�s'-[vwr�-&��=�x�S���ȄA�<���v�z3GjH��{`�zU�}��#$ܩ�����~�%�c
�����W�Cf��$�j��ߧy �zTm���\��ue!�̷�X;?k�K��g�&��&1�<#���u���5�%afU�^�"2pƾ��c$� ҆Z�
�I�N�3���Z���� z	���� g��r��2D�KY%�m_����KO�Ftq�!���~�ېxn�~Uh|!���z�ПX:�6e��Fi��:�/M�����g׼B��11��>�5�C6����r��j�����:S����;�KE�s��$�#�aZ�+�����(z��Uj����A5���c�YA�Q�2T�{�R�b�@[H��R��P�Ui�6Q~�����N)�Qݾ�:�rF�m��� Lw��Q���ʮ��G̣	Q)�?*2֤_a��ҏ1�m�o0X[��t2��]瑴��{��+Z֎jYή� �DS8D��y������ �|����c'6���K�Z��������<爥&�\��I����}}�jȑ:�F� ���*��2���-��Zc�+����}�q��ӕ~7	�&!�AW7��9�r0�^����Uev EL�K[��§̭Ƒ~�l����)E�9�݀ì��Wp�2�k��eI~\^�ܺ���-msT��>���J��CN��%@��n�-NSg�'�o�υ�ݴK>𒳭��T\;	:��N�@�aa���[P�kv��1} �R:-vVǛ�7�C	52��w����uhy$� ��j2����W����X�嵒��*Պ����8���-\�7���>X��:<!o�XػC�a��G��
������_���Li�Ћ�g'�0�Ls��#-8�s/��.��<u�T`i���e�ש�-�<z>T���j�%��5��ԉ�~�w�eH��R����dA�%��T�.����js 4]\�YӒCi�Y�� ZV/S��Nl�c�?��j���c�����lC�V$�&,$���&* ޤب�������U�������}�g�d�������N����CЪ�>s��S�=�
	��Ҁ�u8��Ni=����{R��2*l�	ր���c}�y,a{ݖ�E꛻P\��x�cC�`2���(;��#��q�F�և�E��w�L�H��KQ��ߘe��d�G�I�q&l�
�=@�?n`;�=vMq��c�b�d����Drq,8�z��?��0�"aw���?UX@��	�"AQ��kw A0ᆸ*4oh:%��U���?���Tp����MT"�\$��4�}J�k1{N6+�Y��g&�\�?�" �h����/}�J�p0��wo�y.T�,�7�cZ��7�c��wE�-k$}�VG�o N��7�T)��aY�;<��,��A!|�ԻE���j�L�;���˿-J��;�}��B�e��#�%���Z¶-u��K����ɬaD89q��Ms�:��W%:��=bz�W��K�a��
��-qs���i�e���I/ƪ� ^"�2�@���Έ&ԧ����������\az�:�mٷ�-��]K�e�$^������cѶǑ���ա�� �G�V/}�zZ�/
��W�����+:�.�U�x�}�[�G��D����EW�`�|���V߳�)>8�2^�Ja�z�w��O�H��n�$��籇�aZ."��i�%{}?���!Y�_2q�0ѵ��Fth��R~��M�/����5����56�L�[1Z���v%�%_P2�oh��*p]�N��h�������y�{��O�<����(YM��e��3�sMwt���.��<>"s�J�s���ZP�I0�Xҙ*��[dhHyb�� J�tK�\?G>���3���pz����u�vs+���]T_s�Lc���"�*§����7��T���K.�ԭ ?0p�b�c�t ��N ��C�ف�@��i	s�Vg�"�h|h�	��))�����m�`i�<H$����$���z�0�Z��>1��d���I@V]�5h(%
Ҿ���D�|�{S�AX��Ꝉ�����$乎֘��g5 a���%����V3௽�v@��h��ͯ���?��9���E��6,�xc��w>��R��������5u�!���D:���F�x��wO�(`����s%�킋�L�k�����Z�^)�Ե�7!�q�C.�y��A���dZH�*uP�N��O3�R�j�/�M�[�֡�K�|���X���nA��a�t|~:I��R �]�l���`9��<�ڂ�~%�^�̹�68��l��*ٶҌ
]c�jr�<�
U�2�k�`E-L��!"�Q�mT�`ڤ��A��\���2i�u�m%���]�r�����r�D����b�]�%B?�k��s1�/�IW�qJ�t�S�Z���9�zV�L8��T��߲[)^u5�,�$�Z�jH�F(s���$m?/_����!�>���zV!��H��liZOr����]�X���V,�+zl��&� T[c=b-�Ä>�X��.��]F�u)%&���ѣ��
�����R�hh������#.����&��N})#U�[$��$�C�t�[l�r��3*߭x;�w��:a���#�DRT���0�v'i��;���7�\s:i�*m��L��2` ;2��GQTA&����5��f:e�cq�M����/�+��B�T��3���+�j�Q�O�K���e ���=�!�?�)�� �~�_�x��<��z���N�9&0�J��O�^� rC%�c*����,�������S���i�0��p�*y��Bo�*�u�Dd�Ynq] L�]r��8v��Bk���D�8���d���!#w�m�a�����&k����x\��̍^m �Z�yN]#�U�݂���ڌH|Ν��!$�Ȝ'v����b3�UrX��c���H,���ST҄�؁ .��ma�{�w�q�.諀g�/�i������qVt���?�J ,^^P�!nU�]���$�ͥ7�G9�h���	��y�g�]�I�x!G'�wB�t��aA���̒��'� ~�q��}�p���N��~ͧ�#~��<]����]�F4�r�!1%%<��y��� ����iL���^LU4"�����c��ױ�ĝ��M����^K�C��L�����#r��4�H��.��k\9@D��`P���ڂ�Q����i���ط�c��$��U�ܬ��'�M��O�ѱW'�Ba����Ɣ)+63uŅ��k�ѐ��~��8��MCK�K��	�|Xs��T��>�
�C�x�t��75�[���������5Q��8�`�K.�AQ�n*]jO/��^�q�&��k��L��{�������k"ĚҴ���Y��l�T�JM��w.�EJ��%�Ԏ픤RfRaX��*ioq.����q��訩����O*�6��II�x~�kRL)y߿����o=�<��CM�z��}�`��:��D˅�&#�1���l'���Rt��]���䎰�6OLj�M�;�1`?���'�
�C���3��R?O�� �)ml��e@�5�-�%�7+@-�����.���r����F91�*����th�V���Yѻ��d�Q��?��&��T�P�mE�c�ݺ*N��~Q�j���Jާ���2s�B���S��&� U懕��=��%��kl��7%B�����<CG� P���t����p�s������ AJ�~�
�70��C���������÷]�Zl9������4��^�ˮ���-4!E8A1Mp�B;	�ظw[Y��N�L^�.Zz;nY1���<"��
�'/�����9~��l=Mv9�������'G�ۉ*���YI)S�(Wl����~p��]��،��@�^b�+�����1�'�X񖘬�iȷ��;		�;�L�^��#�=q⠮ (chH�ݼ��[��w�%��ڰ��.��N��B�-�:>�]�l|$ݷ��E櫦vauM�X����m8H�TL��>E���p�¦�*���Yʝ����P� �@\T뼌t0б[��h�@�QԴ�=_��c���΢��V2ߋ���v:�.������>t^��j?F�_pu�YO�����
�0J�*[x?�=540�Ɏ1/ť(k�g����KAjCc�P��&YS��,�bYK�&��A6ub{�ʠ�Э_Q��������S%�"e���$V�#hC0E��۸:�5l͓���E��+��:e��J
�w���{�����Oɂ���#˲z����N���3�����'�z�n�Y ��>a�ƇW{��N���|PP�0�pYKF��^?��r`���jӃ��]�/rG�wt�gn��s�z�khlN��,qM:[%�\U�"Z�d^��R�b�i�J��􈂺���_�?N���Si�i��k�����x��"rN�9��l3\)�C�g�X��;�><��[��.B��+���m����g"����L��۶� \9f�)�U�N��!'ŝ��|�D�h$�4ͦ�G!��xw���=�-=e6�.q�`�gG��Wj7G����Ӕ��g�k����إ3۴d���<M[9��Z���t.
ܬ���a7؄�	"�����u��D�t��z�Yl�OfЌ��a��|��)	+%�m�;s/��ρN����t�$'џ��91��J�y^�V&
�$����d}�c�e9L�Ua���!�Y55���/C������R��}�g���wKL��.`r��by�+:u�����T�S�������;�ւ���$�4��)`����;�>�y^e�=%hF.&���r��%��dC)&k}��k|ד;Svk�ʝ@�����I�o�8��3I�F�J�ħ���Ts�|?��X�3�Z�n�{K#��X]��)��z�M���J�GI��lv�\ꧯ��w�m�8z3Sg:Zؽ�'�J��l���7~�n�¡V��D@��bk}+���k�`���.��+AE
Տ6�=x�Vi?{Vz�A$��ՠ���	�7��=��O�#�]�c�I�Z�d��&x�M�BZ׍(d ���{_�b��&�]`Rp��Z��a���g�a:v=ntY�F2��������HPn`����G6�0'��Ұt��6_��y�n��)��3�Q]l
$D0�z��D��:IOS0��("8�5�Ί�����C��gRvc8eBڱs�
S��N�8����A��n�-���J@#���tnI'[��&4Vs�����{���1 z�o[����<�:"�r>�^"�'_�nJ�'��G)�����S4��De��Y��4�uŨN=��i�o�0�Ӹ��B�OM�2-�}۬w�u�HϬ�k%����<�8�>�Mh,�����E�$�Qv^jM��v��j�}c�Å0]���Ą������>����ig��טݏ�	^0��e�_��5�œs�_�G�R���w�{_E�'����t����D<�!L�l�1������,��t��0�y��n��K�.'͍�%�\��A��f�*͸um��D$X 2M���ҧt���o���(�]C�K!�]�XKZ�<s��KQ̔,�ڴ��a�)��#i�Ç\�^�X٨I*6�ʊZ]/��Z�?*M@4�*D��Rt��:܈�|qq0ϲ��3,ӸƋ�3e�Iµ� 2�C�m7:e*���0Z��,ä����&	e�L�E_0}��� ���w�:����3�����<ޏ� w�[�Vg[��٘I�4U}��֣p�ʾ��½��|�(�+��Wo�_i�@��cs<	��[����\��\�R?���{�������(S�jۭ�v��]��xaP��uI�];ξ0�v����V����+�b�^jó�4�_���$�?S�͇��vq'���F��#@����ؿ`LX����	�%]�tQɧ������o�&�w�M
�}��bC��ϝ�WYF�P��}�z��oia`�~�7`XYO�`�^r⠾������+�Nx���管7M�� Й�T]	ɬ��
�sy4ߺ�S���J�w�)��_�ӘZh��|�]XW��Q�؁�oyX�*�M��Sa���$*���6��W�当��ê�Cm�� �=Q��J�"�W�IȆ�8	�p�r�V�?������5�ltkݥ�$)����"(��j�������,�<
bap��)J�~�����p�e	U��C�J`�ٻ#sE���-ɍ:u�A�>]� �K�7mDT刷��/X*0z��$��s�rBv��f�@�v��k��� �A�g�VJY��}�����X�F+߹���a;$�����3�H�ˢ~KZ3w]	](1��s�c��l3��52ں�;�'�7m����Vʈ)Q�����>$�	P�JO_�nF�������/>����r�o�?9����[�{d߶�
��("�τx�\���X�����bn8\���@�5��"[Ѩ��?T�нB�(��%T��������*��9r����dB�C���¼w!+�B���d8�ڦ����Ͷ�D.�\-ǑI�����:�EO��d���B?6��&{@3>$h�Vq���h~��2 \�-q]��q�3s����K���:���{��i\���h��+-��H] uQK�LZ����

��l��������%��m,oD�����)]��3��FXz���=�|0{��n����8��`Hr�mg�k�Š΍Ox�d����6h=�0��R�򐱔:�N摨�Fu�c�ۨc���xZR����f,���������f܇��=�-�Tee�N�|c�c��V��
T�T���1@$c�U_�[�m��f����:�l�`f̩!c~�^�Dk�;��D����:�nr^����� B�7��W�D��:7�|����Q�j?�z-	����	��i��}���z�K�8��p
��,��y�op�ɴ�m�����Y�1���I��yxC���δ����D�e>�y�5ߨ�_���o]뱂�	K�����\��@���7��Vo,(�Sy�J§��(Y��~!�/XS�v%��!� 0��	��W}QR=3i_�q��m_�8�~��~*���w��~���-4�?#umW�A(�gc�Lf˶zhj��&I�Q0���?P��'
[g���NC�J��aY�\���M�p�[��_^-�%��S��3��V'�Eŉ0:�]��R�D,k?�}�W~�6Ii�� ܒ�&��ve���a�Wq+������'�/pxV��L� ���{p�֫Au!�M�F�L�tǪ'Ƚ��4��c��]{j�W�����ko9�#�IG���$ Lo,%����S��Cu{͸Nj/����f����72������P���N��G��T��د�n:��Lц`iň}֔��˼M���ԟ'��>�3�/�"��r�)��*��5�UG�����|�pW�tn���ņ�,7��d8��K�L��e*�+F��Q���@_~'�C��,݃�O���vB-�`G����\�z<��������-w(�p&?"��:�uG�_��{hM�j��3�~2�ǘ^�[�8�H�Ot}�F�3}�+{���P����K�seU� �!�`�����q���>�7�s��f��|�K,���*�2�z6��@{�Ao��&�9�?�������-��h��`� ^R��|$q��M��)V�G+d�p�0��ˌ�Y�B�=��g�+�Q����R�Ev��T@���/�V��7�F������>_&j|W*?��!��Z�I^��?��6�����)�A1@5"���Na�i����_h��k<�ًD�@��� �\G*��I}�l���&(�zn9�x��V������{ytğ��5�
��:�ڦ�D�e.�Y��ʙ�B9p��d%ׄ�b��*ζ�`�/@?Mw�� ��@M@�BvO�̲��Q�Їo|�������?�̟B��V���kLQێ1�Nb-���}��׼��<�]��Y��՟���a�m�Yw�^af�V�[e�MB����Ƌ���\�׭�6�;(�w�|�kID���i�Y���"�gq�@܁i��z�B�u3�Hl����IiV(*Hc��0%����ޱ��x�<8q[�%�G8è��o$��릿R���PW�=���1�u�)8�nCq܍�ؖZ�  P��%,�BȻ(�W� �$�`Xj��u�u@>l�3�}�y���lL��<;z*igG8�1����E<J��W1�@,AD���n;R��Y#��Q܁\�ش�ʪ&�+�Uv3��e֐VŖ`��c6]%6T���m�*H���d��Ƚ���80-\޿���g�v�q�oy�N���	�w�i5�)�8\њ��&d�o��8=Z��nr/�#1��(���K�����M�I�a�E�u
�a�`�".;�*���s_ۿ�04\=� +�}H�F�p�;�p�(e����7[�6)$׃���<g�c�,��~�1 �^]���*���r��9��ړ��kr��b��i�փl�:�z�bo��aҍ2H��w�vND9��-ke�dS� �d����θ���Ks��z�	Xj���֕�;M��PB Ծ]�,"�B���u�'lq%~\AVV}�����ЇpAs��QJs�k\� f�,tz6vh�ݬz�dnh3���v��qZ�+2���
sA��b��̴i�F�p3yL���Q0�L�}/�^���xdI���h����i�TAs�f���ԛ���{j�P)����]�����X4Y��"&z������|��|#��p��u�J��j��՟>����&9a M�H�ܒfP�+���/a�����ZBzׁ�?�4��~P��1�����K�&��>h�{M��?Øx	5#>���ˏG�`�.��q8��J_d�%��/�z}�|9EZ.?��d�*V~,5�O�ڨU}�=���d9Ȁ!��;�MG>G��lZx�@�<��c��Hǒ�v�/Xr�f&����R�T�����.6YW.��٭� \O��3�^�ݦ*bI]VdT����#��nc\�����y�.�i�/F�7��ɡ�R14$��oN���Xo�uq�d!�e��~<�'�/��k�8��f7|́d��PRf��I9Z��k�đ�9"A*| �����(S��^o�YG೘ �n�@1��rL�PX������n�M����=7�\mE3[@���)~�����~�S���@���]�qt�
K-3�4sL-�A��G�5V��Vc�tCHg�\�|�l�pK����WC��E^�\T�����g�a4}�P0�XP����N�o�(�u�a��Y�����n�D�;ºM����T���p)V^j_kb>�{�İ���ܴ�����m���U�A*8���Yq�<�f�4����	�gb�#���0��.�S���/5ۡ�"fN3o0�Ǳ�!�i��썟܌D%6�T�Z�e)׏Ù#�$�}$��69�^�;��-�^ʶ��G:$�g�^�;�s0Y�<�,wփV)�(ơ)O��'X���p�K���_���������ڭ��Zx�t��O�w����ˡ!b٫�Aߦ"��K ���I��5�r|����`�{U,��֖�~�t�ցa�e���G���H�#���H�rF�Q��S�W��"��!@E�E��g�����7�j)L�~����̆��)��"�F`>*2X�1���
���i'K[�-F��(-�ґe[̪�\	����OM,�Y���7��0R����_�2[����ɮ�S]�j|�>[�3�>\�h��j��&!�r�/4���`������6��4�5�V�v|<�iGd]����a]˜B�	���j�1:6��d�gv��&���ϼ����}c��F�q�|���Z)g���y��Ќ��#N���w(�^o�܇�#0S��+�����1�'��D�xP� C�D$���O�Gվ*��sdV�A�bX��9���v܂W9�EI�.��2��5S�$(���=첊C8P���@�Ǳ���=��?p�Efy�/��E+/�W�s�+
�s�h�׿N�/����$�˳��Dc[�6-����(��J�'i��4Y��T&?R	��lLf�e~�޳0!��Z����M� �K���3+�p�Nl����R紉*(�m{U�,)�"+!q��
�r�sh��d��n��̫�d9MRUǂ0#���^����.O����uQ('�x}���^��Z�KMYf��P��|�z�Պ�x[l��I��� �ξ��%�O(q�p����1,���Xv��6�
�O4��e81��J�{ʧq2sߌp6#�����4J�.G,�B�����&~����~sh����2���HG�Y��q&��y �ֿ�ه?M����La|q:#�*vu���f8dQdX�=����W%��\l1��?�&�����q=x��t��[�tL����������o�]��>*rb�"�
�����z(�
��kp���c#Ǐ���X(̱1ݔ��z���2�U]>� ��9�h獅՝���f��V�zL�̤n[��+Pq-��L��E���I{Z�9����rkb6�A���J:���~�A
S] 

�@p�bfK�Y'�+��	�0��K�W�������V�m�qY�� [��i����Z6�{����v��l�h�.�j=�%�*��ۛ�!�8�g�;�[�x�J��=�9�ЖYѾ��>L���憹����I�zq�I�N��M~۱S��l�es����m����F	��� [����:�85��TLj�Z������ddr���ˉ�{Q����P���p�Y\�/R���%�d��~3#,�LG��=�����BH�@Y[ 2�?$�O´o�h�K�Z���~��5�R�SN��x�-(<��f��}ǥ��$T.)D�nԧ-���X+���fB, ���?���\[G]+����ٿ9��:#�rx
H����zE����xE���q���P�$��"��-�P��zq�Q��;D���J�QrY;���������u��13�%-e8HJ��	�2(�a\�G�AվSn<�"dPs�������8��J��z����І���CAk�jƓ�ۓ�%�孟>��ݗGW'�F-�`��
�3���p�/:���OU`��&�to>E����p�W�L�Pۈh�[�3���ϓ�L�~�<�6��� +�b���!� Qg��&��c"hyD���D�	t�=u2Z�og������wzb��eR+�Cvu-<u��ֵ��0Й-��Їj��C��B�=h��i�S'�녻ٯT�1*�ʱ�zOpԛ\�}�u(d: z}��v��;��M�c)��r��e�ҵ���C��D[�����^��i'�.�s�	6`�Ύ��3�]���k�Wo�eE�"a��z�d��S�d�2�ݱb/�"�0H��*5K��~G%���"��8=|E��X�lְ�|���a�tf!�>
y��L����u���b��7I���Gx�s~H�9)tb9ݔ�yK��f�H1c���P��'D�%j��܄�]��B�"��:	�7�
4��뎰�!�����&�t$�m>��P3�T��s��x�ZG�F[#��;��zd��ٶ��M0�>��+�c�V��"��j�m٧&8i��3��0�<ߕ�:���k=P�O}�������r�^�t��}1I�V����Ӡ�4��ׇ�:$<����z�D5s��K\w1_�H�γ5ͣC����Ge�'���p�-�:労D��Vi�k��8�4h'+fW�N���C��>�e�'TU���.T+&q��U"jgk �=J�vӜ�]	.�&�1���	��u[�/��nxe�Ms���P���v��r�+�F��eu�@�0@�*�v�@JO�L>���%�S�;Ѷ�ޔ�?	g�MӬh5��5�H�]w�26� 9Q-I��@�!�`���Ǵ�vBu��<�Y"V._N�����19;d#x�!�D*a���F�e��@�EBNf-�q��&G%\Ż�$�mC�-�'U��eh�4�z��}��iLG=�\��ò�`��t&�d� 5&g2��S#��3���k7���*i�Οm^+��b*������p #:xs�<�����h�i�r�'�KR��f��)o�/6��ZqPO������\��6���^^�65��.8]w�:}�7����β��ld
ߛ>����]���I��$�!�)�1�-6e$L#��_���NKmM�yu�-.*5�0�Q����"G^�%>>ϼ��/�p�T����*��F_�v����#��P�ݹ~��!�G�A"�W���2�i������BU==�ؽ��~�)�F<��f�r�m^���@ao�_��z,�^pa���VMꦂ4�4�� S'_@\PZ�5N۷6~��'��	�I2��n-�_���	a��6�������7K��k�6U�ځ1�)
���p)�)�cRj��Xo�T��$��[-�-�^��ml�-A�J���$���H���]�)0(@��[Ր�)�ƅ/�y��0�����ǡs�O��u�:�Q�,.�E%���������_@v�!�H"���BSj