��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��I�ɖ���˽�+]�Jf��N����2��@����甘������A5�N���n�nD����n���p�+^�T�������'��������c(�Lb|?�0����gb��o�YtJ��%-��8��7�A���*qТ��m(�ϯ��@�?1K����!�5)X�tc���F�:Ǘ��� �M�z�ឋW�p�{S_^9oӵ�H��и���=S.~��#�ևd�Vί�%���j�ão~�@����=�e@�L(��\�C�HO�c��;dS�3s1�)$FG#��h��������3c7W$9���>��|�Y)�[0�ʫBx��p���u~xݚ�C�<kdo%��	��u�>���]�35�����aRr�H�4I�/�>��#^�[I	%D��c#e���b f����ȹ�d1�V(�I?>���1!���k�Y��jV)��[�w��qjt������A!c�G��m$����)s߾^�_���]� Кg�||��-�T��YQ�ON5�S/�֨�$l�l�}c�/T$Qr4͛�O`��7��K3j�Fڊk�<^6������,%���W-?
�w�Y��u��M|�%�9���\m�:����y̭����(��r �n;k��	TG��xh���ȃ�������Xu&�GTdP JcdE!�F�;.��S�}~�t��RW��j[̇6��RV�+OP�W�1�ߥ[u27.�"E:�v�O�'l��D���������~Ġ�
%e�~�Pu#V��R1���7�^�ʑ{�܇��{yD5��5f��:�Ux��h6���⺃Y�5��8���x��c���E�)hכa7lkU����r��oA��>�\�U�Gp�\��5ҟ��SR��2>��֜cp�Z���=�Db�A�G~���}��3�ȝ��cH�O�$���K���q#D4g�Nd��D�Ó�&H4?��p�]��xf/>������!���9Gj�[����D�Q<�<mR�c*�x�gI�G�/F������b��0�O+�����{��gྴCs�,	����d��(�v7�������X�`Y9�5��[�	W���##g;���F(n���5<�[�9�����Mn�K� #a���pi)(׋��/��^0C���T�)*g���e0+�F�7�6eM�י��di!��@
�JA=��i�RdI�?���!Bi,���n8W�_y���=��r(7��,l�������8��3��VU:|�ĭi�L��R*Yƞ��-�b8 y_�O���l�����O�o��z��#�8��+G�'��ES7��|1�+$l��BX����D!�ꇂT��Y��� ]�+�Wl���B�����v x���
�<���yEf��l��0k��Q2fk<oR�垶�3k��������ѭ�)N�Ь_�߃w�:,�b�[PH&f��hN��1	,f�f��N��bc>�,���T�AÙ�DBx�-e���>��k��ؾa��jh/w�,p�R�`*:S�
_6駩i����eȚ*�[��5*( ���!�==k�S�x�w��K ՛��c��6�'��.]��l��0J	[l�2n,�^���H)C���4%~�
L�۰��$o��T��_&ە.H
o,��5{G�����RRL��2VKF� ���������d�F�Mӡ><�-����־h.�=^+f�3Y��b�m�,�A�o7f�!xx:���� �	<qn����Q�)~�D���P��E
m[��S:1G����0�A�o��!>��f�J��:yE�,��y��%u��*{ޥ�DόGŴ��?�S�.4�a4���:�L������1�o�#�����)u���X���*hUk���*��{��¯^�.͋�ډ���e9�n�.kp���=m�V�a�k�{�[�t��	Vd5��a��<C9�H`�b��禴?n $��[�≦N�c��@+�En����-�-��~�����V�<���#�����[o��R���/輜�@|�_�q"`�g2����0�D�C������FL���.PU�������"�3f<�*�o]�*�D�]������B��c$l�qy�Z�
?DF�飡�/Jq2qr$��j�k�u��0�`=�T0LUb ~!Z�D\���L69.�-h?KLPƐ����ngV��nb��o�;.�"����#�Mf��I�	�~}��W��RɷZS��f��M8ڧ�q��V�&�S�rm=K� .�~�i��.�Ϫor��.�DT�3��YJ�Q�2�J4�;��K.>g�Vj�=��!o�	��AM��T�1'r���v�!f���3I�'W�>}5m�E%5���0Ì�a�<��a�:u�]�0tA-Q��j\��]��3���.�t+�܏R�	��E����7_0�k���L�$,
��q��5(���c��Q��~I)���Ǫ�Ȉ�{��V�����z�	�wm�����}e~�5{��KM���7X��0�O�e0nZ��g%d^��>�P�K4�C/ /����٥���#��8z�<���-�����|�`�#��n�+�w��-*G��X��	�kO9`V1�j�ۘ��$�P�vO�gz�4�2�S�te�@�-��^�'�JBʧ�M��-�3��ϙ�Q^Vf|y����� �`�����3��m�ׅ�	�d}-�k �.$19��?2�L�v��N�W|a���؁V�� ����]��t�_�Ӹ��@���Q�?����]���mc�ZZ�dq���9U"���TYK�q9��~�_[ȯ!e�����s��E��޷�f+�8W�G؁z��w�H\��/�\���WZ�QL~`��U*w��9Í�*t���b�J뻫�[UD.#�єrRJ{��7���N��\"~����h�-�T�Q"=�4
!��>ލA9�Q�����àI�����\�i����H�Cs^���x����.U\l"Z1ƒ���[�E��;��7�"����:��f�@�Tp��;�w|�͕�Mh�ȕ\5��zK�O�R
z����@�z��3�h䟉��)�:,��'bPPK���4���V\�.��e �m�	�ƮT-�f�H�e;g糍u����&�kXy��:��}�?Ul��S�/`d9_e둜S��먪]Z����(�9?공C���S�H��<yGZ��$9(0�|I�4]�_UEG�Tn�\-H*���� �K�N����(�Z��A+4C�@����3�h��jhq���/p��y�W|Z�Y(���胶W0uWY�nϟl��i?�i,�_��R����L.���w�c�n9��AC��)��!��n���׆wdl������?�5S�����-��`!�x�<%� Ur��n}�ئ�9�����6*hZ�MP\*r�_��.�Ѫ"!"�roET�����qV"���>�����Z�lm @w�}ɀr�+Jm��v!�̞�{�6J}�-���^Ey����+��� ��
A8s�H�����E�����x�Z�;Ңk�X�brf��#���j���&ˢ��ORr��q���x�M�Z~cʟ4�a#���� ����,pQ̥�(���sl����UR��i,��a�-_`Q\h�n��׊�`PE����y�v~h�e��4��4-��@����"�(��[����s����vח����^�I�\��Μ��[�hh>U
��)���l#~|���I��xL2ȶ�
u	6�Va���/�����D ��ղ\+[��ɹ�y^�)C��7���H��H�w��L����g_b�4�\���X���1;q�ŊFs���s���eɌ`��f�n�vw��