��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY�%��sߓ��<k��OI�x[��<^Q��d[E�H0q��[�'��>Kj.��7���M"�J�o�2a�g��vQ%��|NvT�q�
&��W�m�E'��pW�zѕ���Q{W����vL���pU�n����E
yN���ݨWj]ND]��:��z��-֨�pX"��e� F�;��1/H�!���/�� (s���=,�A������`���h;�}7�t����oij��I�w�;�P)簀����F�r�� �!�v�"C�����PR�50�	d,THϣ�#���E]b'HM����3��`���TX.<y=ͤ��hc��=aV>�zF[�����r�B���E_?�h�X����KW+�5�-Ռ�̡�=h�%�3S�� 4a�S���G45��6��k���"0�O����#�e�f���x���')�0��f���{ܤT�2��ک�ߖ���$]qr�ǥ�π׆Ki�k@��5[\�nZ�g?�7��;�i��/^�gB����	��=�K��WR��w�h���թݻ����rAQho<R0�KP1����Q�k�2=^�Il��P��
8#� X�8�ڪ~���}6�C���wx��p�١A:�5]�{���Z}��^?zw`�0s�2C����5�d�W"�*�C�K�M#uw��u/Od�?ɜ䥓�� �����ő��]�Dl�U24�&��A��{�Og>��4d#���ٮ�R����Af�f���+n���%ͷq�F�^KZ�k�|��C\�@wy>+��J���U�Q��CW���z����	���# �y[�����^yE�,�Ja��ưg��ki��h��w�f�<d�
��!�|�k����x^\�
#�`�:��M�C�����D���h����ْ>o��'�(�I2SER�"� �g�T��i�t}z۰	�1���x���Џ��0IyW]�:���1=OR]1y�ɽ�M)����*�+���6�l�f02��%����j��K���씝~��m2�R�g�ö�V��^�U�p]��sۚB�ωJ�47�	����&�cp���h�*�Pv�#t�U50�3����ٸ���<��Y~���pi�	��M�F�g�EY�Q���aOf[sQp`6	��`{T����nD���N��ʐ~3��E��>��t��A���9�Mk��W��|�V��|�`��5����-8�^s�$�[�^9&�ptI�(��@x��EIIMI��A �V�V�^���[�ܪ.�����8�m���c�t�����J��
��΍}��QwG+�w~�g�D������,y��$2v��'�all݆'�˓'4"�x�:��t���_ W���~#����t7��;���@��~��E>[�{���K�4g�ˣ� ���X������Qߓ��v�8a��ƐXxԅёB�X��\�8B��D7A��rd5��Y�#����'v��c�ɍԖ���/X[3_#�_��x�3���V ��e��Cj�H7�O��G>���&�r!1.e�#�tֵ/�^]����&I
����΍�|��e�4�WQX�<�.����JQ�\�������N#���d�ܚʙ	�u@��y('�nTq��  ��*��cz�ZXJ8i^�a*�f�6����_�җ^�i�p&�3���&�c�xQN��a�C'0���<�0t�:Q.*�������	֪�'��w6�v̝��X�]���S%x���0'�u��R�02�W�������7k���P1��i���;�xu�F���l��{��raVU�Su�Q�z	"�P�ߩt)�4��m>&�Lںh[���Se��H��� ,5�pct>����|m��em�x��e;d��%��Ѹ�A~-�L�	�(��2���/�[����QV����M{�S*J@l���*K�p�iHR��0$�K��#�V/����c��ub�'k�ڄ�d�^6[�Z,��u��{������� �f����8	����_�"0��[�2<C�кհw>�����^V=^ !�ά�nt�h��Q?ʸ������k#h�.昑{��/;^&�W�ɴ�7�e>ÇRF�=�,�5,nR��BvRmxJ�����O�K�	���Y�~�̣.��-������AU�x�Z�'C6�.�������z.X��w��C� !��rH�`���C��2��cM6��~�TW����6?��D���%Ѝ����N����p�����|�.��~~��*�݉O���+Є��)ԝS�'�8��'�:��{���鸇���"7��H��x��^V����l�2Yhv{[z��Ţo����z(�sg������4>�r���!��B(�>�[д�L���
�Ι�H���;��`�T/9Cn��DВ����9�ڒ/DOM�$oA�ѥҀ󂮘>8@���I+����E_64��ϤGs*X� Df���v|@*����������~�r���\Vk�?s�*�+=�ؑ������$	������
��u�p2�JqL'%�`���]��~��_�§*�� @*+A�G�`�}CO<�S50�d��������hW(�Ӈjz�����Yv�ϊ7/Z#q��~��������ɨ-J�)�4�ς��5����ڽ-N6�g[�}MD3T���7׳o�tr��F�"v*}���%�/[ܑ� �c�<m:形Ha`/��E�aǢ[�+�M�-\JFbIB���̬&�[���TU�3肜?q-N)�+օ��<��-)�\\�Q�)X��09ZF��y1ʡ:l�ژ�x]�u�֘��$T^}X�KU���3;X\rr�8����C� �}�v4������V�[s��KY�S�6L����z�+��ND\z�%�<@�6Q}�할e uu��<�@^�g F�HVi���?�F�9z<Xِ)9���0q4����������?ś�~��	 fT�:�;]��z��^��  ^e��fI�)�a4V�h ���Y'��u�H��O�A���������F���v?���݆���o}0�zK��!�q�ɔ�=��_�6)(Y�T�'�
���j	Z�xa������~MFv�ώ�� ���+]��>qY�Z'���43�-��C[�2��`����v=&A<�#��D�{��d��]�jaFg~?pb��P��-;�f����)D��(d���!\�Y0�;��L��?���[D;�K��HħdE��9�c�:���0.��1%���WS�	��4j�{Y�x;� ��F�9IzX�`(B0ŉa׋Lա�3�e���
Pj����{���U���!�ÇA�.���-��!��܌�Nu��-" M��H�ky���=�+Oߛ���b����B��~���ţ8��N%�,��*m�;$w����Y�e���׊?N>gXA�B��A�*�Z-/ $��q�z�mrR�篙 sۭ�3w_"d��x������9s�N���R	��y,]���Ѥ�
Q͹��)��rX�_U�aMQI��<�dq�h]� y�厨��C%ď�~�q3	�j��H�f�(r=�f��)����m�����~6�X��>HMx�]��6�0_�K[�(D�؅��֓����Z��9���bjM����'3�����yr^Db"b{?���!J����p:�����%̬Ƙ���UW!&�o�+jQ�ҹ4D�*�MھW��Rz3Gq�W�S+E�y��=D��.vM6+2��Bk�a�pWg���ŠҮ�����l�7��$L�s�DȆ_���r�8/~ڏ%lW��7�:�Y$�UY����s�і��	����wݢV������S
jp��D��C��orÌ���(�Xn���4�����7�Vβ5��J'���'4*4�9w4����r����pz.(�	�4_!u,z�U	c�-�JP���cem�{����y�"gpm�r	�@�o��̸��_���Urve�'C7�n)&�_��l͠��ڊUN�|��nmH�=�����?t"�d�%���P=���K�EHy(�9MIZ������鯩�I�Ů\�S#V[�;��Ќ�L%v��ökp�3�<moB��긁�1q���}�c��P�ĕc+���V� #f
潋=o�
n:y��$�M����P�`U���e4�i�`D[����M(c��-A�w�3����i��3��I5J���"�<�����L��.6'J���sy@O��kϮr�p�Z]����Wa��"
>y�E�=q�aS����[�����р[���"������=	�z���/ �n�Y22����mGX&�w@]�
�0 :	%M�.*�H.�Yв	�߸��3c]Б�R>��j��kf=��������z=�T��Y�'<�m{ƇR��s;9q��|u��<�:�q'5�����3��3$6��KW_�$�'/��V��x�mnD�}�q����� {pU��u�m9��hp�×ҼM�ǡ]ٖʢ�Jz��RM�D����d:�<��s��%�8A;$-��8%>g�����/����P�<�JbJ�m�@}�$�u�-� �gI�lS�\�P»X���J�Ӓ��n<�j�:�U��r D��"��w�C��k���?���D���sU�hL�R������?5k8&�%�uEݘ����%5����v��kh �Ip�� ���@C�R1(����'�8#	����B���U+a�v^3�2<����b�Q�Yy~Ƣvy�~���-�����%�]Q��0ZB��/�]�t�������г�1���tWLC�u�]�"#�xXy�c�U��[jO�‟5�nНK�6Ҹv֥2φ`'.p�XC��a�ޞ �o���%�O4A�d�OP0�c�k햬nWr	{��B��tl�RBgE�5�:؛k����:�̄�M���U��C��	��8�71&+�il�)m{>Ռ���R� n�O�Z�ޓ��亏����8���c�iC�*4�V1>���ck�p�BwX�O�
��ra�໊��21v*�w𦰢�cc1�8Һ��gr��ᵹ���yt��*q�Tb��g]Z. ѝP�l(�8%,1FĆ�셴'�w�	(���>`K�|����k����V#�:c��_���H�{�7���n�A��C�S�9�虺e�� ~]K�F1��&~�I�V�7�d[�����KoB�m� w*a��e!��*����|D�u�>�~��.�{��q�����J`��:�IÜ����/Kn<�S�
��\*���ݙZ�C��b�[/'��)�Lh�?O�ᇇ�k�Q���+r��`}�X�I����~���6��*FD"�+��P�z�k�1��ә�0�M�d�z� ��� ��wX>���+��Wq\�r�CX_����$q<äCC"_`1�8s�0ӕ̶�{l,T�?BD����)^՗���-Y*��R���^����Cg�vfZ:�G��=F	V�k�����V���:�E�]�!d���C��.��@���<Et#*J��$'Y���U�E�'L��;I�\n��M���D.�{/�l�kUQ�� ��f�H\б/<TS8���@-W�"�/�����ܛP��U�I8����̗k�Z�xI�%ރ�wHJ�{�?>���\;|�ݐ��	w�����iB'���yj�6q&P.&$�w�h+�̓��O�� �x�8�cN�&n�� f�Z:d ���*&��oݯH�Tq06���\~�[3�?%39�C�Vع���%��T]y�/V��臠����N�v���l��墠` fjᖜe~%��<΢V��C��%��ؚ�n_΋�(�TOA�z�t�G!׹���+��-�Px���� �y&C���]�RZ[h(�r��42��p�p�DF���	�t�Se��)�0����#��$m�(q/t�[,��!