��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,G��U�	�oJZ�@�z�����>�� �F9!�/_g�T@_hm/a3^��(#z�dZ�E�����v�h��|���-�>bkgá�G�j���zA�;h��Ċ�k��ׇ/�gN�3ӟ����i�� ����4��m�"��]��V��W!��J乧1�u�M>w��;��
�̗�E����@<S�ǿ�α�7C��8��B�TGEM=[���b�#@sr��C+�:�]d�}��.��{_e[��9#2�_�IQ/���*���ڥ���Z(4:�	��k~a|jg��ӹ��dY+@y��k1%v�J��AW�m&kT��v��	���lT�I#-�T��-�L��kRv��ڄ������s��.����``uc��
���ˢc�����Xr�+��ů(~���,�k��8���3o���'�����tM���B��~�V�m^����n������Ȳ���b�-�~B��=4���
��.T!E�|��+7Ik�P���.�uA�Wķ����Jgd�,%��u R�*y��Ŧ_���,��I~��Q�I�$�F�����S�&Q����ǝ;�AS�V���h��.�M�����Ԁ��x"��Q=J�?8��/�Q4S�������R�P�#���C!!8(�0g��C0�\<:yg�I*�{��Ur�p$ʧ��B���\um,�`�,�n�w�wCG���ec
�O�����Aa���6T���`�c~��#���h��׸R����k:m��ϞLy;Y6�*V�ڹ��^ǣ`3����G����ߓ��N)G��pAm�ߐ�=����e�փ	����(��)	�a$@�3Oj���UqOe���[zC�V�i��5������޺���@��D�s����A����ZO����7�!q��h��>Vߞ��?�@��(���:͔��܌�oJ[��_�B[�$�M�"�|��!x�0�te�F#j��2�]!�	�gS�wE���iKP��E�[(�M����kd��_k�w~0��h�>!���I)\��4��[��9��W����bj�����v��h��T��ݣ�u�!��]�x<X���F��6��~k��1~�18Ӽ8zyX0rS�d��ƌ��EGƞ�q ����j/cڞ���6�����˯DsP��4zf�^���r�>?�X3
���Ίw;��(��mw!3��0g����L �����D��O�ћ�l��d\1�SO!0�E�Yp1~d���!k ��I�c�S/�\gΩtH���[i_,#��}��N�}���/��0� ��E�pg^�5?iG��v�h讗5���t��-��S��|7��vU�C�#�`�D�,Oc愕��yy�Tp�1X�A{�z#��4��I$ަ^��]�V{5,�}�2�}F0LQd�|����N���눩&��=j{��a4���v��Q���.L9���D�$���MkoO�@�D���Xb�y�NRT�|���fN�[�P+9Nڷ�~{W���,j�_'mK	}���c� ���֜����~�6$E�z������稼I�PS��d�+�\v4�������J�[OG�U�p73�m�]LIŧ�K�Ȅ��A����,�+�����+-��]���� �ۭZ�4���g�ӾЈ _?�8sI27��mL�o��K~��w8g<^�}A���+���^p��m�~��񹛏_%��ȈeVth��� ��p�Kvӓ��(xv���"&?4bW��mQ��	���&���aAeL� ˈktu;�}vEm
꫼X��W���	�C�MM �[����б@ Q���+a�`s�D�����Q1�l��y��ä�����J�C���9�vg�O�[�.�U��e�}��o3w���TH{!�T?����=�^�8T���s�<�F#���%�#6{�Ġ d������'y��$�]��0���av�jAvi�	���祍��9R�2�8�$�p��Cu'C������7JB#ph8͔qt��~l�)~�exsz��w������y��Lv���\��L㻢���W('Vh��������P�5̊4Q̄oa^Z˥�C�+<�c_�5r1d�CK�_�|u�D��nf6w��a�H�Ҹ��Ċwn�������ᰌ1B�V�C�$��r_�]�@A�ņ-á@���W���%�	��|�:�����e��\$`�����1j�������I�����V�Ăk*S��H��X�B�'o�$�I���|·8�re}��=��7��_�c_U������B�>�:�]��A�Ɣ���>����o.)�ރJ*JH|[��k-M���B�}�r��7�� �QEf���P��ʘ
�yD҇M��/�+N75�yN��6�	�emмuU�>l�E@9�h��aT�5k�lj�~b��_'���tw�� H�z<ᘛPHD�cA0�x��f���:��,c��Ȉ�yT*��ڸ3�7A��!�73W1��Y�V��2����]v�t�16�&)TgQR�1��>��LQ�1}�v_pf���m}����p1���1x?tg=ڴ���W��'�����hN�P�Cl��k��������(��a
�7�Ʉ!͚��8}D� S1����{�SD�G��Z��D@�T��/��B�}1��ȊZ�:`gwj�!1O+�KL[y�9�Kt���j�B�qDћ5�S�;��ھ+V��E8f��9��h=p��6\x��tg-%|~�{��l���_QB�ѴT�,��Ng��Ey	4:`�i��M��iK�+gQ�fo��֍�t�K7�=�G�NJc?��7�^ӃD�܀�/�nwj�ED��G��e^�S��ř}��R���Rt�B���y��S���K�T�ޚG*Y|�c����X%_�D�&�hA�ɔ�'1�i��fXX��7��N�<V�e����n;G���u�ҿV��5x��(�6ʝ�DWO�r^���P���x�d�0��Viם��.A���c�И��Sõ���ڝ~/,L�dE���'�[�$�ړmY/V�Mo^�Bj^��nȻB�u���͐�	%)��l-}��j.�0rb�& �s8�z@R�xK��%I,פ��BC�Xa��A��"e7��	7|<�,!���*�d�Iϙ;�]��
�T�l& �V�<��|�
��,Kk����(�mg�s���E��_�J|�R�M�I��7�ԓ�x��lJ�2��/t�Ut�;$�(V�!��D��R>��}{k8�� D� �n#��\.{�2ᷯ@/C�Cx�+���r̠.�^>r��A��R�M�Wi/��V�?��v'�A�����T�ӫ.~��wY�[e�404L�/'/�9|}`�^\EY��0R������[/>C1�f��
S/dl�4U,�a���O�g֎�8���Meaۨ�^D��1;���iǇ������*�6c��fqpK8I��c�.��'rS[��tҩ�-}a���T4s��ّ�_����R�vϤ���n����d���lAp����w���q����&c��$���[���:=���g�L"#�P˯�M�7���(!Ջu�~���þӁ6�%�6��b>2*�w&AD��%2˾�t��_�������:��c���(�Ia�v����:n�,���9�j���cf��P�ݙ�S�	 o��g���C��W�i�m*��ʣ<�#ϔ�`���������l`��Y�(���뙗�R7u�C_6A�#&h��͉����� 	��*�R������