��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5����Z�Q�!�&��^�����'Fdf}uQ��z����*��>1���	��k.A_wa���Dky�G�#�,��*W(<�����%����۲Ȇ�������J0i�}6(�� ?Rvt�=�8{����dR��冖�kx�BZ{��$̐�,�?AvvR]5�Sڔ�\�4����j��>,�5>�-������E=���Q b���k��s ������c��Y��E�̒;�[����5������A�k�R�U+IM�"�JGp��w��Q*�|H��2�c�o��MP��P�W�-�0����9�Y�� �~~'A�wёO��/�ϧ{%+�)�8�B�F�H��l@.��Z��!;OJ�R	(� ��P���P�C���^���J�yӵ�����)7�ߦ/�L�������vO5ك?8=� �$N,�N����C|��(��-����l0M��Hs~��d�#:/ ����HjAEMi���~������1d;�m	��ԢvO�|��H�R���v�ta��;��j-������6�,�Fj�Ͽ��9�Q���T>*���	��B�\w��������!*E	f�z���݉�8̬\	�v�ܥ�Bf��PO5d�9|�.��e�E�]��/��F@ķ[��՞�Ƥ���RXYb̹�}�4c�:{�U�m	���	^�.���o]b��BZ��E��V0��+���R
��6��������פ���N͛"��O��	��F�Z!ޢ���Iȃ���B���0� �����J�T�2nu�2�M�)�!ł�n Ŷ��t���t�����M(��'�sg���g�]j�z�ɿ�e�얱g?ջƝA��Z��: ��AA Y5�f��M2Um'(���ρ��R�e�1����L�<vU��e�&TD��9��H)�2�V��{��%g��kl��[���)t`�ȣL��ni���8Ж8
ԓ���KS���4��&6�������4���~��`o<%�!�qK\_< �8��.�l��u��$a�v���i#��_�0��c������
�S�GV�ْ�	��k��vT���0jZ��#>��ćW%�32?��m5�kB�?]+��V{:x�du53"���Y"|�>�Mny/L� |��c� wM,k���(&L�Z6�X*x������U�IU��\>(hW$��M��B�Sy�0U��w�)��_[a-�U��X��y�V*�����T�.��~uK84BIf x��H�?���=��M��xU�&�fc��b:y��6���(�ޕS�F�{��g#��e���Z�㸎8ҵ�n�g3qD���/�ĮY��۵���kk,Q�����U��|�]���B���K� Wt�u��H�g�D!��>�0�����3|i�:��I�c���#��
�J�[�'����Y�����uH3Tt�~�~�'�b*C&&#�l/WVի��n��=ZZ���D�O��T�-6`�b~�F���k��@�`WQ�i�g]6��&-J!7��E��B�	ܡB=z��꘩X8A��x�tm!(��l�/>Ԝks$�UI��I����"��"a�G�`WNP5Uس-����,PE��J"�cr��
�D�����R���H�jm���q}$��w�a+6tB���QϥR�3h�s9R���y_�`��͸�O��O�V'�'�����R��9`4�q��~ĸ���7��3��iF�<S޽2��� wܐ��>�mK��㻇������~:��5��ZNi+��(As���zl�(ϯ�/;Y^���[���:�E9K�XB5n����;[��vn2��_g�K��TJ�b�<�i�io^e\i�ڱ��fN��Le}3�T����1���8VKMξ�L���_9��i��1���3��aI0����{hO���^�D�=.L�.�U��Z�fw�U��Q%d[Ep�YZ�g*R��"[���7�����+Ȫ�Dի��fk�I���v�o�
c5d���u���s������FKs�uG��°	����=���*LX�6��!���ӌ!�Y��� )��&/���;��N���us�14�ξ��X��!�._�J+�{�,=.��d3�,?-��/2�D]s��8D͚�'�����C��ĥPd=���$��h�2#ƕA�U%{�)�Ֆ��4�̽�� ���ti��+�hU���n��)��l�I����Q��d�@�W4T�ٙ�O0Ƅ_���	�P�v�IٙL�K.�&��y\.T߹Y�4Er"��:�i>�U�����4+y[:%��
[.3�T15TF�r�V�^��+3�v�,U]�)C�X�8x��i�Hԩgb�Vl�*��L
�=vb�����X޷���5��`�I6rX2dQ'��CA:���B� 3���q6l"���|�6��!ѐ�v��v�ͻ̗ALHE�}���v�1=��]ݮ>c_�µ�GU��$�����-��������q1>��BE�VR���$2�]rq��/A�베f�qA
�TR���3Vڹ�5Z����hq�A�0��z�i~mv���TЖ���J�C-�1�b`ߕ�f���>�H���sBEm#����&{ї��_#jowRІf+��I+I������&\�t��W��&����#!L��P��E�2�0ƕ̜�Do�]� X}i���'}��U��b��U��fS@�2��R�H���Nm
L�j�*�IoK��{���w�^i�igL�%&W5�����9? �v�|�����m��e��!�|��HwÜ`��+��WF{v�ڶ�Bf���@�v��T_;V^YU:���*HT�K �� �X���K٩K�/���5L/	�3���k�QDk\@��C7xQ ��ʘWcĬ�$��\�@�k*Ex�W¨B��R�=��$��窷��&���A@���h��]�J����)%�Z;���sd�����3���HOr���J�}��YG��˺�l
�٦U�Ю��<}�UZ�n�+O�(^?w�̳ni����ꛖ�:��@��>
\~�:h�N���[��::���i{�ǅ��o��>�����|*{k�Aׇ����s菇�ߢ���ظ��#����?��x�>2��푼���շn�@�!=ƹ�;��J���P�͗�LF���*��)���A�LɮJ�$�hOY]TI�&��1�H��'��7C�o��a��S��`���ʎ�{n(��=��E���#O]��TPY�����sf����ڂ$u:�x/�C�X~Ez�ub�^���/
p�?��)� JF�[�E?�Fj����C+lR��*�;Xϧ�s�̽��ܡ{~�r/m�:Sz���9�
�.�5[SB�_j[1v�B���dq�)'����47���W�U���fo2fw~�-�г���P�����X��~-y?�0����裻����)�%8J3�>��]8�����_�+㎂�1�-���6��m�LZIf�f�q�V����>�?F$�\�+O,!�x	w!a���%Y��/�����;�6$3����k����V�.j������%�8�`\�w}��K$!N��b)DJ��W��({!����`����{$��Y�`eW~��U�~��j�y�r��V;Hm�,n�J�W^�Lf�6b2p�?��V������U�� ɞ�D����_"8�@H[k14M����d��ƺ�ܙ��Ȁ����}xƷf1�H/4�N�mͺ��Y�!�@�Gr�8Q�js�B�"�b�4��9E�����f����_4��8����L�zb�L}���MT��E�n��CԔ�ь��N���݀H̠�������]U]����ov Z��p!Pf��IMqU��ʊEA�cq����(���}�pI &���[���#L0z+���O�.��ܻ�k�QV:ʹ���g�ߴ�C�tJ|s~�Z�G��J��R��D�Zg��q���̰�Gh��q��U�mt�[��yM;�UoLH�Vݾ��)���P#Z�3z��@�n?,�ǿ'���r��8��H�9��}��@�G��(����z�%��i�ܠ��hk���י��f_Gy( �4P_�c�]gf��W�<�������nldx9����R�CNF|7��a;� ��V6��j2R�?�U�NX��ܚ��X���� �R���ݜ� �ݖ<�;> x�M��u���]
0���7��s�<���㥏up�m�/���[�����|�'M�J,�'���01G�m�݉��8�ݍ+���½e����T+����s�ʋ��Y�iK��c���_�����Y`י�6�骾��`<�iO��v6T3(j�+f2:S�)g�X��fȂ��6��D�En�4޷�J��4s��fc�0�`%�}}�k�ڼ��E:A/�iYA�'�!��Ӟ��Y�Du�a	@*1$A�Cs���w*pgҦ:͹{��4J-T�)��R���-�����p`��*r�������I��Rk��v}[�)*@XMI���C�{��\����]5��bm�
�V�3�HV�I!*�[�ϸ7!��������mt+�(o�Dh�N�����g���w)LF���{�-��Ax58�a��8����N\Vr�2,�>:|mD�zJ��c�c��7��&[�Y<*��ӛ�@��d�k��.�SH�Z����"e+��J*��_��=7���Ul��cx8\��_�_�,>6�?���E�n�C��F���|��ݲ"ǳ�>V����=�j�{qğE�LB�B�[�3���ϗ��P�o~���F�7�m�TW?��&X�P|�_/πďn�t�;.���.�R`eLJ��9�,7�BKXm9�n�=Y��8�<�^Sh��V��׫Q�_�s�Ǹ��f�z�ߩ��sq8~}i'�y��n��2��YG���g:gQ�T��j���;������Nir`�e�.XB�Z�4A��wU|�˥�B}�ғEKo<F�W0�b��\P#~Js��)Da�jO��h�ݭ��= F��_Ě�텑�1�O'���Kf0����v+M�J+�-4_���?8'h(�L@g7G1:�|M��:5<Jf�nc�i��t��ey�U�
���y����iq�~"GM�@B	��޼́٨㒳�L{�I��!:�����H��<�~Kє���T�Hp��M#F!���eWP����v�f�M4<�:)%���:�M�����m=�F�&���v0�V}��;W��(����֤��� !%�-^��:��@Bh���on6���&�Kˏ�NP>#�#*}H◍q@H+�]6^���²�m�a�-�H��<��n\R�#�r�B�G�N4��?��� ��n'Ŭ�e6���sq~����|����V�_/ i���$pt2Y}�J���e�������:�|�n�N,�(�=���=�bqg�,�2��٭��..�ǯ����%Uh""�
-x��c�p)l� �j1�3�g�z�aN:�R��\��t'�����ʤ��sQ[����9>J�nP�<��j��]'E%�2e��.�,�̖��-��q�T���hR����D�X�����ZHNi�G  �@=��:&�4��p]f�/JK��]��[�J	��Hb�j��X�����3.Nٜ.��kC)�|.0�2p�ll̅��H�m�q�U�Y��Y���ɋ���B׊��3�{zۊɁK6�|\��V��+}��N<�A9(LD��v�vߪ1�3�J�Ő��j�����Ci%?�cf�&�Ca��Ф���i"����񍝲gҡO��p��m�8�E���{�a�-kGf%NZ1&i���T2wR�Έ�u�`���Ѽ�C��D�{u�W�>�΃t瞈G�� �C9:G�?K8��YK��"]Bq�b��Mv:A	�{��	_D�Y���B��C�m���)TƯ}p�`(1�h���F����O�7�:7���A{9�2m4R�!d*{={C�/k�+#T`^F��Fy�����a��i��]�-Dt�(��-qѷ���o3�k�<�����~
���,��T�*0\�]f����4�����
����Y�x�R^����S��[Y6fB��4��2N����\Q���N��!ט�x�K�p��][6J���}�\�)6��H���$�vFZm�vv���ꁎ灮i!��u�m�+��G9=��|�"���4]��_��>3�S��f�_���9�m=��v}��Ղ�� %`�4�����\�Ƥ60�y�	B��7s>��꒰E��U·�(��ɸ]BC7~��j4f�dƤ���r_���vaxZ�=9��D�|��I����G��uF�?���p�7Ne���#b=�L'�Ց��P�:�%Q#��'�a|v���0M}3&�
�ڐna6�[�XV��i�&֜����,�H2C�ˠ~��kn�c�v{�5�սF�L }�Q�E��A�}Y^z���ޏ3|E? )է׫��9�$�/���F�]s�t��v�i� 8'1M�2h(���7��B*���2�G�z�*�����"�`U�m8S[�ܜn��=6��D�'�큞�;YG��e�gZ��a�R�A��۞�)I��^{�Q�o���y'�;5e|m��m�v���q	��:�?��5�>-�h[2�B�}������vH�;�y���i���Z���k��6Pw������G���hFwOAP��>Ȕ��P�O��eK�pS�}�{æ2���e�]�VSgDc��1�ʠ)'[����:��j�p� �� ͙@��s�d����0�,hF�(�f"�9�O>5�Tp�^?ܑ�{}?zA��߱����^�~Aq�>�R��+�I����]z���g�H'x��r��W��Jy�P�h��:�64����J����{��R���.D6�*W&y�P��@����t,�9`�z��O �P�uP@�T��r��8:S'w��S��/����>���rx�!<jp�y6߹�M*q���j�YD:�:��L��E$���tS{�8YQmV>��q4�S�+G��>��=~.�.qP��k��)j��� @UΕ��6Nz+<,��m�Z	c��dć6���1����t�Z|=�K�gk@��.Z�O�x�G��VZQD��+,7䛽'��Dy\۝� v�ݯmƉp�Ē9'�i���Ð��{0�ޗn�*��T' �yN�[�F�����<���
N֤�}!s�<8�֓�B��6o�*�f#�PXb�z�ܘ��M�<L .�����s}��؎�&(�5|f����X��U�1�XH����,T�M�s7=���jw��WmY^�pN+8~0ϑ��+|.����y�~/�� ���5�ҷlt�[v�9)k�#i��Ҽ�;˨;��l��50On�����#k�"�+�?�:Y^5(�AU��]����m���!��
�E�#v�	b>�@s���a]�r*�LM��U��+�-���ӟT����Qm�A�1	�^����U�'����+�\�/�7Y��8_�Y��id q�ݢ�K:�� (I���$��-�ί�0
<o�K#`�`�L��`�A���&k�M�O	8&�E�(mi\�Lev�Ziej���L���K��� ��� ��믛�wxE6�O�g�u:��`숭��*	�˜}rWj��ʻq[��.�'G!O��՞��D�	�8
��y#e҃)���ɔϐ����Iݶ:B�������h�b&���ȊxR�������1FmGs�O����X���k+�
�}�{y�傓�g*C�}n�AT"[�uG{�^w�����}���V��}g�݈��z@W��;p��|�mU�Uq�:h��%j��Gja���/��v���,8���x1Z*ۛ��AO��\�UK��:U�vXÁ�M���<=��O�'�����|k)�U}��vҐi�{d&��ٔa��I7'8���kXbF�?Ǩ��~N���"�����	�"�$ܓu�Y>X�nc��>����͚Oƞ�p?p��"^��}@:���S�&��[��l2�y��D�ԟ)�Y�0�z��^+�������Swr�}Z�2��1 {�di>�H�R�,I�e$a�PA��)�-��^�@��5٠|�g.�rN0�,�r�`�W���:M�L�F洞{rc2$$�ª�i@���U���b�����͏Ǒ��ó%k��N��%��n΀P�j��l�`���5��� ����Z(w�"a�� 7?�+ ^�xPK�8�aSBiD��N7;��Ħ56*]U�B���7��MpG�\�0��-�ύ�s��f'���3bkTز��4�Z�0����y�Ʈ/�$Ლ��Tk>����۞;�����+��cÎ]�R�_!yl�����%��4pIx���R�ɪ@A�����i*�}5!��J2�׋�Ym��,[��9�!���X������z��-�S��ß<��XX&�|ﵝ>������
_����d��8+�Q�����m��b�����O��'JHߜ���:bL�{��ָ�EΡ(؉"Ư[��S�//�#��Us�7=KY���.mڄ �8osl������k��Z�0\��T7fT� b_?Z���n8.�A�p[P�󨓩KM�[���V��ln$�BLyB�ټ�q���B�Hn�XC���F/�ǟ��4��s
��r�#{A-A��-ͽb�-�V��Q��S7����-��P�bt"�3�7���!�mN�
3˘�b&�l�+��
�6��	��,�4~���Р�E���T׳� C�	��I�z��\��M!�����5D��9�?��O�e�� PpLw�q,⳽��F�0Irg��}�p���*���5����^M�H��~�V���X�c隐�!�L1rs�}ڿ�X�֣
P�4a"�V�0��;W��D8e[�k�}-(��QV����Dx��J�x����$��(��\��[��� ȷ���Fߺ��
F)�t��7V'!��p�*'@$����O�1��$9v�
,����A����`455C���x�7��PtQR�m� ��+F��F���u�:��I���'l��r���_�E�؎{���#|���ɢ��0�K���mGh���k"�8iO��cz,���h�ܼW��mi+�����v��"Ϋ>>���.�r��!���w� _�4!�������by�13Ŵ{@p%�Gip�Ď��%��-O�~�Ib�Y��^�on~h������� �^�ԗ�gasI3��$v�@Ϡ8���K��3n��v�uDs:牥e(Ѓ���R�@��M�/� �Q\��Adb���s(����Гl�IOͨOh��".���7�8����'J��^2=��K�dw�V�U绌O=V~��zo�}w�5�Qu�;&J��犀�t�y�G_�6_M6�7���o��D�ttq�J��ău<���*��,�U�R�sFݜwՏ�(L��6
�
�:�6�����ȓ����H�-���6��U^2���{ȍ�&���cŚ��y�ޝ���#vp�P�������{�d�P��pG�5�
�$F`�,��J�����f}�m3��T���f�SOi��[4��}ܱ����.<�ٺ{C��H.�m��b�(s�M�a2k��k���6��F'E�6�p0?yg�t�%9�{���äW���h�Z���G���;�U�b���[y��Uj��+���;6�J�B��o�GԊ#�:�
K��3r���0%lQb�2�O�n��g�2���!��.Q����J��Xxœ���Nkr�f5j�#N	Z;j���Mؔ�������uł����>���{_G6[W^�y
m�G���x����I�5�����J*�Ss�7L׉R%��|܏Q2�;'�h9O�Q�bt�4Oi,T>I`{~0H�
�7�dU_�.��s�)�M�/�兾�mʠ��f��a���Ka�D(�v�Cv7�:lľ�Wf�u{���f�Qd>�������H7H�HJ?�1or�g��r�x�Ϟ_!�~j���I �ٲ�x0G.��/�Z��8q5����t�/��� ��O+��v9�V��.Xuf��)�%{P����R�LN߾]�MnP�@�p�/�,�-E��2aQ�ҕ�'����79��=� _��}q$4��/����J�S�q��� �-�3Z'�t�-g1l{�xs
�nf,7���~I�lu�T4!(Ő�f�ve!����>����O�f��"km�<Q���1j��6~��}���dO5x.a$� ������7=����B�����.n�F�E�WW�.�}�u�*ֶ�r&�T0(m�.��.�%��'�ä�n�Y�A������~+�H=�-�_<���H�˶��͟i8	㙸l3�I|ݑo!�k�`�{\FA�E�>�-��05W��e�olF+�,��K�����r��r���#���N�s�)A�0s��n��y�C
hW��u��_��C>���5U�vΖ9w���r��IM0{�4B���O�����W9�Y��x��Kɂ�U�L�?m|*�����Y�����s��a�D1�)�?��ǅ��:3=sK�LM�����,����,��F/��k� _a���{�����G��)mӎG�����H#���IE�F��Y�6x��yM�O�F���3gr��A?=��d�O�u��ҩ2G���P�]v���O:�tA_���b��ؖh��t�~����j� ��h���mhX�a;C������!�e�9����gS�ܬR�Lڅ��o��c�]�+���ECW�q��	�lx!T�٦��*�d��T����g��B�TK�t�`����q����;m��HWx��ح	�NHpY�%��� =)ZS�/�d5��D��DK���P ��(��[�5.D��l��,.�Xc��A����ErI��R�7yED"���[�3����%��0o�=vӠ�۱�[Z-9��+��1p��e�9��p���r"��Q�y͂n���k��=����PA[��0�B~�<r�����F���ú��C�V��ؓ�27^M/�K6W���廻�]9��>LУ�r��	�l0zS߇u�e�1� J�6�;0�},�Irν�:$6�2�p�s��q9�TiA���O�跒����`�اnOI��;Kc�M�~���|D�[�K���V#�Cp����V��h���}gI����m\!g����=�>[��� s�;p�Ajo?k��	%Q񟏚�6������0$��RxĠ��-�O���E�Y+t�|B�ì_�&y�o5Q8iF��=c�-��8�&@��h�BFDe:(�5�vx؏�o�Q�F��Y?�s�.��NU4�į�%��.몋n�s��ֈu"�0�t�N�����RN�SS�[�m�
�����[��9Q���p�c��=�7nQG̊
K�qa����i���@x��q�l�} ��{h'G�tk�"oE��'��t\��'xqѠ#ǵ�3[T����Yð�.'��\�;��(5hc��
�ů�&�-
�G���^7v�j):��\GS��㜨�7�}�������j���?LF<2`t�e:�L��{����嫤�#땿��i��*E�a��=���ЅDQ2��}�6t��AS<Tt��50c_����R���/ZJꔃqB���]�m=�,6_':�(sheb35�S�g��|�4�)�%T�����m�
l:��UC�h���3���`��ɾKh� 2萤�L���:�ꓶ:���u�F@Һ�ؤ�}�/{d��\Y�WC5�̒T`�%u���XV�.}�:�G����-a2��l������KLBÿ�#-�I�J�|�b���ݩ9�O�B«��B��\;�no��Nz������8��Ģ�@��[�b���h�K�C�4�͗�\�=� ���K"��|�J�ш���'Γ�BJ��+�ΨK��&~�b$1p (}��o�Ƶ(J�2[ܧ��HL\��#fC	6V�1A�]0�Of�w?�bO//�3�Y��~.������ae�ӝ���9����śU�Us4�������x,"���j�$���K(�䛣�΂��@xʣ%�2���y�ZԪ�	��R���K�8��T���*���B�pз�k�A�F�u�ߊF�I����Ѱ�����>J�E�����{���+�5���6Э��J�N����z�*��m�ac�l���{9��EU��k���c3�z$)��9we���%��5A��jD�>��Aq��F�.�m(:N��];t Mu'�ɀ����y�Au�'ߕ��3�{��G�(�vei�Yϯ�,�*�$��	�^�U���l&.��By�{����WBue|��@
,<Q&������ב����	Nf��լ
~��V�ޟ)�Sꃸ�z������ݕ&���iq8�c0�� mƱ���~ܡ���y,e�Y���AT�����^��x�1{ậhi�x�B	��@�5���g�ؐB��Zx�+G�59#�1�?{V�`il����(�8^�a+AH���mhFrF�ay&j'��/~u���!�������{��߉#Ճ��n�"��&�f 2�<5��}��gv���}ɇ��*# }��P�|�#��|�s����������Y��<��)�>�m�*G�>�}w����Vj(@�Y.!��LbAyn�z*�.8�ё���q/����pN��׫u|R��At;_\�� /b1�4cG�`7u��-o�eј�㽸S���R\��ߣ0���l�z�3W���	�EOz᝼��w{Ho��(8����$����Y���J�:����uK �����H�<&����nuy�Y�(C�D�e���)�!��M;M�~�G�����sD��[��~5I�cN�Sd�?����QVEpO����:��b�+���(z�#�9z��3��0�����oj	��:S6�%>��oUa����b	Ⱘ/��,~ُ��N�HLfVt����p�>	G�����2L~�.���ѓ�c \�i��;mg:�_����>�\=���L�x
Y��V���00M�r4���M2��!1�	��P	��w�S��l��1�/�����@b9(IQ�;�q|� 2��̥��P�_D�u�y銋h@@| ��DàM�o�S*�q\�#6)�%�ae��맃Ccl��F�J��.��\8�G�%yL�jN���-*|��}j�:����H��
B��:�:N����,6��'��|�_�e��qBLZ�J˽���.n�^Vf�p�|�O���K�>_�s<��ej#C��QҼ���MO��R<s��Aї��C�JW�)|HD�e�-ySD�n���'^�7��m��{�� I=��L
�|�'ʏ�� ��Tw�Y�oDc.Q�yz�~�,Ky�Դ^�<���4��D��)A`05.0�K�G*��\�%ŋ�6�wj B�|^H��
�j��ed{<�]�ųJ=S��Sʕ���3��G!`= ʜ�e��Z{����y�A'�;�{�0}U�jL���Y��=H��9#���� ��M�0�ɛ~~�-���'Qe�.�-EtE,�{����w�Q��}��"`����ZF"���#���)��D:!c���>�:X(����4G�uv��F	8ԶV9s�y8���m��k趷�38v��9<}���@�ɻ��Ut���)W���C��F]UQ�
)P} ��ͥ��i��M��Äψ����[��ɼ�ɜ̯��.�T
M
�6Z�R�Zf�nz��E�G�'���)_:�̦�������W��!� �9I`}��H�$��8G>Y������	�>w��aL���*�n�kg��������qIu��C���b�L��!ށ90u3O��?�}�M_͸�#�w�(�c��(Ŷ����Vj�UŴ���'��5,����l�Ve�
N����G�$0J����Ȫ�4zAp,��l��8��#Q���\Cݣs����iZ���ׄt��Yty!jZp�;b
�J����'t���K��&�]�XJ$ŉD�K����}�d&��$Ê��r�f؀��/�k�$��M��ٿxX���� R8�˂+�,Fi-Wqm��t���@ iH�HY#��X �F��t��>N���j�Ⱥ�O�f�J��mV���O��������Z�Js
����m�e� �uІ����d��Q�DOM*��	:���"=�2# ��S�����8š��^o�3J��{kXi �C�sp����m�n��ѱL��E[&�P%<	6MD��C�g�{��
��;Q��iE�su��&�����r����LH�J��П=;�MR?�.#�uQ�S�$�t�DL�Y"�٬�����^�;:�=�\�
����}�)a0��1��!D��0���z��0��K������{["��u�����Ch��.�rx�E�3b���`c��c�7;wh>��6�{� ����V��Q��d2C��)I��������j|3Ȫ���$f�C�c�D�0�*�<^ǔa%�ʒ�y? BX8��6`���E��L7���a�yU��2�l�'!#oL�sI��[y��6 �l]��"={�'��X���JH.ɨ�`�-C:�$y~v1Xo*Y ]�f�Ԕ\�V^���N疊RnM͕�C<�h��|0��/��D�=��E�_�}@~�
0H���Kz��<�x�f��Ug(�]}��,��(��Q]�VôG��:
PmO&�ib����e��x���Ff�o��=�[��B��-�����lp�����{�j@��h��`6UG��+��������k�Ceu�������S�G��WG)"���e��E
w޴.��)����EVp:�"��=�,z�A��� >7��b4�<xs��M�u��4�z�P��H��LL�µlՠ�5�%�)�A/C���#l�ߞ5�2w �S�&�����}c���CtJkG4���}��7>p	�Ԝ2t��� F��6��B���z������}P+��t.m
X����y�ۆ@?��	٦�XzV��D��D��kj�ݯg�-ñ�87�セ��|8 �F�7�!��pZʢ�+�܈�՞/�'ڠ������i��מI=��+r|6|�VH���D��i�^������;�Na���r���?s�Z���/���1R
�b=۩�,?��h��5�"\�2?T���Gо�0W6�, B4�癢S�=�n�˻�0��"p��#�3�-�AAȰv2��Yܼ)�M�+�Q�����<�3��L�0�����^��j�D]������b�QO ;چ��j����z��˷קQ[�+����MM�?�'X�Fhk$��ì]�E��̒�N��\��I��uh�w���<`)&�읓��4(��S��M��>ā��.�e}�ўPt閈�D�Wz��H^Ab%W��� ����/�e�>���UJ�����LE���|����;����5 үr���J�Dk7oH4��zz#k� ���en�
�j���{֟'d�&�gx�W�ѣ�+X��{���򑼺����W��e�����+�ZA�F �+���a٭yCp��@G��$wi�T ��A����?�X�ZO$�q��۳|�v��k�&�,��\ި(L���y��T7��I:V�Sy�*��{
��]�Q�z*�/�(R����g�_�;����g�HI`"N�UVP�
T�d���y�Z�1��fyWA4�٣���	�g��L��Q���߫ͫH���|'D��Ī#�@)
��?���)Q�\r�SJ��z�gc9ܸط��D�܄8���Ƀ����	?�TJ�d�'����C
�p���Y���8G�#�P��BoK�~z����pGn�V����Iq���9r�a}�#��r�?|��$q���̵Ȇ[��CMƎ�sց�/q���B9_���8`{!9���z�c�(A|����m��ͼ�56R��J��C_?�э�>
��{N�Oρ��`�9��`�S)�O��>��������K<\�~�&�� ��ʵG�O�K���Xa< k�����'��C�"F_�^�v���/�;��%�Z��a�š�(��P�`Q�����K]�;�TOǞ_��,���K�������M��mc�yS��'Ü{��5�wڟ�J�����aICş�fP��pAc`�/��`��2����zo��F-����KhP/GK,jt8�6z�qr#�-�S����	E)U�/���B8ܤl^^�e]��vQ���)������mP_�^|��l6,~�%vO��1�\��G<Erqf��S�aX���a�E)�CKGiX3�6*�vw�:F�����4 D���SA�̶0uڐ;Gt���q�QT�UyM��`k�QTSGwp 
�Oa
���ԧ5���
�D�Z+Q:�C��OU �p5+�J�I4Ś{Ӗ�5��+S(�����JT�E�/ �,$&����π4˟	MTF@�fUC���z�r�a�w�~�&<��68��P'qқB|��SF�,ٹd�8�-9�;n._�8���Zk|۟6��l��X_�v>D	Iw#9�3.R��5�z��x"�ToQߚ��l���f��I8u4,��IUa�$�YhoO���*�`r��B��wk�ʉSv>�.���x!�ZhR�\�S��A��:JyW�f�(_b;�����l�=(�]@�B"�b��ͨ�!c�"�6��2�'��_B@Oíf%�����&�е����U*�3R�j�w�o{���������h|;�[��p(�}R���������&/:TN�)�T!F��faж(�a5ۑG�X��"U�j][�?dZ%���xׁ\&mD��m��1�O+�O��4&�p�_D������-��¶6Ge�b�y�R�Հ�FR�/�]��êe�j��rί���i�V ��(�y����^x�Uh��������[gu�����b�OĹXF�����'g����<2�7�/&KF�9�YmK�WT�Æι�ȯ�K ��%!˹�
�n�pJ���&�Bx�m��/λybS6ރhsI1�0���wg��=�e��@�@[=������\��F�e|K�ǫT~NG*͎�i�j�~Y���V jH��L2�'���􃐏�����+ �
�j��E�{U&����M�n��Y�+�t&"	/��3�t:|S��ob�K҉0X8�YD|!���qV�~ĺ�F�qH.�7�t^}�6��V�úf�*kF����+�_5�07��bU��@ڄ�o�DP�C��敜c����5�gȦۊ�g[� ��h ���i���63��/�tDR]T�܌� {�#�����HJn��{��8&f�����d�� w��G����^G���L����I5^zv[��NvA��/^�����~њ�$k�՜��Ϫ�HM��~��8���ww�Ю�?�o��O�W��ܲ�>��뙛�`:L��������̰�Z�(X�[?H�T
��KP�ei��%����b��C4c�'�G���`��Ǽ�����n��+�kz���%\@�Cz}�&�|9�������������H����F�P3�Y]:���3+�Â�Зu*Q�nm�O��,A+���,�M6^���<k��?���V"�W�Ȇ���늠��_2��B��D�侅��:R`�,F��ٗ?���e3Ws=�fazR�R�5�[K�f������?�e7/�Cnx�<8�q�R`a驿�D���{�٨z����H���q�B���2�+�@g�{�:U�JF�!G�QgF�-��n�O�ʺf.�-���	&*�mS̕W7���D�b�a��hۡ�/E�Ě���@I��=?�9�^R!A���5�-mӘb�&����Y��v�C�
�Nb����.�V !@�7��ڔ��rڂ����&��P[֗�u����vA�e_���|��|�	�ۑ#�_��Y�'Uo� �����v�9\F�a�<��;lK]�5����4ev"x���м|�đ�X=�kV�q,R������Bٟ��P���!S�P8��4�	�쉸*=��Q���cq#6���u{~�	=��(���Xq&�TP	�&�ҘA�h��CT�0�ʔj3�p��`f�¬C��'��/|�%��.��MɖzuZ�YM`�v�� ʃV��R
 1�e���)͓��/:n���B�:���!3�,�~��*SO�ǕqK��U�z�1VI����/����
�0��;��{�9!*lX~1���d�|�[2a�O����oyu�Z�_�(��4{�w`�g�.}]��t���/����Y��l�3���+я�W�
7��~)�Ӹˋ�I��?�ڄ�\;�	�,�{�5�B<�G�Z�{�F[���ڥ$*u�UrC��!�xw2D�+LP��	7�cbǕ��5���g����1N���c���t��5����.! (�h��3\##�w�v"��
c _�?�d�Ay���$w,��ip0O��O��@�lR,��0' ����	Ms��X�D�Y�U��'�0k�ñ-�n�'־�BJ#�7MX���D��S�Ax *6G+~%2-�:J�z���>�}^ᤔ40���7������c�C��Hٚ������I��ڎ ��
��
n�����Nk��?��Զ!l��^��W �E��^?���: ��b'����gA�Q���e>�hE[U]owt�wKp����ė^���zS��v}Io�"O���˱���ߞ/sh��zݢ�Hإ%���Ad�?�NJ�4&�R�1�Y��0��7@#�>���[�[ձ#/�{�do�������2�'\�GYv�Ӣv�wc_��vBl�<;^�e�h������Ψ���f�ؗ�R
��z�Z���ϯѿ�)`�{W�Qb�0]��T�w��ؐo�	?�/��bT�B$�1��8�k~0��	���_š�Zb�i���6P1o&�<^6𼏷E'�O� LG�Y��.�8��=tq��8J���
�v�,���6��We�S~	�4�+���c���r׉����qM��Ƹ���3�5x*!�PxHT��z3W���|��)���N��>���a�bơ^�;�(K����z$+Td�!*匆�����n���u2���>D���2�cLB���J!
I����R
���|���N�\�|C�l�|"Bv_q|����c���L��c�|��������Ws!���A�����C[��\�ɠ�&xr�)� ��i�ǿz�����
�'���xI��B��!ڽ�&��I�ۏ*&L��@���eǧ5�z�V�X����hӤ:�t���{�-���3=���MBW	(5#:�{�	��` Y�n�!%U�Ȇ�4�{�]Ku}�f���ݺe�;���>�a��P�{��νlE��+��e{�� �Yz`��{3�����࿩7C�w��"tQ�|a� 1s�Wf02N�!���!)�����p��ֹݾ.wF$o(:�Y��k��	&�09� n��
��u��2��	�|xpf�^s����
w=�dǤ�	-I#������;�[g��3�7�	�¿,2.e�� �D�L��"�S
3��δ�& �jI |��v�S}�>���B���8�^�7]A5Py��n�-gV�/��u�n�"*]F�w��N�VZ:�N4�[ �WOy���M�V���|KlӐ`�����{�ߖ��E���K�pr=K4hHU�mO�?U�c����ܡ����=����l���`�P
��7E:���`��.T���I5�o�j�(��-�����,n�˲[yܽ-"�Mo�b�=�WӞ�,�BX�#�?�ˊ ]69��.�K��G�d����}5Ud8ZL�9�ԝ�́#����ٌ�7q�A������>񕗎_��:ZKdP�N<�e���� a�y���lƓ��m�� &���ޝLAQ���T�J��/�־���g�wqF�$�ҧ�W����> U�F�>���n���Nږ)�E0`.y�X3K`�<�wv�*G�w�0��8a K$�JԾ>~!�(,y�.�#x���big��ʕJ��Ҩ�nvʩ�'A���Gx�7Q���� �]���/�I;�{�߽?<黯P�{֘VV���M�yR~z�gP�d���H_.�8�JP�j��XU�d��Oe�8+�w������q�����v-�y�bB��%'�UD�����n�?Z :8U���!��훖W:��3Ej����6���涠�� � ߴe��}3���y��3ЈA �Hå>�=��,}ΦK<�jb��~B�}Ab����.J�N�V�߀XL��s~\.��τ�͔p�I$�H<����D�/	EP��F�Hux{d��oF�����_���Nt,p����ł&Z�B�j���4YoG�=N��w�	�<KX�1R�8���o)���yc��Ou�^���}�G�$j�Sw��)j��R(�gދ)bE:^�~����EU�Ԓ������R�_V_��:Z�=b8=��v6�?��}�H�-mи��Z��V���=�_o�jU:��.S���J2T
��t)�M�ne���.M��n���6��^��Խ��3�4��e���^ih������ߪ�9��`��RV�!dJQ���F0�������ƛ��]������ ����6V�W���ˡ���G��h�&-fC���f�)�(o�5$������c�,��sy�8�+���m�`������VK�"A�^j���ʅ���%��b��-�v��I�NQ�}�gQ~C%u��w<e�ˁ�	��^�(~A��`#��eY�%�O�W�;�������P^n@�д�HH?p��h����aAc��K�}gKO�{:�[�ןN'oG[I�Ɲ�)���K�4�[���^��I�h�璮�h��B$�7֘���i��I��fÜ8�=E�9L		��C�W����7�j�}�Lr~���?���A�5��|����S�Y7��L[G�)7��Sۮ�HL�}ڙ���d�2�J�k �O"n�Ѿg�LJ_h�y�ɐ"탈��� �_�.^+��h���P�us��5�$Y���B�e��i�V��\���e���)ֺ	a�-��&4c�J��.�����czw@QCm�u�i�%}>�^϶�S�%1e�c�`���]���K�d�d�����ͬ�"��Ղ�����[?�0��vʀ��9��/U�w� �����	�J0�^R[��1��fg<��S8�Ҫ<�a��fz��h"A�0I^khSuc$7;��^����� �E����]�S��~|�5@�w'�h�'��+�����9�����ج�%~�H��Ze34���a�X�����?B�:$i�]�il'��]�:'�I���7al r�A�f�Iq�����m��f�Kֆ�\��d=��Q�Kw��z�	զR�0*m�1xL��'���#�XZA6G&8w,��E�W���`F~�XL����]���h�#���scb��s��9XG�������&�����	�F�a��ۅ��YH��)�L) s��(��g�<oq�Q��H���q���LX�8˱�1�`N�;%� ����Vp��M�gS�]�<�p%�W����3	
�&g:�!�F�$���5O�:���vQjM���{��UX�Fh"�]��<����M0�Ud�&�ՙ�0�?�u��&K۾�����w���,O���)PI,q�Ks0Ej�8ڜ����8�t�I4� ��ې�U�����J�J@+�3Jޅ�y������q�u����DZ(��@�p��3�Kz�#F���')�M�c�` d��FB6؆���!�����⢧�챁�����`]�9<��g}�y|��;ӎ����#R/�]��jU�Exu ��L��Jx����:�i�[І��3���1G$��.�C>X�H�^<��оD���IH�W6���y�K��~�h9W,]k�O�VUS���%���%���7q��A���F)�yʟ2"�[�e����Q�0��K��`��U��"�VӴw=�S?i�	�n��O���D��=پuW]E�V}wm/�cfEI��B�����Y���\���"��n�|z�؀BǓL��e�[�}|A���ACϗ��NU�ռۄƊ]̓��M	��)��[5��F�G8C�6�{�_�Ƹiv��.JuC��ԱP���`�-w���+�q�U*�P���=fI���yee��O_OW��R���a��""5�5��t[mV�7犽?��V�3�����w��#E�`����4��y<�m��k��ٞ����_.��_d$��7L��-h�v=��E�B��X�.K�8${\�IV���=m�t��Ϡ��'o垔BXlb��}%����O���sx8�M�<.��bv�5���7x:�m{�eǬ�b�+� 1�ɥ��%��WQȻ\�|갢"���T�L<�p�vB�S=Q�v°�)����3s@w<o���{��[�']Q3cn.�>Xc�!�CS��v&�;�VÎ_��Ev��VC]�#+9��b�[(DKv����Vn�& *d:��6��&Q�0���V��B\���"v�i.�$YhDl6T5�qU���<W�%%9��\N�����H}| ���9Tb�,S��y �P.8�Nͩķ��9Ss.8��]Y�:\ƜK�:)߸^)JV9���0��Ԛ�>�f&��á�ʺO�T�T�H{b3����S��u�dv
w���ڮn����&���O����!<Qz�ު!T_^|�Sj�rP��)�{��x�JgM��I��e��i0�[�� �Fᾁ� ����7�_*L��m����������h�^>}�**A뀔�d�\,[����ئ<ފ�S�!��S>+p��ï���9⬌_���N�K��~z>j�8,���՜ ��Ί�/t���^�_~�q�u7��9:�%X9�!9�$/��=�����y$�5�<�wu�̭�r�$`���7t�3G�����K(���Gv�1��TY�&���u��y����ȶ}�Fx��>\�M髳g�7rƠ�|bp7��W 3�m��*��h�+`)wO�I�2'���*h�����͊�[x��{�[�n�% 1J�I�J\vƂ�%H$P&�^Dl���]j�|4�ҧ������ʧ~~?�W�AE��1�9c�I�2X�抭=�o���E_{��ұp�c��y=�����Y���u�c�ʍ���B~-ݽ�GyylRM�c�pd[�8;���������	V�#�*,~�Y�������s����P*�k�Q�Uh��r��Pd�D�֘��ޯe�Wb�8!Vh&��Htc���ٴ#�\� �_zg�~�P�$���C�܀�B/	����::(��r:�����B;����wl�yv��vӪ�v�	v����QhP/�v� |���2������	h�i��'e��rm������@<u�b�8\�����*͐�c������K�[z��I�w0�Y�[���o��#�k�4�,��E��g0�oo�}C�#��[')l��\�G��M����"�e��O��i<t�,�ć��EG�M
�S�0.G���Α������I�zO��f2,��R=)AK��g6�.��Mx�B@����cE��j�{ӗ�'�淵s�����S���\5ؒZ�	���������0$�4�DƷv(��+{�����| b��ߨT�7QN�nK���[P��Ml�T1�^�S=�)cR.��AK+�.p�z��*-A7+��b�J;��m��>-0�ۼG�(��	��&���F���h��DbÇ�����&�x7���N��)�4����o�]٭Ew������Kw(��00��>�����K`�4Wo�(��U�si��pI�{D����h���&
FB�M��B���3j��Q�e-��a�?O/�/[x�i$�H"b�@��Z�z��+�EML$�q��l��:��L�6��W��jz�PuS��[\�'�����+ ���%����{JLd˩�ca��;�.�%������A�������E���������jy�ʬ�B��p]�f����:м�Lr�P�H�&@bC����ʇ�{=��Tb��RZb�(s�& �bK��XX<E���5,�< rS��ץ�f���HT��ڷƿ��Ek1Ѐ��JE�j�8X��e2����y�q�h���W�|��umbR��5+��Ga��a��q�+Ĝ�������gU�5o�˷м%�~�jl<��,t,�Sw�[�)q�˹wt诱_�j�1&�|ь��cB
�Ӧ�����J�c3k��i��X�m?�� ���[H!�h7
�Eś�ɜ�5�Q���K367����m�}�² |��//���T*h��V��ْ��>�zIK�)���s���Yl�B�p��$�P�0�wrOP}�	Y,x/|�����[�ɇ0�h��!��E]|����m��2��:�K$K--��ƿ���3��H��q3�ŷe{�K	S@�98�n<Y�:�z���˳2Em�Q��T�N�F�7�1Q�g{��s��-{`}�r��y�}�t���fL�v�S(v���3)��	�^_̃
�����N�\�t&��K��<j�t����,�ѳ���B�e/;9�1��n)�&s�'f�����0D�w
B]?���9uc�/{�H}�nJx�Լ����(�@C��[�@��N[��g�H&V��]�jAZ~�٦�r�|_�T�X�B��kJ��*�M؉Q�,W�o
���b�T	��iLa�ߏÞ������=�e��@�� f��ĨQ/^�?:dU�2���y84�Cn�R� �|J��Mi�\����}
�uNd7�3M
=��Ium|T���t����i���]S)�||�#X�M]J�K�X��^$�I�[�>�n�Z>�띈}
B��|�٣h����|s���mzۈ�h�-b�FKI���y极3Pe��lzE��+��u#ۓ0���ղN���5���(����8�D�C��G�vm-[s{�c���m?��:vY
E*T�]@[ߔi�����zU�=U��� ��'��l2��J��X?4vE
IzP�uW���v̺u<t�8~|ȇ�\��NLĿ�v�ᩛ$�q��t�Q6=��={��c����쎩��8'E�鹮O�+�{�7�����υ���֢�ŏ;�C�2�os+�<G=U@E�Qh���/�������t�r�V}&�V��Y]��x��-���~ ��)�l��+�hWu��R�K�A\�;��JH!�G��(NJ�X�i|���z7cl��\��+��IG�G�%�|���A�%+��A��h�;лfF�^�!��F�.�.���~s����������M�A�GS�m,�"�;_�b����җ�PhĥKr{i�F�$�"���R>F��*G`�˾����e�\E�@e���P��,,M�q��S�i���5����j��e�F�}��3�Ȑ��r������x,A������x>�� ܷ�0�An��a}�L>�hU� ��[4iᦕ���x��iګ�]Bl�@Sf
;� Z��h7�)��EA��p 'ǡ��x~!R��1��Y,�M��ni�K��� �ŉNO؍�o��(��Ї��NO)N��Y�Q���.�zdI藢C4�~^ƺ	��T;��o���u�9A�_���wc���K��&��}�����|\�NG7�y��q�L�D���M�sUY����>��f�ѱȎ°V�����C6�\|r `�����.��w��ۇEuw ]�Я�s&�6$�q��l]�$Ⴅ�PQ[���K႕7ao���{t1 !9�`�2�MS�>kfP��Hf�Ul�^A��;d(0�s�3�$21�ZBpD�b��j˧�7�xs
=���v_�D#o�Kl-����O�%��K��ܓ��R$!��mp|,־�_�4�c�92�U��vH*���ja���[�Jǖ$�c�M</��)sێ�>~_�~�%KKV���*6��`�h��'�i�G����7�^q0々י��D/�u��/V3p}���gj,p��E�\�R4O�&�._�i%�_2zE+�"y4��(���<�!fZ���LP�߃� Y����	�C��v߀��e0*�����������Fݩ?iN{��f>ԃ�J�{^w�C�d�x��#(}��W���T�0Ҍ��g���phee�/
K�';��l
�<���Y��^-�=�3�I�^#��N�q:��0fm|'���?���t�GI��X��Į�K��|u��7��␸~�j�����6��G�t�Ip��/��UOvI�iG9�T3֩�P�u%v����K�����kf����!��P���(d�TY��@�$�Qa� ���m���ɼ#ڢ��������7�裎)��w��u�o\G���u��1�f���ښgsfd��]qQ�:��5I�=����
``����ġ��]t)��	o��K<���&nH� �k��a4�~��;�{���l%�|8v�R�~³�?.^-$p�U8U�[�/��{G�6�~��q����H��T@9�k!�1m��z~�b���%��bqt�C��O���lӺ���.�@�B7U�O��>D27�T�~�ȃ��'͛�g�+��8`�������&^O��R�	�~� �-�ȕn;��$%��%�C�|�\k$~w�n�:��� �v�Ƀ��4�����y�ؘ:7��i��~�*t�UF_Zi'd��]`���	�M(�3��z�$v��*+�'��Ù^���*�QU�»�q%O@�n�|�5gR#�5��3�c>��7Ocʜۦ9��r�ḁ�v�/-69�5J5I�;�4f��~���l�����e��ç�C��nqN��GWק��ro?(�ؒ'J�ۦ�~V1ZĒ)<���J��D^S�ec��]�{��->���G`�Q���l�
u�C�����t�ɴ�l�Qj��CZ�f�Y�p������5�B^�)�hakq,����_��z>W���Q�s'%I}��n<`$�;;3�<���}�f�X�ZU���|��$|�vyb�w�	�"�\��Nb����Z8�2��1i�����jM�	!���8����}s#���b'27h�g� �s��el��y)fI�̌�����2n(������Yv����#r� ��A a+\��L�'����X8n,�<��r�g�TŚ��������;,g/|(p#�<A�}����`��%@��l�"�s�qp���S�e��Uу��I�`^\��s�7��8kܞ8����6��@M8�O�
¸�mϛ{[ґ�MV9��X�n
��޻-����_��
K�C#ڜ�V���'M�F�=���D�b�/[�qB�j���E�^�1�'�I�a��G�}�p_D��u�7P \m���]8���P��.(�ŝ��ln`�(JC��>�x8g5`�����!�?+,���J���٘R!f�yڌ�u���8^R���[j�F��X���V�y<�%x�~��J�y�	���4'�7��Ϣ4S��۹�3Ĺ�ۦ�����Xܬ9pZ��r�1٘�O�^����OZO�o�]�w
`���o��B* G1
�z} ��=f:Y�?4r�'�q��s�� �&������(-�O��m�L�Z�2��ΙH�OV�fI��K��|I3�1aK׍٢w��eJ��3��G��L.����o?�����0x+�:x�{F�5�5���i�����c�"3��Yw�Z��rʟ�)���r�'^�`����,&�C[.]��K�� ��_{��:�:���FK��+�3�h��߈�w
+�s<�]0��X�ڊ4��Sǽ��/�_�����������'�\���܊���d���V=����}��uK	i���
_8;~7��<1��\�Ø9?��9
V��EA�h%hn9���_��@ʿNo�ւ�j��	�u~x���4i�KT�)d�`d_> ��A��t)�q�w�Nh�sx��>ꭷE����e���Ú��!f��p�q-��yE�
����Y'�n>'Y�T�LDt�����]�\��_��nD�wY���c ���f��܎w������P�F�0.���@��r�o��M{2.�������a���G�n7����x�0��B�'߸,T`M�7a��<�O��htE�X�P�<��H��{��5[t�|�<��lh#�g����63��e��ON�B���c��7X�xBT�((ӀT����[A����N��]������T��]�+�Y��R�"R���О1CD.��qb�)z�}��W2:5K	
, ��cA��ͧ���o3/��/��"�]�ѽ�w���t����:~s����)-��Az�w�r�/�`�B�~a4p	1�h{N3l�P���M\�!Z�BP6�u~~��Ǡ��0\��#�,��Z���qi�{�PZ���@sv�����L�ܮ�c��j�I��m���@[o�����n�#c�A�=����XU]���`�-��V�I�l%P������2��W�`��*&�7#�R��yR���?mXG4��t��bZ5`�o�4�sG���z߾^�G�0����f���逶�Ԙ�ex��s���.d9�Uh�4����_2�)to˧:o���7u���lc͍�.�Wmݒ{��O.�F<�(+7W5;�%9ǿ�.,���:}�b�j�Ԛ�d�g� ����g���Z/Z�����gI졳+fi Zr�eK��3�u"�dz�ˁ�;��u)�f��ѭ��U���3 TR\!�Pd�M*��y"��K�u� �ڷݣF�2:�xq!>mI�C���nE��W���-�{�]�W�l���h�2���p�;}|�%�\-b�m
i$r
�^$��I�z��s�G�!����%��Tj��7^��7`�@B�S�4�gǓūW���eĭϚ�we��Վp�칼
y�О�n���L&���D�.
:N"�<a-� 6J�Hs����@26��f��h<���11C�POa���b��fJ�nqg��\����6�o�f��4|0�m��#�#�?� �! ��-L���B��E7zF����,�+(׼,mC66�o0��S��P�5�<D�{0-���4ȫ~8��[H�WVꡈL���:B���qɎl��^��$�V@�)�$���bg�z�R����(����x?�!c(31��+�I̕�"
@�$=Um<�}E�8u%�� ��L�,c,i���bfm��?N������cBi��9|�t����Ph�N��L�3�
U�#��`F�vԀX7<{X��3��y�#^7�xZK��wCg��S�O(����&)X�=R�W��E�G}�l��H���B�͏g�2>��`΂���r�2i��dр����a�0�	]����j�?&u���_�܎���ރ�m�'U�3\U{p�z}�s���6)��?��=�S7kkܛ���@�0�)�_�©�r���zK�V^�����(_D� ��Oݿߋ���<��n���wZخ�Pi��؍Q�Q�w�}�7Ğ_�X�\�dڼ{v� (s�M.}�\��p�8�W �z�
8#��VY
rx�'�63хF�fS�� h��!̉���/�
�hSG����!�&LL3J	��O����9�j�S�;r��o�� �Ҷ.���e|d:JO��z��#\K��t`n��_6.���|Ëj��}���L&�ܐn���Sz�n�&$��y�FD=�����?�o���\ǾW���נ��િR�;~��Bqz�[GD��(<�S�<K44����;QJ~v��z���?eM�6�c����,JH�	v#D�g��nWݭ�2�G��Kn %��)��_����VY�z{�s�]�&��)�}�I�U:uR�:K�O��ߒpm��ޫ#3C��g|g��G)!q����$N������F���(��<�oyʛAC�<�R?3B8h�껿K�%�/�L��5���J�`����5q�;�-z�v���e}�\r�/c�e�>������T��9���7)�&��m�1�r��="�G������d��uR���w������ş���Y�� �Dh)��ho�3?�E�Z86����A�ݤ��_�f��ݽ��,����.�E���>�u�H^�&�#*|�͈>Y��ЁL<�HQhj��K�:20���6@��Sv��oCR|��n���^@�,&���	�͵��(���h(��)BoЊ<'yL��3����Nv&\$�R{�=���ڒ�!=3Rl�Kca��G����Cd"`Iȳ�����Oe_�'Sk�R�r�����d�kyBKe�w������#�=�"�Pgw��0��p^�|�(�ZPϜ�I����bX��C��->��[ ]v��&���]�K�.e�Σ�"����BH�8�o|_Yg�_�.��.�Q��B 9��=�v��ފ�^\�v����R�ۤ�4wV�G��!�B��@F3�+a{���z޺���8��~��zK[�D9*�XX�E@-�TbJ��nb/��r��.�cq��m�9f9���>�O�y9hd��Vm���"pdK��3��K�A������o�rE�q�H��2h�%�r2J=9�2��?O�Ƅ�̂�����z��g�kZX��n��$��h�1'�@�A��fҬj�A�0鼳F'y}��g/�i�*[����ެ�J����A��d���ʑ�w[�;&�2�'W���z�#�V=���$Hb96ڋ�;Nb,6���#<}&���a�XH��~�,�M�!�e�z�z.Ou��@e��D���%5)���n��1�? Ø�Y4�³�E�}n�w�'��@�%��  ��d�~�(Dm�[�Ԩ��K��t��ܾe9�]ų��4�DW�?{�;��lI�D
������
��).ޙU}����&�"5%1�;��eސ�!*���`cx�y�f�G�e�Y�	=ǩK�K�f�.b�$$���	6@kH��/͔�*	8���-�Y�M��_4x:��5a���E��HB��=�$Ͼ����Y�C\I�8�o�=�kk��mz@��iĘax�d������+N��W�����t��ac����i�e�$�8�I�@�������@�p1�	�]��j-���P�Sr��(�s�ů��P6�~��;�ٜ�CF��,"�o3��].1���+��'��`��2��� 7��fŐ�*�5����U��j�\@m4�L	|5����hڀ�m*�S�������_+j��aކ"M<P��`���F;�W��[��A.�����s:Ŧp3"��q$��qdU�0��C�X�Aʦs��ΰ��ew��j�1��Op��&B	J�{j�86����z�crd<M��g]p��vX7wq���Y3�h�"w��#P���l3��-�������]�0ja9��q��!?H��� >ۖ͋<��]���2⦂���.&Pa�D9��@[M�@6���K��;�Ԏ�:�`��Ĳ�X�?'�;��F�����1_VR�ABֿ��� K����>	W)0��td�_y�̙��C��A��)zL���}(4�­T���}�w8�t�К�]>%s�0��@�<.�����rD�,���}I�;��{�������"���y�Wt ���kU�~�Ż�)�2���s�<V������T�s[C�K���埐����o�֚���Q~��y�)���(���ĸ�pg�*�}9Z�D,�c��skV3؈#&D��Y�����v��+��K^�1q��y���O��t��U��z~�)�۶����z��p X�Z'�_Y%�eܮa��/,Fl6�j(����o�eh�/���i7�5N��� ��_/&g���T/ܱ��2�9�8$���Zׄц�Sn��0>IF��v=�s"[�w�b����!r�{>��a�(��Qgf��AX�H~�߫�0:�݂7��Ҿ����3�Q<���G=�P�bލx���9�r٩+	 KmS��p��	![y�R�K�R�SL�zon�ƣ��J��-�uy\�g��v�&aY�q�1|�Gr纲8��h�2k��#�I����:�MN�T�ǌ�Q���-�g�Gy��6V\�x���	�/�.�i<�X� ������H���LЏo��(�ߧP&���3��. �p�9.�62��ﲒl@�R�b!/�
o��W��q�נw������m�uj+�.��s"�ȹGy�x�z���gR������hcxԣ���Сk��t�>b���� Ð�'�#��4�y8��)�W��v�AS�L�@D���,��/�W�A���ؓp����1��[��J�����Z���W(w�@�%�ƴ���J�4��LN��_x�ߩ��n�ίԈ�T�VJ���
u ����ǔ��(�Kw("��&vM�Pq�"Y?7pl4�6m�W@�i�&ww	��'5BvI�xa��vطt�io��$��I�i�W@�g�7�5�pK�/�]s����L+C�/�̏j�5��n�� ��Υ]!�3qp��ֆ
�'=�M�1�ئ'�5 �`��ׅJ���	�\t@9s��n���3>,�C)WQ����Uҏ#�R1�0��>0y�-v�2��"aK���bv�.�\�,�jb[ I�a���{G~]��7��R�2� ��	��W/�<���J�_S�%#]���t��Ӊ;C4��3�Z8��b���ὒ�~ 쀂��F���%�gN��g(��u�d��`�x�}V��ג#�<�ܦ��++dSL��LR<]�n6	n7��>[�AI�g,ؑ�m�پs!�����~D�ek�K1�C)[ɮG��^8I�{-)��>�6�@�Ӽ[5��_��U�����}��[���6}yc$ �s)�ڴZ�s��
�v��tC�k�j��Nd��l�?��H�E
	sK�K��!TK�-�B5@����f����<��(M&>#��� ��Tuġ~�6F�]�Fp��z�~���;�]���1g%��'��'�'vs-�qW��8���N�B�sT��ML)1�+Kh ��v����DW9p�E�Ŷ�(���=�I�lc	"��x�+�Arg���`'��#�|b?Aߚ������Ç�;��59�'ٷ[�!�R�g����.�e��ռw�ĉ�x?���Y�A��7^U&نy�m	9:���()l�h>q$��I�V?a�f�גZ@��~���杊n�����fT�tV�Q�k���I�Cx?�!������j�)
.��q�Y`��s���}��W���+a�A2�,�S�+A.���^�}�Z34�3h�n��`&���O�����e�	XP�Kȃ���$��_Q���j�٩�}Y�k:'�~S򱜎2d���ݝupv�7�q,
� ��{klE~&�B!�2$W6�[�~+���W���!������:ٛ�`���i���O5y�֚��[Q��0�8����<d-+�}Np��^C1L`!���K5eB�J���m�;"�)��v>��4�����ҡtk4/p�~��2�zJ���ӭ4 �I�)$'o������$�B:��ۍ�~��/w|��8"�7 Qx0�v�[*{	���#k¦e��)l5��wm����>.�$��&���h��{(U�gP�D����b1���Gj-�m���N"��zs�>��C���l�C�U��@Z%�)Ӊ32g�#\��*uI������jb�@�'cT;^.��i�T�֯��$AtG���_m�n��8����f5#߱n��z�"�(����{pB�@2�_4m"��8t7��p���,�wr�o�yR E�b,��Q =��?E*�-UY�\�z�"M\�;�i��x�4�����j����{_��Mr���E��^bM��+���w��8�M'3�c��o_�Cv�𝷔���w�����M���/��,�B8���w`G�ˬ#V�f� �o��E�H������[wN���@�1K��M�fyG<���J�QY�=��*�}^���<��LG�)���������;�6���;��m��$S���]f���?���2���%�x���޴�����k�<*{��*zX���P�G�Q�d�=~[�fkNw�S��;a��.�kĻ
�����)����}pp�e����݌��/�� �i�Z@Jyr����j��ێWP��V����Ҥ3#� Y=[$��w��(���A���N`5����$@����.*�5�P���i�FúD�I gXw4� �2�@���0��S�;�BB����7�]l��r�|��5�	�4.�!BZ	!y$c�*�[;8���еy��|1�CY۪F�B
��M��ez���ؤҌ�i���0��tb<�RD�+�{,�_R����yCb����h�'Σ�����K�$�Ȕ (;�)�wٛ[D[#ڳ��=ЃZ�w�7x�Qx(��3�_]����-�0&�X6���p�S�D��W���Ʌ���,�Vt5�p���P�
���-�f���O�5	k�Z��UK�d�~r�����s߉��� �ê�x�J���d����Pc�nOo��%^E�x��V��s���3������#�B�wr����+F������JΓ �s&���0AeR��>�yR0���E�N�r�1]�y�����;T�a~�\��c�p��El��1zƑ�&�oyv��g�u �v��DY%+ob�d���&�W�d�8�h�숟x�mےu�F��X)A�qMΉ�唔�Nn�ׅqr� 
���E�r?�����4
�bA��E�1T�h�FU}] ��y0�
+����/,P���h TN!�p|�|�����3��#�g�JU�L�$
��c����W3g5M�Y�n�@��=���s�ģ�����w�?7���+D#�`
���x7��ݟ�#��Sz�;��`e��7�T��s���@H�Z��r,��,L�m�ic�����EV��8�1�Y�)�itV��G�=o�a+V���H���#��b�X>:r�Ԉ�K��}�&=�NFw\���f���ص�Z6�9���t�!�hy|�6X�˹���*~ލ%DGK������CA��	�� W���3�_\K�9��?�B�}��US���� �����FH���ĸ��fA���i�\ӳ"{Gp��S��\��vqT8�-PP�u�ӌ1�ăDi-z��*.N�+� �Ng��2��X��b��a��_R">2is�6������j6(�X�h0O��S�F(��1�38��D�Ԛ���ȧ	G��פ��0'v��g���j�L�e�#� ���e��El�L|[1�㡂u��I�Kg���a�|õ%����5��V4���^C�l%���0�@(���ޠo��Q�.��5b��X	��oۓ�;0�&����pH6ˌR���К/:�7ɝ��r�;�{��:��Į����0ցw�d+��l�*��l$�1_}�Ya�B4���D�0U�S u�O�S9�F���V�7��R:H��C:�z8d�Ვy�k��%�~<��}�J��fZ������M�6��?���*fQ)h��0Q��{|�b]��Ơ�yT��2A_���*T�Q�r�;5z2	p���|��v���q��ƾr��i���._���H��J��n�ԭ~}8K������RG��w>�M�'����X�7ئ1�6EK[Ey���q;O��,�F��X@�a��^�}�:��F�����Χ�R�e�ǿW�yf���4k r��Ut�'�b��d{y�0R�\W��"��zk �����lg�N���"����k��ˊ��,LK�� h�#1�#$��̵�!�W�L�d�Z�s_��^]�	�R�l��;}���¼����:����W~iz�@���IJ�q�����>���1j"P��*���\�>A������H�C6����H^��If��F}�j
�x,���^��l1u8���qS.�x���S��<�x���(2�h���T{�sV5�8_h��(���^1���W@�����}�?����9�%�=�tJEEn\Fr2	��-��F{9�t_8�d�v���2߰�����wW�CA�%��HY�d�a<D(���0�8֡��C�rO�v5�ˤ�t@Ea�3XI&d�Wד|���E�Pnt�AM9��Hz��8�u�K�d�(�O�6��;��)�si�<6�
-pJ!�[���3
��l�h-=n�S=�y��l<J�����A��Ǉ����FH�F���[�7[���7�&Gb��Q����I���C��"�~m�
�Xe�����n�m]U��T��V�'�Ģ�c��Gmf�=�{�]��8�ނGB�t�� &��ɰ�P
uB
�&��a�<����B�m�KO)2J�\�����2��=z�<��S��oB�U� ��Ea|;�8b�U ���H�d`r��y�L"<����jc蔳@Ryw�vD�cG��� $.2��:�^��;����O�'f!~ :�X���K��O�uU�T�~y%!є�pܽ��Sg��yH������s�W���Cԗ"��3zurv�f�~?�=�ǽ(^ɳ�����33�w������KV�5��,չ��15����!o�Bx(�i��Yc�,��*`�a�h"Qm�ʧ����zJK���s�M�H���0�'�)������3�O�$ɴ��Γ���4)	!�7����m��b�Eq��.Pw�"׶���� (3��{�L�W|���/G�Lq�Nͮ��R8��;��e��o�p�O�������:Ѹ���ƒ�;f�iU	r��W�{8�9aV�	�����9m��2>�&����0�e Ą����L��k�pA�����a��\��NFs�=P`@2^������1j����:��_bN�+ M��	q<�T��&��}�"EB�����'+�s�Pu3�6J�/|���i� w��Lh�F�&���� .��k���l�K`�D7�Ȥ�9٫|]QO��+7��N��Nx��e�	L�K�vir8S���A�8n�ި~�)��^�q��"�g �D���'�F��-��O�/�m�C����,T�훋ǘj�a�21�*?��2|m��a��]:**�1X!������)U�%z��&�c:juL+<1���ǯ�PvO��!���~��u�3�?���˱P4������f(����s:v������wr���;�F�ÓVZ�A�5��eKۇ�̉f��^�.P+�N�6y�WZ��}q�.���T��C�(�wL\�Z�����/_ Ais�d���ˮ�̂(ZI/�N�);��E���(�� ��\϶�M�����vB�Y@�؝L��c�Apg�*C׉�M?�ay��"%�t�d���Q��n��m'|O�rd��nKd}.�Ҁ�ݘ��a���q����/�W&�8o�YN���2���+N�<n��h�쀠��Ӫ��guD%����:_�<�q@�y����:zmm�*�వݗa�Qvg�&�J�i(� oǏ������@�z�|k������G��;ק"\T\����\8���9BC�WV���p�3��~*��?��^4OZ�̺�N�	�Nn6�g���8�P����%n�� �k�D�A�ںU�D�:f-�y�=J������s^�(�<�u�&F6��4h�d�:d);�=b���>0��jMJ�,2��<嚤�\����t*��N--��li
� �Oۜ��lT0��B���0�*�.BWR��ܡ���`�А�]�-�^�sE������~�)'<�iE�j��0
隝���\r����+����3Q������]�7J�r���vB���x�����)�G����㨹K7�Sǂ��/e1��˗��Z���"�4�K�����'2ZR�+
��i�Æwpt� ��X�$���; Pu�*�fvf_k�m��#@�o ;��5��������I�Crʤ���Qf�� �҇,�Z�CS7L�W�!��l�ZIO��V�������k��?6,԰*�	�.9�ƾX9�(��'�(S#�� ��*�*~RTAu�(w���0�/��y6��*8�'�t�uK@`��'o�VO���@-0l%�ђ?bH�E<5Ƒ��	ᰬ��I.�Ez� �1�|@۠5��vx\�wF8ќబSM5���3A)�/�R�dp].,;�P;�B�,n��G�U<�RN��iI!N]J{����E����a��Vxq�����/�k����D�M,�RY�sd�>���xD��ӵaўC�10c���)�ǅ÷���W{FT{A�y��ڽ1!ge\zK�����u�ha.��KS�k��/+�&&�E�0��Rg9��e��k�����j�G�5���^x7'|�-��Ñ��UR���J������e�c���w�d�*�?����7^�:�� =@������[��tE���7@1P�R�����ꊸO/=�6O�aۿR-�@���"r�S�ˮ�-��-�,4ɧ(흤����:s���+�^**�:xe��,K��و��e}=��G�mYC�ek TM(S���f0F�o<>E�i��?���n��K�urR�J��X;�m������w3���pQl~B���W�1��)�g%����/�rF�Je��)�e�{������$����9q����A�w�#GM1���}�ڔ��p�Y�B
	��D����9+sT�Nl�7�F�+�?3���s��Į�k��-�]P(-EfrIr��ZY��5�W�m��_�4�?��3�O�Db�.�ot��ɜ��LlH%��2R'Mr:j�Xf��p���{V5У�,�@�O�@c�[��;f���4>�`{T_�q���� ���|Zd��PS�V����(}5�Ȥg��cV���8����I�4���2PF��R�-
�_hW�^y����=�Q�ӽ��8Wj�rd_r�؛����I�T.+�e}�k��.��,��뵩��3�­����!Y��dL����w�ҷ�l&��hw$�����3�p�T�A�)�����;o��l���7�ʩ��J4A���K����V��Ե��Z�М���A-Cx~��&�m�v����Uo�@?�ќ�6���s���b ^�!�~" ї��B��?\<��g���˯t�ŕ��/t�S�@5��E��%���^@ �
�Y�E� ����)�#Y�K!�h5N�ïU�P����HO.-��dg�cЊ���j}�aaux��[��$�6�>^F����]~(=ߎ1N�xT4�(��|�
t}�M��S��&j��B���M��MM�(Q$����m�C������ˏ'�8��������Y���VG#d��F��Tx���
u�Ӝ*�Ӭ��5��~ER��=����8�k��!�'�'�X֏��
��sPEW�T�S�*S�+��i�H����-s0|�������x�I�c��Ui"�
�Z��p��C��?-t�����dh�?g���_�mr����Z|�ҽL��P����7�X�Q���O�;{�p���l�Z�9o�s�z�ו���#{F&����R��\�+���s�j��sS�;+:�