��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|����z=+���v�����p��6f�z�3��w��g��ķ�H7P�\Νg*�.�%F>�vg�Ԣ`͙Қ�y��&�L<��Đm}x��(�di��N'�K�π�wգ&��ݎ�30,pŉ�$[�1�5� ��_.G/4�w ��Yʖ���(�E�T�OH��cN�{�:sT������mi^Q�oϲd�,��}7#�lUh��L�T,u0���T��ԐJ���H*�u���5��)r�7��/��ܵ�A��h�Ul���Aï�z�ȵ���h�հY�i3q����(-!C�k�|ʿ��C,D��yW��+z� ��)���
O� >�9��o�o����mD��"{�5y|�Y�ҡrx�.��Nd ��  Bݠ|��F���\d^Y<�W~�>��|?�QN���lLЃ�����潑 �W2ϔ�^�L������S%�@��oٶ���R� ���'�_v�V��	Q�[?����t�̙�
wA<���r8lߎ��s�U�ޤ#�t��.�|嬿L����BӀ���!l歭�%.��j�e)X�-!͏P�j[;г�FNS��٘��S�)�4*�P�h)�˥��$��!4�4�7{�k��=}N|"�����ʧ��W''_z��� ��ʆч;ʍL��jJg�$y[��E�^�S�p���F���SY{�4U��y7�֭.�xH�=Pd��z�����B�g���B,��?@9՞���13,�wQ�V�����&�������v���\ �+fKG�i$���d�ꜘ����ʅ<8�J�?���=��6�Mk�&4�l6�P�`�;c�SG�۩�h��:PIRn�a�N��a0KS����R>��]yZ'�s.�(�@�z$�&�� y�/����EM�-�"�W<h"2r?n�1�$bL�kP���*�����k�V]�n��%�籕A9��v�y�Yi8�ʙVۓ�ݔÍ���-�x>i�S�^_��4{�լ������r���;�N�g#$p01箈ΰ������
/YS��@bۈ����u0WOꌓM�"�
�e2N4l��ItF�����d��#h�a�m�m�lL��ҾOg��:�\\��2ϱH��+�@�� �HN@i��5�Uȧ���J��p�}p�A��P�:ac�+oE����`���x/	��SV	�L��GH��`��5i`�h��Gt����o{t�)�i԰�}��ۈo���,�"�
?n�.C�-��^F�4*��՟T��h�V�\k���j��y_�#Tۧ�Ne�L�TZq;���D�9���u~��X��2�G�9,���O�\�O�l&	�<6�Uj�m�p,-$3P�R��;�D!׼�/�j�A��N��U5B��������e� ������aK�)�Z&-�dJT����=�c�[3&�m��^�Bk��L��������tO��
�Ĉl���Ũ)z�|�E����Hg�R(���w�
�ǫ�3�;���e����btu���p�������>��t�=�n���^ݏe����I��)l�C��ذቺ�]/}X�O�O���J��WJ��L��@$���t�}.@.Zg�1*b����L`� �̊� �7|yx�BAK�/p9�N�L�'������5�޷�`:��a����@G�	yyΟ?�>�r?,�8˗�S��p���:�I�sSj�J
 �5=d[�=���^�G�U������L-���vQZ[h���y�_�K@֖�7w)6$�0,G�� 8�'�̤3֚���(�w������_�O�'�a۞}g��m�
�z�t_ ��Y�����&r,�GBl�����*��X���L�����Ј9�хJc�S��!�3���8w���< ���	����=�
)�) �؄&S��9b^@ ��`��Y��M2w�Ne��P�"r{�G��CmO�BL������M7N����~����}���1���B���7�o��b�;�����;ʾ�7X0s���fx���
�n���J^O���ͬ�����_I�^LP:p�KG�+0:� ��0��F@�E�6��D��!eZ�S��a���zN/)p7�c��E�;�؟�3��ukn��`'g�+�Q8���s�6d���=�}}�2������d ap��0}=�p�̜]Q�,@q��gq�|�?�i�#{A�M������ ����(3�Mv�t]=/��/>�r+y���$8
ic�E�e9����E�%�z(��@_�M�	\���Bϭ�t�F�K�*x����� ծ�#�SV��<	h>�S� �I���5܇���4)(�e�xb�w:�h5_apy��B
4��f7�>��=:2x����*�;��m*�۳2�C?�df�<��7q�����(�.�G�>	G�7�by������Z�Fk��N�}6�j#����e8����䑝�K�<,�^M�ʿ���c柿��ƴ#�7�)	d_%\::�JT�.������DC tVr�(化'A��+u1m�H+aM�`v��ÖǝHo_Aw* ��w��P�P��@�T��\���]��g��ç'k�!�q��y��Q�������Z%O��a��$���=(�� ��Y�R?"V���=���ҳ���-S�0ɾ8�C:�\ߒT.�bIh��-G%��Y�c��g]�j�Pw��Ǳ�w�R�01cb�vP��Z.������,�=�E��P���f��p���7�s@���R%��``J�@a6@8�ܜ��Q��i�������"4Un{@c�~o"J�G�� �����!�o�� �:SBq<���d˪�)���B�o��B�$������е@+c��j�Қ�����v�e�+;b,̠��<PY���nemG`�9������i� '��U(Y:�k"YJ"+��_�'r<�'�l�G�}��U��2&81K�cE�bH������Qӏ�� .B �w��CTV��9
�Χ��'�NVW����1Pɤ�>��z��E������|����I�B�n�����S�j;2`qO����W���:Ƈ��w���!��Ƀ�:�.Rm�O�˝�Cl��~�'iFP/�^H�*��g;f|��T�
c������O�m)� �*j�b�3���ѽM���,�9<��[Ԡ��K��0�H�Ba_0fl�ƻzs�,�E���
t�d��@8�� �G�"?l��Goj^I�7�c}(�exdn+"��ڌm(�@�1��\z�f[�I �;�s�F�,��H����}>��ͣ���ڞ�8��FY2���~�vY�a�mX���B�a�c���Ɓ�#)n����m���^�B2UE$����(M#+�?�쿒l�}�
�Q���t��8���C���o���c��(Z������ ��"��\򟶺6X����^o�Y82��}�a�Ee(
�����qi�\
��\>vfT�F��{nV��{,�9&��Y�[�F�ʒ�DKEu|@i�cTc���x/�x\�gۃC�3��&OO���PW�^�Mm�clτjSˢ�nWW�-��9??���|T��o��a��k�XH��E-7���Q���F�ܨjMe�2�G�d�p���:yȅ�P�^��}x����