��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� f
���O�Q��Y.#�d'���J�"����4���d�"�Ŝ9͜����
�~�a�rN�����o]y����1���nJ�]s 3L!��,���zَaw�{,���{�b�[;ҙ�u�\��������.7���}����H��ΰ�&���ے9��y��y����͍2��ё(��7q|U9��1���i��$>�[�G���^#fU����S�"_a[7B��7~ez�#�5��-������>[{Љ�v��G]��Ew4��5`�|x}��4�y�z�f�|#�դ�e��5p���1��L��d=�㺔��y���h����V���Q���t�̿�rբ��6�j�mcP�iT
���c�j��5�j�KL��tlV��d��x�Z��"ks�kCK�|�i(�;�����6��12�XTeP��[��'�0u ����r/X�<��/�]Gȥ���%N��]84����Uwp)
���un(c�Åf��J��f`9Fqv]���+�<�w �N��fѧ�h ˞�C;4��#�i��T6n�Q�T�����ڸ}�rS3�*�x�٨�j���y�~E�s�~+s�G��'��%`+�w+.}��(Jľ�$SL�2-�M�M�W5~���/%��t%���0;��3��G�rq�Ħ@];
!}ˬ � C_3ZjT5�ъ���29L��>ԡ��I�#iDn=*oB'R�؍����v��< 2<���oc�M Yx�R5��ܡ�����2=ړU��oLW9oq��4S�um줂f�X+��t)�a��� R��M�Ć8��,=���LIQN��wJ��̩��O{Bi`g�.�c����6T8���u�������_=�����L�+�����{\5d?D�_&��Ju)��R�$���R�⡔���7L��"�PM�\��DRR�0/���j��H�z�H��?jiٵ��W=1�!��ep|ۿj�Cm=�]��Mlb$z��ł6T�M�����n*�����u������Ⱦ�qG���r�x�f�&l�)K�?ft65�X�!G��m�^[y-,�� pv�R(ݵ\H��^p=����	ß��P�6~�	N Xfy%X���*9Ψ�sn���3��P?0� ��L�?���Q!9bR�
T�z�$�z��,�����C�U�3��ö}�?v�7CRL�|��C�&J;wZ{K���ӕ�̩Fv�0w�I��X�F�D��ZY��ѹ�v��b�f_���u�"_���`�`9g��'MZ+�9:��yZT�(�P�bKNK�T�Ɛ�ZGd�V+n��?_b`D�#t5��~�O|<�C���}�ǁ\9���`p����C���ky���fi�_��©�Ȓ�_��{�t�a,�/�9��B����F��D�u��.��@h�[��֬�0n�ε��;�n��O��{s�[����o����V4v��f�� �/L�D9g��w�l �����7�w68�����	º9+�����|�g1 �mi*�Sa$�P*>u�h'�c������s�
-������k�"���Rϯ7��Ј�Q�����{F�3�L;�
����km'ѓ����r&R7w� Qz-����ډ7;p�]�}���'1I�`wo�2��'.6�39�����z��	J�����k)��N&Щ�m���j��J����wO���ˀ�9TKs��%��9b�2�4>1��v����=�%T\��E'@�~��]s ��1s�������&�f�ڋ�
��3��{�8���	7I��-�!��&w��R�@�
�U�)���Z~B�
��9xXX��o��#��x@���q��(�L���$�j�[��ݷ�[�"0+M�-����h�nք!Yۖw'��� ���-U����Hh�Sr�"c�tC'>�z|S7�Y�\.`|�3�m�En�᭭Gobu�XSWVS��c$i��dR;��t�;Y)�@�"+:v������l��4����~�إ�P���T�A4��W�)"��$O����|5s."N|;��AJdQ�U��>��>��MG�w�\A;��A������AD�O�ٔ�2Q�vU��g7�8LĲ^l�v:K�t�o����s���.ˑ)����-O�q����ܭ y��F���=���x�x�N��4L�z�Z�W5�h��3Q�ޝo��7����	��+��|���z�o���D�	fo��;�`b|/�l-�����#��=�癘�撱���E�T�{@����r��{v��_ą{`���f�W���{�8�-�Ezu�ި/��.�X����`�H�ꖐ�
k";�X�3���#�)����H��F������r�z7�p%�h�O=�s�2��� ���l���)|p(<$Mw������ȷ�y���E�S�&��8�������U��w����6����
�z��Ӟ% h�B�늑"�2fWH�0Y-�!����;V�ц���3:�}�^�\�����$º�-l�)J~9dr���LH�3ɐ��������heG^9:�U���OJ!K�0[W@�ܠ b�K�(�h���7��񁣁 �PZ<q���1=���>f��ڪtT�˼A�S_ ��rCU*�6d��&�zP�Dd0�|&2`�]�Uˏ�;�T���16����t���X��d�B�/}���(�_�RQ�F�b �u4AY֡��6%�H̉-�y��尨�<�O��+�:7��dS�?�&`�v	IǠ	�����X;�m1ɯ�L�CF2������1d���<|᷃��.�?P����*�ri�%���I|�����Yu�ѳY���4�mSŸ�,j&����:���b��쵅���Βz���jB�J�^��?��u�r���&�+^�3�z�{
��c�qnVFgW�o��ֱ
�(|u[B�M�c��jf��|�TK7�W[]��r��A!AP�����}�by��y�{���U\� դB˺��T�'﮵@�BL��(���$L湑:�~{��jd�w��@-:i�;4��i�'��u�s�*�2����0[��?�z��g���HR6��nI��VZ��!�3����og,.�q�߱��
�Χ̹B���
���4