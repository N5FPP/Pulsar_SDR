��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY�Ɗ�����5����� ��o���*����	���b�Q��'���Z��߰N�
�t��ߌl���U z�9����Þ�%|Nؚ�*�N.��F�+��)�YvnX����\v�S�]���	mKi����@�
�V}�Mv�lwj�Z�6O{9L����ǚq�?0O�9#����憸�H��\M����6-�4���L!/(8{r��9��1�f��5	��-$���N�	�f�H��uرmɤ��Y�K�Z��K��Rb�)�}V:�2�\J��>�j,�6���=�M�q #� &<p�mS*c�,]��W���DV��?�#E�b6�d���Zn���Tᑩ~tw����pI����(R�_�X��51nD�nψ>-w6�fs�ʍ�RZ�==�#�p3����&���l�[�mM0���1`~��p�����@S+;&V�隣�����)�/a�kp@�+:�<U��t(>x٢.�u ����H(��N�>:�]9x��QZ� W1�0�VB��25��/*��9q�t�𧌌"��_^q�+᭨<<"C�����&�G�����k��*	�.{v�6p��c�	��E4}[��#��D��a���+���ֶ9X3qųI��)	�4Pw��׏�ԅ�AI7�}��W`���&8��#A.`��۞�'���2t�%��Qz��0݁ �Ryo,!����9��e7��7a�B(z� ]��>ZX#�s`�ou�k3L�lg�s���q�C�_Ѫ��K�da��>x!��h�O|:Vc�i ��lhƲ�⮼궈tE�D]XX��)��EW�-������C����ͳϫ ���n�`(�C��o����%� �$5^��j��ng���U�yT9Y���o#��1��岤��ݷͿ�㽾, ���]v��A0�ÃjJ�j�@�a?M��]x�d�VCu��>�ĥO�ب)u�;����֟��G"%17�IkC-zx��[��+u�B2���y��K؞F'��_u���))9�U���=�C�
{@��C4В&�%c��P�n�e���]pا�������۳�h�3����}�+�HxUBe2������Q-�cZ7/zi.�I�O8E��]vu�;��ŒߧZb�ZU�0*ݏ6{�ж���W�״ץ�b>��#��Ƽ	,��Һ�Ų����G+{U,B�MW
��#x����M���m����,�iM+"#,���+�D1o&�۱gd�"V=�ȗ*��Y��W�h���5k޺?�RǺf�%͌R] ��R�?���2��_�ьCeNqll�kT�,����c}����;0M��ȃP�" X�(�b$"�RmI
��[���p%����"~�yX`�;�g2�h)���'��jVc
W`:��#@�9��l��J�D�p돢�SKث��o$]������?1�]|�����!t��s�����.�v@cR�{S^
@���(DKN�#4���?�"�,���G��ߡ��
��J<iЀsK��=����͢�f�J��E��Ǖ�R������dP��(�����.�� �0
�e�����{b�4��<�8�s�j��5Ww$aӸM D��A9&+@<12z�6m͚��X6<�,C߮�P��Y����31��V��!�����Э�f7�DmB{��q��@�v� �%�M7z���H�1�G����x.k���ύ� �;KQ����"ĳ�ً\��Z��b++������>��p�|�De�����B���X�g3�����N�~Z�+[��D�EJM���g�ʶ��
^�v�w1-�ۡaQ�j��,]������:�LM��_/Pq@T�\7�@�U�f$�(2}_�5>��ݗYX�Ih+�Y(Jj��Hnͅ-�����g{+uR�H;|��>y#�/T�h��Bڦx���N��_�M�«{�7�ݵ�����0����cG���ʨE�}�:��.���W������i5B�����=Y�^��)��$[��LXЩ��=��o�x��1�FԐ.�N����G��ӎy�*�D�i]C�~	�m��$��u­��,`͞�"c>�9��oLx(,U&��A�?�4����	�P^u�Y;� .�����oGN5�KL�����Cf�z[�����BT���5�ĳ�ݗ	)aW-9ٰ���f�'�b�$����pt.�y=��!���a���S����*.Rx�?�:�a�-�ϗrm����u{W3HA��N��:��/z]�}�y>'�����(�[�|�̔��A0	�q��^[!����4�׳4�q)�[�>c��-��R�u�����Dj�M�4�{Pn�V\�(������"���D�߯���c���8�����֞gB������+�?��κ�$%����O!q�Ʉf�6e�F����~��jkE s�@Zـ�昼�g��o��ώ�]XĈ��?n�5�b����A�(�H<2=yc��t(�j��\S;�0�=4��;㇙{��P &��������lh l�@ ��� W�1ג�'D�9�"�����=
иk��M8d�}��\�E����Ӛ�cm�=���VH��K�	���67w{R��aS�#���M�3�gOǷ�'��&�z�zT@�**�/��R5����H���c�)`O����Kv���d�����"���x���U�7���c��u��h��T��qX��4��a
�޺2�c��<��.�At)��KŐ��B`�Z[@��ê�5���͓ ��y����O-G=@�9P(ݯ�5�|ڋ4�u�A7�"[	l��q��T݃�!��d
����=�Ph�vg�����O0�8B6�]���[z"�}�t?q+��
�5�i$��Đ�4�c��jc���4�E���Ȋ����3�xE�;Y�/��(mZAq:˼��}�Q�lX8�����p��5�x@إ�}��������2�o�{S�"��x�T�X�=�s��wӍ��I�*9yH�^�sf6'�my�Qt?{����.�Oor�ַUkh�Mb�>	���k�uG����?���,��&q�5�z{���9��M�V���� z7U1��� �۠x� �����m�zfmNL�N�@2x9帞��4X{���.��� P��5$�;	�p̯Ѷ� �� �5�㳯�l�3�If��F.�R�\�Hu}�Ɨ�z�S �W�����)m=���Ʈƅ0�x�{�@_RSf���^q��_HWP ������ĨU+^M�/�D��x��$طo���^jdB4�9z�v4�o���p0�;����slGX#��%�
L��݅v�L�������U�+�M��L<�����R�b� t"\�� �
,�G}���kh2����_��U��������C��^gn<#��^�A����AF)�~ 1M�u�1�>����a�~���`n��
 �ُ�S��X��z5aK��o�B�P���"�g�4����-�r���4f�r�ZCOK�O�-M���������2	F����8�������Q�9�R~�ZS��yBP���f��n�NqW6�I��+Suy��]����/酤�T ^�F�x>)*���W�N6=����C��l����*h}�:a_ ��:�p��"	�{�P.�n]�{'���U ���GR����
��G�qcIjK�"�e��]橐�pBK1k�>�BxUY�羿�E2=������ $�r�Co��G3����F �������n]�B=�h%k��ưk�
�kL~����]'�tS孁k�Ĵhi�Ʌ��B�60�!��B4�>ٸ��Q���u@J&骕�4�`&��{;��X�l�jSgZ>��.�Vs���vg+��ȅI��HR{���ꏻ����3�7��RQ�+�:(�[�[�~'��Q��F�H�1�ߘ��[���T��d��=m�wW��{!����<r���LG8�R<�Fƶ��F�t?����-���Ės4S�Z� O �v�!;�/E���-oB��@cK0�w&yd'[�bM�����.��!��놶��4p��a��a�/��9Jt�����{g�T�]��<��D��
}�}�f\����R��Q��&�W�ٙ�]���"��_HM�����w� ��\�T	�L5�7�T�l�k|ϙ:)���&Oޢv<�z���+�](}� r�v����7J�Fbeg~��TH 
?{%�澒�8�@��](������"�� }�������������Q��!�Lb�PԱYoz��&S�R�N�]#Yu�{Xg��AN� ���Z�<d��!(�����*���j�AD[�ٮ}���*<��=j��t���p��鬢��7�w�(ӯn����0<��R:���ts�[%юZM���@�g:H����*~U}ܦN�0XYmF�n�b�+����z�wWP�?	t�1������{�B��_��� �C	�����kȁ;u�քI��XVe�H{U��D~��t��B�ɠ���|��+�� h�m#����?�~$��޸�Oa��v��)�j��-�#N������<�;#��\Bg��ہ���(�Z���������^��Z�NY�{XE�j��Q�f-����1v���@�&����E2E?���l<���v7�t�}G'ګ��Շd�)>v0��(:�}�CF(L���	6iH�ޟ�o�}��^f�^qYέ���R��1�$kg��)L��l��re%C�t��w|2~7V*W�-������Y��ٟjD�$����|�G���Bֳ՞��s��@Efǃm�1��,�Y?˚���瘫݈W�<��H���q\'Hx���V��Ʒ\�0q�D�ǋc��~m�J��U9�NRXS�CJ������4Ъ��hO�P�)Е��B�TaXY]��z빠�-��2�E>H�d����8�R���A�v�gp�tMʟY�6]Bģ��	�S����{.7�*�u�Z��OH�����$��V�8�O9ͻq����9$��Zz	"�}(l�?��se�Ŧ�h�:%z�8?�1�����H���+��*��9�j��>��>'�X�n��@YH���c{�\<��K���C½<�bc;F����6'T�	ؒjĄ�>v����4�)f!�g�W��; ���̨�@ev����6��{ŋ��ow�e���\���;R�3��#pC��Ie��5�&K%{�O�K�Q�d&��
��1cs�Gw�LZ�ƥ�;2w���M��4��/�FD�5��O�߷*��"P�I�k���.��+��GAt,O���2?@�}�y>­�g�K��1/��������ꃌMl�v:�!:l��&j׼
�ln5T$.�p|ű,	�ڴ8�8Y�?i7���!
(#끎���t��w�"�OZ�� �P���#�i�ނąbM���b��0k����Ck�[rF�R�� n�;��"U��-��P!�,"
(�	�z��s����*�7>s߾~��>�'���~�C% ��]\x�i!!�76N�p�y�/�#�ͯFs�
�d.��ԛ}�	�cm~Ap6@uC�vjl��I�&�QU24W���Ÿe���`b6}�z��k!1'C�oɛ�ФY��=b5����u��0�荶�G_�*}�(G��3�F��5�W�{��d���� ��?������t�J}3�{�3�Kz��l_`x�⩩�BxZ[��/P��ʊ���w��@LZ�GJ��N~�dN�3I�S[;Rd��f+��.�k�G��:Z�us��;?~��$�o�r�K��fr�;�	����i�.iVX����Xh"��R�ܽ,Gؿ�Y˚*m,9O�{�b���?��83���]�C��/�"���g�4�Т�j���!��-,���9_fYܞ����ՏB]u
�k�@n���@:��L�f�eJ�X���S�f�0b�m��Vx�2�@��$�b�M��֯Ĵ���j'��	�k5�e�<R�a:5�y�4�~��_���4m�WI�oB�W�0#�'�GAPWR9�GK����Ȉ���|��>�O�<�el��L_�y8㻕�i��0��s�3![:����b3��r�|�z��������@j�^`�SDZ�T9B# �� v뭐��%��CDp�����9�F)n���MU��;��-�v�B�I��8�D��u��=��"�F�v޻A��v!r^������hp�={�$,�t^�)�@�r4��%�_�9/ܱ���{^H�}6�l
�`��^B�לa*�˄XY�a�C�֞�u���t"ď�~�����l9�Vr�ۦ��ۛ�}uA�gf�L�^]�B�RLW�^�5�d>Ӟ"��0�Ɗ�-�;���A�$�f_�x<ӑ�{�=6�a��P��V��jЭTYj�����PӴ�����f������LS�M��6�~���¦]�Q�p�k-��Vry���إ�t�s�_k���WL�)��E�kG����(#��I�sZ����Ǖ��&����n\#����D�+����f�S�,��G��g�&ҧ_%[�An���AU���� �(�Ljm��ڼ���-�\�))�8Q��KX�����!�4-���MFB�9�Ķ�ԭƜ-����BCBU�����T��ZB�m�|Tg.%BZ�r¼]>\���Hx�5��c�����k�-L_X�G��e��}ْ�Ҷ�f�����FS�Q6b�@�{%rʿU�[߱.�.�W��ŧ��)�	�6��*j��+����u��%&L����`�*�]v�YsxD�g�p�Od`ph�5|ָ/G�Zykα��'w��β���������bޫ�2�,�"?f^�.�
�¹nT�C�M^�ENztC8/m��tw��&6/VΨ��+k��^���my#����Կj���!�բ�ze�{4�<r^��r���HJ�O�jw��6��Ib#d��D�4���j����lR֣v�����.�z�^rwU&�5��`�Q#ov�=X5���H
A�J�(�X���uY<�M	Y]�6�D�X�(��l,�R���p×��6|CA����ԝ����{�W/�
7 �R>5>`���,�LQ>l���}l�3ɬ�f��)x��E� 0�r��*iт��R�����:_`���CN���B%y7�����1d4��`2����_�����4IO���C��K)�D�<���N�2������x�+��^n��cͺ�X�A**��5A���� v��
�n,�T`08�6���"��µ-QvňSv)\k���]��էh��w�L� .�x��� x	����{@�Mbo�����De�0�`�ULCT����cEx�hέ,ۛ���A��;g.d��.���B��.�Y�amِ�X�q�z+_�Yǚ~����,:0�"���v�d��X��a��'�@[�X������Q�ʕ������KT�aD{Z�\uY���iģ�UCv��^`�?��ߜ^�};e\	e�s�;���'��D�F����R�^�����˘~~��ɓn{��xx��\5B���ln�5�5[|򜈪�
�M|��jV��n���n��i"�[Q��V��X����ɽ�����#��6�*m*�1�j*B�t!�>u?�1���ʵ^��}G
��M����|~Rr����WW(�Ui�-�7���*�o�3�����;E���Kd�hV>&�1�q繊2	�������n� ��y���I��IZl�,.E0��Q��屑�(O�嗕Ɉ2 u�ǼB��a����j����M����ф6%���P�^����m��+0�"$X�k2LR*l���C�����L�L�����mQ��;��4�T{�V ���6V��]~�7�=,2m�p��;W��b�'r�_C�Tbo3�����T�}t��]_�ͬ�|'_��<a�#�GRi�f��9~�2���l�?�/�iDЉJ�Ejt�͵�6[�J{wǟ;��Y��ڄD�2��W�x���U��pxu@����v	Jml��
�-�b�`�l]v�s�o�O.5ؑK�#\sfp����}D�iج��������c���iƍm����=b�����]Y��9ģ��7������,��N��f��б֛C��, �A��ܡ�|��d��b[5�Z��cz��K��x�0 B�QIn��|��&���å��*;��.�)'�X�aotw�n�w=�	���k���)��`�&U
\ �����,���▚#��3D�5��|�G�/y{B��PBP ��`���#X1�� �$2C�Т�;����I��]�}�aޢ�V��{.�j%ճ����.1�ɓ��Ė����Y��V�|rw�6�5��<���T�6XW�!���˪���E�_��d�y���$zX)��Џm����<���7̳-C����B�<1g$H�=QÕ
�$7���M,��'�����$X� �y�HHM)�O������"�lm�̩��b_�hZ b�͠�1��i�R��i�?�;��q�؄�~b��z�ʆ�H�k\�)��l�h��n;6E�tD�[y�;�TlT:�F.�e�MS�G���k�7A������&��Mn���2	�cӖ@��D6dȳ�5��.�da�a���ފ�z��6�ps�, :,����������*ʅ�ow��1���R�s��e4y���y��h���3'�p�|�9�m-q����ڔ����nF�Kp`�rQ��p���1L +�'Щ�{�DC"*�M%�r-�x2�e��vC\X����Sx9���H)3<2QT�6�~#��M#SL%��P���0?�����_s.���m��{Kh��t$���w�S[��ى�A���xן�:���C<W�\���.�z�)�B���#�m������;�>A������)=e:j+��Ϙ�P��^i�h/u�6���Hq�b�c4�G�2�$�'�6�hr
![�}��N��Wؘ�7�<}N���rV ��A�G��l���bz��<���g�ۉ�%Ħ�<E,P���ؤާ�8K>>B����i�l$�Ň �8��*�-��1�������{^�kz��}ƣ��x����
EBCQ�;�X��8A�S%u�ZgK�k ,O� dv��$�r���8
��_-��_R��e��E3���������-��ѹs����P�*^=��5.���n\5_��b�Yh�-������ߠ����7�W�f^,�qoq"�T2Њ�G-�$���[p1(����xt;eVzě��m�bzآ<=��],{�U��I�l1j%�S�َ��hv���m�_w�y��$���J9ݭ�O� kΦ��{럶�79ȫq���ݤ��ՇI
ge�Lufݖ�~���)n�3��bD�2�6�JLg���ڡQ�oc����Z�j�`Sރ��q�+}��-��x��.���}e��A�&�-�5l�)!F|�l͜��d����#��靄�x>�OR����+C��Ƃ�W�7��V���e՗Õ�}m����;r*B��.olXT����0��:h��	��T�ʴ�O��\>����*fE7�y�jH=��"�
[���18�� r:G�|�@��=���I���N/r�B�fE��7�bH��&m?)�&�!�߬��8��O ��,�X�gf/qd.	�M2��Bm�)�_\Ŧ ��N(�#Q�M�^�A��_t �㜯jB��y3dϻ<B�����CQ�� �C]���x����fb��ڧޓ�����y�!��<����T���_��Q��r[�������@���Ӈz��!�p_?��!����b�|,�Km�	{5�y�
\%�:Cd��/���5������&�,��+���V����/�cIw�:R�:#�3���O'7>�����r��>��Ѽ���ĈDŅ�(�Č�.o����ٝ���Ÿ4�9o;$�8
d�9. �L���u?xҗ��"UeNxp��
�Ffm�:|�R�5��7	Q��͋��[T�>��2�G��@�bv�$S�Otn�҇��
�����z����:�:�t�x_�C:�s���Բ�&�V���چ��X�/f�"��f���+bE9џ���������i�ED䇈ί��IC�u�6ov�3���ndA88x��/+̀�4)UB�bu:�g��]T��)3������z�0,g,�1/ 5$[�k�'��DP~�t���M��z�E-�6;>�6�K�}��A��d��e���dt�u��=5E�Y���N�y?���pO�|Y,��*Y�Z�B��ш|I����}��Z��9���F뀮�=�P�[y����yY�3�
�!��k�2;2%uw��3 1�U����kcz\h���j��X06Q���rK�fML����z�������\2l�!��to���,Gvf�u�_��H[�ͧi�_�!��#>|�YE�;z�*�m�"0����W���V�.
0�#fI��PQ'�=�y�bR\�ʵ�<��#��R���1�Ӕ:Pr���a"At�nFۂb�`w�ر�!�u�M<j�
x��	]T�}�/�7�j�v:��?� Y��A4WO�=��)�Yx�RQi��D�H�<���OV�$��,��Q�!�H����?�$��O /�	�~�K�C+NY��>�^�ƅ�l��1�N@�J��)�6�����ӊ�uD��X4w���w��#$�<�*��k�I6!��f�'%��o�;)
��p���yh������7pd'�nn����A��y��ľh�yM=���K�bR�F������пH�=�&}"/Ȩ���้0��R��Vvdj�&���q������m��(���/ �x�Ű��d����KL5�������	�'Qn�GQ�yHc�=9HZQ����8��	��j�Q�J�Υ�5a&q��ueDlDd����k��N㭯���"V+��I�M� gJ�Q�pR��^�V�XE�� ��ʿjbV��a	^w��p��8^w�_[������tdv��%�ڳƬ�@vF"&���#&D7/�ê�(g�!�n��E������L�����ǹx��Q��x���g܆	�[��X�]3�����h��4֔;�ߧ��q���Ⱦ]��A�������'��暿g���cqύ�ݜ�t��?z$m�L���D�ϩp&�'ۥ$�X���=�rH1�8��Eb�T��M�����;��u4��0��ߪu�5{iН���8��`�ﴄv_�cS���^�C���/L�V-4�D��TJa[������*�J��=�*�L��_`94!��B���j������j[z���n�O����b�[��% 9�e����"b�F突%�$3��v
cq� 15@hļ���Mų�4IO-�$�X�.�����Ǵ&:jN���'
Ue��L��#�A<G,6!��і�?�W�o��.�v%B	+���~�����:�a���ai-;L��"�(���/���LփԨ�:b�|kj��;.R�ɔpR���Ynb�>r�F�c$ @Nt#�w�iڄp�D��ؒuS�4����ݥ�WS Q ��.Q����⢣�-v��~�0�!��z�𻭗\dZ������&��C<|����{b%���W�l�ͣ�߾E�����+z�0�9p���sՈ�N�gO�|��#�0�R7G�R�4)���qA��A�ap�}���&{��Y� �-�D0#��nP�4Z�ĥ����7&��z2�Jx�}�x~������{̯�)@�ue�C�g4�B����m�RoY>z�w�I��h��^�}��Q�,�Gh�H���d�J�_�9q��#�-��|��Њ�vl��O��KBӌ5e�e6�������ɪnv�iȊ�Mq��`�L.�����$z�����,�|�j��T�r��ɮ��V?�AZƘE^����(�q�3����gb��o�P�jcY��y2�Qs;QB�!4�B��@�?���V��i������NS�Ǿу0sC5����pwoe��|/i��؁���e���]�i��wݭ���f`~G԰{Z��'^I�[��O�)�7E��s�ƨ��f���O�*�Zm&:<��`�<4ΐ)0~ �1���˷`nk_Hn;_�B����qR�5W�)���6�+PA�� p�
E�����s=7�P���H s?J\E'7��\A�Z2���	]�-�D`^Oa�ǈAз)�2�iP�	qNz��]=̚@����J�q����?��Q���u�dT(`Xs��-��Z�4?�.��|� �C���qxf�2sy��j��*�]�TF/��r%�(�GJkeNx��Bc�K"��.U�ٕ�s�5��G���������! ��gE._����Nr��sR"?v$��ԭ���e��A'I�0n��'�pw&��� ����>̚J��!�����&���[~��o:4R��Un������RfeDѬ���TWo�R�~]2%��U�"��M��'�x��e�>uT��df���Փ�����l�RS;'e	\3cc��1�,�]B���i�{��[8�P���_�ʊ�e+ݮ��Av�%�_ �X(��#i�)���8�<��ʢ�6u�	 ѕY�bи��	$[ŸU1ybjO���<�M��eA�9��O�"S�Sz߰>�j�:4���h��@�euB�E��0V�C'�CULj���o�d#��^ș�ʜ���~uyo
�_��D�"Ͱ0�a�E{���c7��o�֗I^��نg!�Ep�܏8�m�N�H���*ė�?Orz�.l�(P�;�;���D�D21�ۉKb+	�l{,F�T7�u���g��KKD>5��?כ��������oH��<A�$�a��X1�4^��<]�i)eub=0���ʄyd�]�3��'��:T��=v\��7�V6��2|'O�mQ��FUc���E���ߍ����i�M��쑕��ެ����Ճ%6��9� ��%5C�Hr�υ�M��:�/,�m=҄BO��p��\�n� ���6���wAS2�z�o>��E�ZDi��H�@<��f��+���Ni_�D1#jc����|�-^�B,�t�/6�6:l��E^�����=���禶���=��/M;�g�m�(��{�>� �F"&$Qr��qL����iAO����0@ܬ4���ZU���$��ij��>|�}\��8I�g�H��e!U�6] <��,�|꾊�g\� _��!p"R�S)��<���d[����)F�� cS�����)^<ƗI2���P�%������ G�7*4~}0N�QĀ�r��C��c{�����q[����PO�#_���P}��y6Ĵ�m��Pl�e@$e�6���	 ���E�oՉTRu�[�gȆT$�6Es�:h dFBX]P�ʝ?�\���9!� $�޹YYW���'��	]�h�~����߸S������E��䮟�K��H���FR۳��YF0#,�����1d �y�L�=Aq���'�(�,��3�p�J�k�D}Ϭ_ݫ�T��A�)?�!��A���P��np �̉-O�7�,Ibߓ�����r��%m�b�Ɔ�~5u�*��P�: �
*����&�r%�0�+�[�KKퟐgXɂ��RR\����6�,����G,<-���i�b���a�L�?��@L�����CX�i�X��eE�~߂
ZAg�Onp��
�D���0ߧLo���A���{�B�4V���}��(�d�eqB*p*�"�Iwτ�PM�b���F�1!��@J���ܖt�ʦ��a�[�F��f�H�@0�K���Cg:��;�� !`�撑�~�����}h}!K:�;'N>1�7�!QKS�x����l�5������Pc[s��:�b}�)$����mw�M�}��zE{��b��(
��;l���yR���?�?G�h�:m%\�!��8��	�t��84�o��+C�b�2�7+��ֳ}טz�Ɏ�p)�Ց��N��6�\-�z�a���HK?;�rVPcu�h~@㯀��I�XD� ��-L~Yςi;<�,<K���Z����ծ��5}8��קܠV��w2$�Á�3�4l��2�������\	hc�Ҡ%?߷Lfgڑ��8���|H�[�N)(��K���:�U�k5f��4C?t~T׈�c��j-iҶ�߃Bu����l}������J뿴x=��j( Ď�~�_U_�՜
x���P��D�k��g4�:F�V��~Y�N�Xt��	�une�I�Yr�U�>}�`�L�� ��k,��B���n+؎�U�&O,k/�����D�O-���]1�m� ��hsV�pa�p����<*J��=U��~^I�}8��M�Jp���C_�uLm��'ݖ�+Ǡ�3���ƣ��A�I��$����V��o5F{3�W�M�s����9���hX�UEe���*s�&i�ctdP���J~�	B˒yޙr�'s��djrƝ=<#3oX�PC\آ�/"�Ü�~�el""�����E״(t��R1�S�=M���&�XZ�f�Z���?�����]�#�Ս�M�^o
=9�(�$��EvZ�vs����,p��mߍh+
�tN����mq�M��L�W|G8�"r�H���Y+�����1���/�Z-�RKr$M� O��z�`�K�Q�B�I�*�0��Â�[c�I�O�<��+�}��lp|�j�p���0>׀x>s�N&�������b=�L��k�@�	v�%"F���F�񤣣պcX�J3��*<Y���,�z�nH�!�.�`y
�ia��������6�]�Z��t��hv_���̥P��.AR���3��aeH�F��$��)j،S-��V��B��>�	�=|���[��SO���ZQT�%D���&bvX#��neR�`-��{�v#ǃ�`�I�s�Y�@w-�P�ͪ7?_�W�7�I���_@~I���?Lt a�m�Y{�1åtT-jx��u�|q1P O������f��ǅH�,�ʚ�"�Vfv�;��&C��MR��p�+D��-��ĩP�>51��m즚�t �{`#lٗ��ߢ�C�%p[�E��$`u�f2R�ȁ�m�ȏ�)&�+deFb�5i��PI.�6�Z��]���I�Q��?��;V�$��[^T�)I�7���G\��קQ� ZW��I����������"ƛth�E���k�A���QG��D�5�	����'ޢt�Y0:���.)��N��u$}�R"�Gه֖�H����~�4�V-�I�w� �lN���Z+s�9SQ��C͸������F���&������:�7�O��ώ�w�yĭ����Ql�H��̰Lÿ{;��� z�ϛG$���^&c=Z���{HÜೲ���8�OF���Z"^�i����WS � R��Ι�D�)^�)�=�A�ʅa�s�I<~�Ӌ�N�yL�E�r������44�i��}����i@�pLL��0��e����R��{ԋӂ)�l�Kir�&.iq���Kwω.:5'�yV�����Ր[��X�y΁|�Y��T`��0��i9���w�����
���J�y5_u�(R�y3�P��� �B���ǀZ�L^r�{X(x�d���Ņ�2�56ݏ��F�Là���I�=!N�1���OF�O��r@4l%;��DQ�S���[��~�k?~M�t)�0��%��i�����E��>���Hx�+,(8�r�#/��I[���)�np��X�-WH��C{����Pǵ�~=3~6E$+C��vR�Ν��=u�~�TUT:��Q�[�B��C�Q2o7C�#<�����AS�?��� 5x.�N,��a[M-^�7�_���BC��C�F��ɔ�sO���Mt!����_�Y�6�7=�\�1����#	ڹ�t9dWF8Z�X����nTc��Ƚiօ:ɺ��#P��5��ˤ)H���e�D�{˵R�U���֙݋����Ӧ�g�9���a:L��:n�0��h]��cL$�q����7�T,����&��xFpu�1��_QAV'����iQ��#OĲ��+��W�������{�dUg�k�#���:��D�D��X�L�8xvOo%G�sS�k�PZk��,opkθT�_��f;�~�N&� �W~�.:�� �er���v���Jq�!鳓q��I§�p���""Ӿ�<<_QG�vR�\�*u��(�</�G�N�V�g���@]�<A������T��}�@LGwE��=�]�s7��
�<�˃x�d+�S�Bq75��uk;u�3E斊�P6$'�F?���������[e�4B;����p6޿�NU����so��*[e�ȟ
�����0��+EMℿ������<�H�&�ֹ�̗�[�}#m���y������d[��f�BΙ�&$���}>�/��siH(��8��Ƨ�����t��A����8�3�=�:"z��~�i�i	�3J�E�2���W���1-g���y�����ﲃ,�T�$e��NJ����6i�N�"��Y�E�vw����~�)A���F &Y��P��"R����\�N�hbqv�Eo�m����Rf*2��7����3|��H��Q�����K�����N�g
V�@��0y1�R�_���V	��Շᓲ�^�*Ϳ�@��ཽ��������%̸�T�:�P�"|���
f+�m���^W�W��{����+�E���67 t����Y�-������1n��,�ӛ≽:�!V 7j�ٯ��"��g�r��<y�&Q0M�qAy�h��T��Y�PAz��;�N��U����:}��>5�j,�k.�	�9:�����*RV�
�4j���_v�2�E!!H�Ǽ��g�ȧ6IS�N��S�t%�߼�Ӝ\g\&T�WZI�m�������F�����h�I�J�@t�J�	�'�	�Z�i��g��V��n_��+2B�Uu�����~�%i{�R4b�/�<UF@l��ř���~:�i���n��(��c݀�H�OF8'oe��]P������mO�=��WO�|�]�}�8K�2D�?D��{��	�S ���%�AԶז�V^�lX��9��U�˯&��?m�������է�]����[Kj�sa��#8R�z�^G^�i5��`�ENY�1b����vDZsXJ'��=�KP�+W�	�z_)�b����Ӈ�;�d�ѯW�$� �R�0�޵�Y���V�KE�'~�������e2��3�`�a$n�"�0���.��}N��Z�F%#��7�)���<3o�B��T�܇���v�}�PDt�̙֩��D�c����w���e�LO��d^C�߫ ���w�{�n�ǚ����o庪ʬ}��_�z5g�� Q�ac�y���i������Ev�L�I.	�ll8��qܜ.��>��\�_��<�Z��m���������r�Ϙ\�l��,u+��]CQ�v��ƈC�a��,���n�)Q�oBp��vnl��ح�q�V�A2�|�g�$:�R������G�j��Qn<ͼ������A�g�hYL�������M�H�4��.WM<�lD�FE��"�T c����L�Z�#�=&N�Kr�IgM��0{����m��85�@�Qk�4?��G���a��@��cI��t�ÓGs���HFA�P�~�K}#H�k�>�^&���|W�I�kx�$s��Ȕ@9�'h<�MY�OJ��ݷ�J	[T�K�E�d�re���������V���4{q+V�oUvr%r�.�O����������z|��y���V��i��\�U`)Y�I0����k�^�"�n?���ށg��_��ʤL�ARU�McB��]~�tE9�ح伮����X�z�s�-����h�D�x����c.�t?�j�B����a�����,��'|$h��g �aR�lA�;�>��JO��se�E����&U��������]�F�)�L�HX�v~�(бt�55 C�����:m�a��+�B@��瑽��Gy^���A^h0��
Ȁ'�?sPr4.�%b��ߋo �8Q%M=ȴT�.+"�Va� 6 Z[� ,���UDl% ��ڣM����u&\0E����`�]��nt�ibT��"�zu�xq��ǿ?ZK���:Dz�edo�+�e].�*6s˽
��6x��P?1��$�쬥\i	���c�igL4E���^���G%��s�ʔ�-ӵ2=�k�?w�r�ѴԺ%�	���rQ~w��x]h���p�ZVB���Y�Ad
����4 ���r+�<#�}�\�����BZJj�����isyDY�q���w��h���!��m`#˝�x�}��F�'���#�P��ަ���x�V"��|!�O��_��d��1@ӕ��$q%�N���E�׋m��t2D��g��3	�I�s�bM��#�3�YN��aO���ެLlz2�xB	AB��]x廉���/�*&�@��#i�d.0-27{W��H~q̀6�E;_q˪�3	�LB4����&"w'��&�x�w���u%b^��r�&�� �q�X�	1lK&5���#6a��߻�1��Tt�;�FIĩg/B������fe��Kq���Sʿ��r+BZ���pI�F^	ۏ�l����.u���!	��x�AO���1��x,�̵�̭C��$¤�=�m.@)���V�%��j�Z_�JzKȁ��A�~J`����W�5lx]+Ύ�U����cs�0tZa9���m�P���o�VRI|�0kQ�a��FaL(�Lq��]����Xk2�pf�
���ׯ��&�?>��;��f���4w	R�8����AI/A-��ZI��C�d��c�w
�G�祧�*Wz ���Y}������E��s�fR�zI�Ͷ<��{��et��v�Х+�ԟ���H����g�y�)�߄QD)�Z�`�q�_/����HZ�+i���N�c��@w
�Ͻ�$C�Pq������T�PP빊�?�>V�o :@�a�q@�����z�&�� ~Ų�1x �r��T�N�pR{�7l[�L��җ�G�rzVԁt'J�!�gG~F�~�h܇�q��T��@?|k�m|�{rݜգ��a7��	W#���z�ˈ@\x�1��i�$�M+1i�7�d�E�;h�S�kPV�}B�<e�n�;ǲ���Hg�q"*�� �^��Jմ�.3 _���`��q���Jay��@�0�pp��ؙ����:6�T��K#�f�=��/#�e���T�(w�,[J���v��̀�"�È`����$*5�� �|�V�M�pS�!���08�+�6��U� ��1����'D�,���d�N5�:���}����	�	��Q-�wx�Vl�)���s|�0��W�X� ��L��\�Ή����)')#��L���fE��H�tp��ڟ�d�Q��P'$3���P,�(�������#o�p�kP����e��r�C�����F6�t.�0KK.�?nԠ	� ��Ѩ��:[S���5"�f��"rZ��sR��mj�D_+�ir}P5��W|� ����Q"<u�ZZ���4`ȵ��8~����2$}�v~���W'2�Q�b�R����W˾��͇�����ރ,��ɛn���A�{ _s��O����ŵR*�8|a�9n�v����S'aS|Π݀�*�[ov���$�md�8ή�Xcd� :���wt8+�0X����K ����a��6���&`���8r�}��V�1	�����b1�$}{�=i��)�6
������@�D|��*?�vS���q�q��w�����^tI�TJ��4c��Ҫ�"e�ڱד��I	�O�Y 	_���u5u>��2ސq���};������xi��^r8�<_Y��IW�}��"�޾��5�ǲ��ӺE_�j��r�^ރ����� �v����y'�$!�U��UO��co6�OZ����cd����%%�5��2��M�ʮ�Cv�\~7���V��k�4���-� u�C�E`geC��6r_S�M�~(�;o3z�}��)��`V�I��7�]d�i�)�8�Q*g���rр<�Q|�CZ�Y����R�M"[ ��i���rx�ឺoH�Z��;��-���B�s����D�_��<�6��%��1L0֎�E��/Ғ��,�Ii��`A��`�XX���(�pϐ��-m��'�G��;�����u�w|
��c��y��ϯ�����o�%AlR%��]�ʲd��Z��hi�0�?t�y���|��F =6D�RVqx����M����.=|�|�R�H�6�9�C���A?G⧄�2`$��Sr]Z��u���tM���:P0sƌ�����P#3��?�s������ڷv�/���ۆ��� Q���� �kYK���I���<Q�b�L=��*Jd��3\G�T�E�����1r�D���`�*�|V+4(�p~��'ݜ$�������ތ�H��P��Ց���Vɗ:�:O7�+��O�l�"!A-��HwJ�r�E?Ox�wBS�1ð�X�|�t�.��ՉN��r�T,�w3����ܸ�K��Vl����G �-��}���7�~�d�=%I)%�8m�t�����.�V�`���(����9��¯sw��K��&�;�_�џ�����=��ڂ��w��Yb�OJ�?���ݓ2��g�l��vD��	9��*_���[h��5�i�
�^gQL���- �@Ի?@G��%gf�7R[�{C� t�}�ؙ�����D\E)��?׍����X��Pf&������W� ��>} �v5�e8C�b&*��tt�zTǠ������<�j,�!Ub��&�y������%�l'�֌,������/j�$O�N[`57�4�e������NYq�rd78@㉁��!Vk� |�\۩��f䐹v�+b��y�k$�A�^c��Uֿ�a����4>� �'OH7��ل-U��q�
*���>�2��^B��E���EJz踻2ļ4�/OD��7���hO$ ��l�5�/�=���<ԃR��Ӱ��'����xg�ǈ�2��m����/�D;�����ـ.�>�g�;&��h�f���{nyݥ35�{�Gp(6!��)-�F�O%K�0��:$N����]�5h/���`U�0`��2�o��*T��O㍐�ӗ=D��4�����;S��<?L�;�i�X�`tՖ�*i�U]n�]*�7�;�F�F$y�|���V��7_�B�aQ�X+d31i�D`�thBS
��E�>_H�g2����D�>D�Q!��#��t�g:��{��Y���L������\Z>S���ő�<it� �&���<n/��|��,U07�m�|G/�������6�(�B�_��㊦��{��;�n�FKa_�a��L�)\�j+{�9yQ�!�X����z������i����Cy�%���h�o�rR�!�N})#�}p�	۱��#�z�#�o`��\���)e% �)ߡ�
�O���è;�������������c_�:]>
8��+p;�:�T]�r�٠�94Ąw`4�J����P�ȷ��D&�F���o�?���[�'Zڞ�r~CY�$<�f�tu�J�z�#�����b��Ǟ�ؗ��a�m!��9�? �b��A��be��>Q�l���B�cv<$+��wy������c ݋*,R��ʍ߿)N���jsHQ�֔dt�S��З�r:�H�wU�v�\����4;.�N�^�$�}��g&^��Ia�#5!���e{Qг�.2N�$����wYҭ��{�� 
d����o㊿��l��,����m(�̜����nل�1�񣬓�8`^�]s�ʦ �x�
&:�E��./U�$���|P`�Fpز��?���W"�9�lta�R�O٘��Rٶ�Z�57g�BR  �z����LӮ�#�r�8p�Ư�H^|�Z'qk���=oƟPK����Q��E�w��#Sv����@H��k��D���������$!��|&��J ����K��c��)3Y=����ѳ���V���H+�mPt�����b,�����&M�,�F����;P�-]/Ae<��f��H%v�k.�!R��'�R�"i9d�k*sһ�,&5��"��PP�Iu�RQvx$4����L�Z��X�|R���fmO��W�TF�2�-g���g�ۑ����:u�7͍���v�(�fLZ�C�?E�cM{/�����[�=���oi��nAL�������ALk�X��qܑ���2��޼���z0�ZҀb�ҹ	5`���4y*�L4��Nc�$L:�]�,*��]� ���+���~�6�O��
�P��қ�)�H�������)�����r��^����.�^��"V�n���yQ.��4��x@�7hxTIv30���<��K*H8����Up)�R\�f<�`�%#�e��݅�!G�]dc�AJ���]��y�P+����S_�u?����Cx=�WܶB;��pN��J�ykƧ1	�8��4�ڴ��)Ca}3�]L���=�X����%��͡�rc��;5����k=m���_��]�T�ԟ�X�+mYQ�qJ~!7��9��L:c�-�V%�RkQ���ںy9$�p���|E0花���8��a�`]���0c��Z%���L�Z`�O!	�~3�.�.s�-Z;0��H
;��i,r��1Z~��BՂ� ��\�!��s�C	|.�l꧉��M�K\V鲒���;�d����^�b1�)M4?�S$�LϮ�]o�.���c�K�TU�'�q�mk�;���|F�8n>NmԄ l{�JG	ZU����>�M�+��0�&k�|,�H�(&Mn~ڻU��B�ؾ�upx*[��"x��X�:��Y=C��ա;�0ˀ����*=��c�=w�M��$��݁�JY.��ȕPڸ��s���$,�'Bm�-���A��aɫ��\H��_u�M����s�`)T/9��lx�yѻУ!����7αX'���� Cm���^��O�U�7��GcJt�C�d�Bc=�W���o�q4e8�c�q?d�"�jVw�M�i�ѧo�v���S'���Vk�G�(Z*�X�489�8�O�I�s$<���?tr�Z�^4��>*t�pP�4���P�\��6�Fo����\��6�B|+p����9�m���V��6߫r�����z�^T���tA�X�<X�����U��e�sZ|��}g1a?|[Z��Fu�u?̱f/hnr�[5#hų�i2ܥ4�9=���EU�vqPRP��)��Mw�Dym7�Oh�-���v�����O���$��\���n]�T���6��WD�J�6�e�8zs�D�\}n�{�e]��6E�9�z�Xi�⫢]����ͤ�Y5��bO�T �o۶��ZX�= ��Y!1�V��G���7챗a���GZ�,-H�
_CB��(8y���lmyrUKo�t�Y� 0 ��nq��Q���GOI ᇤs���(���heO�����H������6����-���Jv���9i�#t���܈JNzu2�c��׺�?[�a�Fؾ���D1���V�%��PW�sW��F��E$R+������?D�k��Z�`���D�5�y�3G��mƬ�Zb�R����`�bG����ƹ m�o~:�9�\_G�f{1G�@1>�6 Bcq�}s�E1����_�S#/�.l�ђ�Q�|�T��8d��2wnr@4��e��K ɤ�Ep��b���0��?[��M��9�k���N�JW�K��d��S�B.�R]H��)��0��I�.�"9G��#����7(6Z���:D���������#�鐽��ݏ=��	&{�T��f�WO����0��$�J22���P;lU.jBq"���m'e��Y>i|�k <��jƤ��<��ge؊��c��}2ͩSH�̒IrC,�:f�?Ѣ-څ����׊(�D �\�+�5��i�Q5[�	Q#Ϟ^>ݯ�Ny�Ӹ�$�`̄Qn��X�PO�b!bc��X3����I��uQD^s��N���`g����A��lw�)�
�u�,��.u�hN���B?fPtr��c��{O~nu67WH|�Dߞ�O���/��(�|<�=;H��>�,c�MK+��V˸�rpp�XC=x�?ʆ�L�l����%�SZ>�?�_}I�,J�!��k*o�$8k�����l� BJ�J�8�j����7:����o�r�yD�d��O@�c�0-*]��5�_s4���=�t��A'X��ED��jQ� ��Bo[_ƃ���^\;�Þ��c]?ԥԁ��Z��K%�$����7���ґpe��#�,����k��[ ����!h��Ҹ9�#�A>�w��I'w%�����X����orcӕ���|-%#4���0����3� ���	�.e�-���&�����z�u��_f¢���>g�Y,|J*	���KGh)���ގ@�t�}�u���&�r�p��Mkޚ�f`�mo�YS��,/K���]��p��|q=J�Lag�d��s��_y_xWi!���%�<��^��

!� \^� ��?^Ȥ�A��$y)��xu('���OrF��_�e�T!�C��,�T�~v�DZ������"��	���q'b����m�3�&=0���(mi"�T�۝���>����'w=�(\'E�/B��?2�P�����c^�N�BL�	��6��|���][w]����!X�����2�2�;��0 b���pFFE�"���5�W,�5�#�Ui����F�n�$���}��
��M.U���ي]��8k��qY��E`�V+Y"�V��V9Z��:�ͫ��|&=�42��׀7FS�x�ɾ�u�`42f��u/$�����;�2�7L?P����Hj�C��d�wN�~u}
��A��.wS���2�y̮�r#��xr���?��/��/~���HHy�[K���B!nx��Ҁ���=��_ֳ��$/&(KL�?��G�ۓ�c�;��ޒ��eڋ%(;	�0YM��;�p
A��� "�֨:��X��+g���u�K��BpA�6��qJAkd��O:��;HKƥZ%0O뗈�L�6�pؿ��J"�u�(�lt�l�<�5U�J#�MV��ftS�ôg��܉5�[�N�?�2�C�R��.�+�J'#���O,���C��K�Zg���=ۛ�EA�T��I���s�,�2#�[n�1a��̖��b;ʔ�0���h�(��/`1��TYE#hb�߂�B�6�>7�Cotz��<�4y�瀡�ٓbo�i�tB?�}Fk�Sj�J����>��_&��Rsu��5[����"�pJ��̋�?�LL��hQ�}h�s/H��� }��1�0G!O��
��ᆨ�(LW����`�~9�*�� j��m��c��t���مA�h���S&��h=�WaϜ���4�o�b��~�+�"��\f1�BRV�����$e-�`�A�V����P�V��C� ��P#�9��5w�l�넳
@��ࡪ��Q�`�q8|�%��Cc�!�����e��\���U��}��_��B�U����� �w,Q�w ��u��L���NR����Ա/v\aaP��&Vɶ�A���,5c���n� )���OD�H����Ac7G[PB
���b_�R�T���"�$�W���m�e*ZD���;�Y��f[<�x�C���I�x2�Ji�7s�K����+\��`ڋ�`?^b�y76ם��Hw�H���֐:e�u�.����%��B:��P5D�d��xk�V܂����N��M$����a��Tn����̚�bZ,��TI4i0��T�KOQ���9�uB��8�`���]Ʀ8�s\<?1G�!�����C�mIl��."#�낻oZ]��Úw'�w�����\�ȯf�e��z�c��̧�i���@'�G5X1�7ѭjOv�����`e4�/}xIy+���x��P��{'�[LΨ>6�?��,r7ǲgV�wH͟yi=Q�^*���Y1��D
w����g'� �t4�ju�F�0�M����L�qH��$�����4�����n"��`�����M���xxw@�vբ%����FeMr������7~�G9��=��+y$kBvn��5n]Ri�fg{�;U������x�J��mm��їH��B�5tU1I.Ep��N��+���æ�`.�������h,���m(;_�tP�\Aճ=ԖӾ4�y\J~2����
X(W�~qj
C�3ѱx^����<�R�$��2���x�N�F���D�	�>�J�sQ���g�t��b�w�I9W[Ɗo����aSEo�x��3��)��l���> ��L�3�~(A��7P�zY���*�J�⫃.\��A�!���yF3�N�o?�<
i�$̋��P�B�u������1(}�0�<&+�!D���HGВ�DW�������b��#��u�f���E�z&��2������U��G�F�ұ�.daR�.��6Id@���)�MԊ�͠Xޕ�o=�9"h�*ʸ��7���AD��a������U��?/����N�!�W�ޖ��}��TS(��9���n��3.(���z����~."0��5Q�I+�x�[�z[Ll��[�c�V�3ҁ�&$mߙ� U��a����S�"5E�j�����Ȑ;{T��\�4�6Zaԧ�mtw��O�낼��5��K@�l=���\Q4A
��A��H*hҩ]�s����W�z��B]�dn���n*n�8����$�D�!�܌" ]��za��!bH悍�w5R�ZQ�6�;q�[��aX�|�nG���T�J��T�ۤ���ޅ=s�Gg@�!l�i�#�Ż���iẞ�x+IoSY�K�"�l�������7��.��C(�>roZ���'�)��Y��.��U	]\�"=�;���Z�"t�U2l��:$���������"�?�τ@�q���C	kR(��w���!�~M�Ɲ�i��s�d�p� �{��;#�P�ZMR���w��PDⶼ�^L�Kr6��xVm���)�R��G.�S���]B:�B�Ukȫ�y�m�8��A�U/�ƭ����&�>K���A���ޭ�e����%�A� �8;�R�{�����&��`.)c�_p���W痹��@?�a���Q� �<��J	f~����0mQ��!�x��euq��%�3%����ݷDB�hb�ڞs��dFiW����c
�4~�N1��!�+n�<����+&�t�3���RL�:y��i��}t�d_t;x� ���I��-� �q�P(^��(a�Q�� �?��ڼՌ&�9Kϡ(�1�z�f��F���ɫI���@��f��3�$�q��ݜ>���}0���W{i��7���;tm��Q��}o���/�/��nC� ]�ucX�H%��ag:�Y���~��"/ba�Kw�TB��ky����Rn���9Z��\٩DDT�ZH��|��k��Fy:�i�nB��|��S\�;����³�z���nP2,H@,3�y3��!3z�6�i��P
b-"I �Jt�'k#��5�����N;����Rɹ #A��{r^��N�?�\H2��c*��fD��7Os��!���?�������ۨ0s��(���.�4���?��������Ȣ��SY��<��o�{n㝜 ,�X�����TX����e�-{��l�{)��P��%�Y&S1���N_@.�d`��2܋{0�t0~��/{N��{��!+h��I4ͦ��$l5�����x�~��|�n=ST�mFB���]�ͷ�!XN�Z�>�m^Q!E�]�}P6"v��N�={�t�I�2�gD5�������qJ~�Ξ ddV�!�3D�N��� �j`z�RN�O9�(��U}i|�z�J�҄T8�}7?-<��1�K���G��A�W?u�����@�N�	)��4��15c����ꨙL`��TAKYcR�Vz�y�)�F&����)�A�����������Yb|�}|�� �&�ƀ�M}��ш�.�jL���&d"L�>�2�����p��A�k���o�ܱC��WѠ�ఄ�n�=�R���TZ�B��E�b�a���F}�|�OLcKl��r��@���Ҝ~�e1,�2��s�$�p=�3މ��~PX7��ˌ� �&ax?�m�x|���M��"��T�����Si�ȅ$�u�^�
yJB0�@Œ�zE��n��j�%�OL|(�Ӌ����4�����C|���?�{F��,����'�ZXx[��QR��mU�Y
����Au4��eBx������@�b<��duQ)RJ-���ԭzAM��X�+��x�⭄�A9~�����p�"���z���f���%��B��>�ު_L��\ ��c��70��!@<@�����X� ��A�(���$�� ��&�d�8(h�t�jY��Q�+e����2ɓ u��&��1j��RK�Z�I����Q�m�G��i~UW�؉=ð�fG�s3���5��vᑓ����O���ep�=TmdL
Ga,�k��
o� ~P'Q�?��?��~�Rk=D���*���b�e��5��HpF#Z�t6P���:�w$���NUY���Nw�<���c�"l�>�[�U�ύQ�k���m"����w�F�ɾ��X>�J��Ғ=����5��*սL,��Q�ky�T�2+ i�(U�\L6e�\��b`h#�Yg�#�A��D=�C�cCl�j�� ������� �R�"_�r�����Ļ�W�5�_��[��L�0��� ��p���{�����������/*K�P
�R�e��
��ə'�5�� �bҽ7���/!9��*�3��)�}A]���d�W�P��&��)쑪�l�*�v~!�]�9ԸcvN�C���^/�@��<�g4�̆mD���^/CG�"bfM?I�kButQ�b�E��M^�҂�z���}7�E���0�Z���Ðu�t@�ydJ���eQ0���'�D�WA�e��l ��� QJ�8�k�[31�c&e�8�#���?+U,K��=%���@�iN`}���� �v��=���M.f�&��c�7j?jR�c�rh�8��HaF'��il�N�2��2
�E��J��X�K�Ю4	4W��|���h�i5�A��p53)�M�4�w�Yt|n�\ӟ,S�XF�ةUr�b�fP�5r��ֈ���@���40Ή���]- 
�<qT��t����y�iy�!�7�*\�d
%��]��Kڋ��nùW0P����FQw#���b�<��G�ܬ(��6�ȋ�}�Y&76��T�KA�3v��7�˅����P�����@dHj�@@���wk����u=��x�B��lB�EaGN�����U���欠��e�4X�K?�]c~�.���-[��~����|�=���� .��֕����h/��n��V�>�>*Q1�lN�f��8:�eue?���G[kR�C�Aji�^n��Ñ���I��&�8J2F�p�Y1.��RO���ǚ�#�9���ߩ|��2�xɘ�[elM�r��wX�^|��#;��8A��$�	�N�HT��T���c-J�?�>|��Cn�_�E�x������@:����CA����P4�ӑ�2���M)��b�{R� �__���"x9�p�.��,,5CX��!Ꭹ>�l'i��
��Y�*	g�RZq �h\r�-S3{�,6�	��:a��uI~�mo���?�О pBw�ok�.�����K��ʂ�[��Y��{���^C�
jk�� F����O���MׄV���+�ڵ�8�2cub����Ƽ�li&tTݰ`�>��������C�'+�4ع7��021��*d���P��^��6yC���c����= u �E�;]aٸġ����2C��v082A���Nd�D6����(�>.���z�b��	|u��S��ثKi�Q��.�]e|)��;C��&LWՖщbz؅���(d�����+1E��10>�0��_�{m1����m~��};�óFO�|���S[�{s��h�-��ZjO �6�:#����f��B7ȥ�z�&���\f�U7�a2�!��b��<�uDA��� x��|/pj�e���$�>��9JC1��<t�4��d�����H!���Ee�*�RI/;aݯY����u�|ײ��#��b}ՋI����-)�g�J���רd��6o��"v������5�5I]�«ZY��d�R�^j��4�x�h]C����U�L�o���-ij�p\ҝ:ᓷBP�S盗?��l�&2=)Y���nB��G���OM���`g��W�F*?���tjʑ������LZ��m�X	��ls��vadT�6l�����ִ����m�S둳w�W!�aD35-fH�ϑ�g�sW��(�MCi2A��Y9�S���*D<��g�-�b���2�ޣ�x�~OD�Bڢo8���g�D�#T� 3����B�p��?��,Q�Z-�0#~d=7��Oӆ{|
�3"�.���͎܎D�!�g1@�r��������ǋ����ǈ�u��L3?��\�?�����Mݔ�a��}D㔁�L����ho7����M��� �KS������@�}��Y��!�Ĺ �b�O�_���f63W�����lEuTt�S�~\�	\4Jn)<dဧv��	0�H�'�:B#��`���<��!�f��r�B�� ���3�� ��e�{F�q$����H���|8|����`Z6�6L�r��M�U�� I�ց���\\~����3�'�bq�ֆ�#!���v�؈��6��z�G�t��oघ���[󟭮����s� �Ӕ�?r9���+N>��.h&���جGN�w�����]&�
������D�N�1Dh�zI�U�<�]�]���E��+�E�G������z�Fg�n[�}����Z�����[���ֻ\�<1���ҏ�֘�w˳�5;�j�&]׎x����C���j��SU���[ي�aj5��߰?�^���:|Pԝ��Y�"�L������Q��J����2�j3ށq�fQ>7���q�k@P��I_}�!�dr�P����%��2e�9MVrj�ģ��P�>� U:�kf.�Z=�N=���R踲l��S��Jb�-�M�LPG�����<��3����'���q��MԹL�Q�E�E~��������\�K�nW�ȧbnd�Q�Ł�llo�]ݛ_��(���9���?}Bd�͆ك�$�vg1p,�Fv���`v��F(���ho��Q����/O��t���'$8��S/�	��1%ymF-.�o�J���l�^����֑s~j'\��/8u��Z�>T�����E6�b�WI
��.�f@k+�/�0v��v4��=�\�\��q��=��?�5!/L�3�����S����>�]g
J�J
7��k����@�!��T!��]$�{�I�у>MP��`lo9m�eO::M}���)������Y@����������f��6���_5k����T�C�#QdWs��hla"A���E���˰���+m>�f���e�9*)�Z`0�K��#�r'�Y�Ƕ <��n{��i-�R�iV9z�#����tϜ�|�������8A�(������g%t��v��Mެ�'u��O����BD�s�V�S�ߥ��H��z��!�-��K}f��gF�������n&&�bJF�+RJ&�������f�|W.�4۽�'�{��PZ��dZWUq�*�d��hT�Ǒ+vm������@b3�୩$4l �E��2X���)��kk�M�_r:�a�]�A��զ�������8r��녕B~b$�)}bs�:Z���;�d�ѐn2�BMO��Q�O`ör߽7CM��~���J(�?��ϼ�!�L��s���=݇���Ir ~��d��̽|������]�����Ӧ׳����膚�p����E{��PRQr�`��J����}j�O�3z�Đ�wJ{ؙG�5�'�v�X��!J@��,��W�ߝ�Z������>��}�E.'�}�S�����wL�{u��b2!	�'��pQ���42�a�nTW����71�	��W^"
�e��|�2�HB.�k�׌��9��-֯e�ż_`
s��z���.�M{�v]8��C����٩���mk����{��޾�EK�}���
��T�U�=�x[�g0�#9��-�qd�X�@V�e��kj�7��G7ᔌ�ܞ�D�F�w�!ps�����Hs8S���j&ઘ�b0����J0')�����{�t�}H�Ģ̫/��V��r
�T���a`'��.C~��!˵ʡ�R���4a%:���&��A��B�Ϫ�9��B�I�K��	XG��c�3;c����܊ng�m��	����ʇ�$YW~���
��3���c���l9yD=Q�	�a��g�C��z�ܚC|r�<�Z�| ƿ鵰	���ç
�����	�t���~���4�.=TϨ8��i����PT����TS#������Wo^���t�c����5c[�9�5B�y��J8�����[S+��o�����qX,����5�+[P�������c��E��ڿqz%rؑZm]���+Yՙ�_�ӿ�,ɦd-_��_W�	��H��s����2}��x�z������o"�1<y�D.Z͙���R�*�"6v�1�S�"%�K��uXw��l[�4���7�9*]��Z	Z�xQ�����Dצ*�*;�o�����󼨵�F����q������g�Y1'�a�F�J�/�$%!�(��(�ɫ�..	g����\�D/뗉����Y�E��a�H�3#t�4���O��~�H`��0ӽ3���l)�b�?>�I�~]�+C��ۄyc��@zLD�J�h�����iĥ�XN�Ju�՛N
b����C�LT��!O���/� ��D�9/������}�w]����4�!#S�U䄗�䱽�1u1eݼ*y�Cw+�uJa�Qh�H�C-�u��j���p�>�[�����f{�ßc�70m�5H��^P�P5gl������_�!GIk�j�k��=�}'�������g�ܡ涫!�����|Nd#,d��U��SJjDkN6� ���'4���y�?�B_�L�Ȯ��r�ҳ���Qk	+p��ZhZI&���6$ +�ND6�h��ό�'~h�w��-��hY�U����|�X�H�=U��gE�6�g.������a}m������ЖB"f?P;�x7����D� $f�l�&�����1*O��[�J�ҋō��x
�P���(w�Op�8�)y�&Cvvh�P��q���iz�Fkw�X �Vp��Wh���`��j�1���ax��;k� �y,7�i(. �$k0��e5.@&n
�?ɸ��v�K|g�Rjr�ᕤ�n��H&���;.|�P~L/�%����p7���"Fj}�>�W:g+Ax�p�f�*F4st�I��/�ăd�DMY`g�'�ŀ�B�*L3d�#M2����С�~(��j����Vti�w�<DdS���ѩ����ӴX�9�9��Ke\Sי3W�!�-AI�ݨ�ޱ6�;(�G�2$�^ުU>'��u"gZ��l�(���8�V�6����͍�@Xt��4��J4wZ���̶�}D�C�H�I�c��1#�g�O��>��+�8Di��1��r��b�Eߓ�# (-���́���L�j���S�i��j�q"$�BwV�Ă�Ex����
)pD�Zh�t1��K�卽�״z�z'!�v|�ڕ���@�����͑IW-�${u�ʯ�X�YCda��˔5z�n'g����̙�)鲐\�\��r�u�-�����S��c��|Ԏ���R�<r��5�P���H-���cfo)��/��{D�V�ˮ�DC�G���A�^��׼��S�+M<����Tz�����ubnˑ�>H���O�����ڊ?�ً��F���@����kZ���A�$�^��3����D递z���	i�5�Ȭ$���q(n����-�������."p���eH^�d�ܧa��Z��ܵV��S%
u�]E�jR� O ��lƚ�&G��X��偈^�V�OtKBp�+��4e������䒋���k|L)&#�~�J��E(g�'��W+B��2�ڐޯ;���|���zkE�ΫcM����U3xS�b��u��<+7tޛ�����7��|�i�@�C0Q��%X�x�?e��;6/y+@��K��E�>%Շ1�u�`&[�j�$�R���)��A�f>�ȅ0����[���m��6^�g��s�`�c����yGV�d��<�V*M�
m�q����;�$��x��N����+��ֻ���E(]t|˥�b�v~-0wSSpD�d-����T�F��dͦ���;�z��U��Ś�s-��^��L4�t$���Qg�Bi�NG�t����[>>2}):I-JN�e�r�=ےJj���E�bv�>?�6%��	px�F�,�����D�_�=7%����V%�%�貐��������LМ�|�cb�d�?�X��@�����7�yz��rѴ����n�ʗ+�����:�=�\�2���R��\I���J�ѧ��.Ӆ��dȼ�� Y��^k��ޚ�J���:-�А���I�m���+��s��?eii/�T�Z��Xp���F�_�L�K���'&cE�A��-^J&z_;}��;������<�-%�e��I�u�������vZ��T�fe�Ú^�=���>�/l�K+�U��G\���`$�3��Mff�e�[t�LJ-yXr��f}ߜ̓��:�-���Z��6-lS��<G<��
o��DW�K��ғ��zr�����͕� �� �D�arJM0�'2��P�k���4�9���-%Y����5_��t�'d��#��bF?ђb$��{]T���t�%v�9N3�v�+Ǌ��T|�<v�ohv�zg�
|'68�S�,���3��.�?h�{)=6�C� 9���9<p���_$��Q��GC��t~1����k������nnIS���d��k�Ұ��H�S����ig%d���V�y�^ %hXDf�l�}}�CYV�Wr�qŀ>����8����y���}M����G�u����	O�ݾ�V�:{�Zsx���Wb�5۞��G�lq^qӵJ���L�D�D�3/�����ơ�r:h/Z���$���]Y�G,�&*� ����'|�2��-����Vccʃ4�����{L��[cS�l����v6_��a��3i� ����O��02��ûU��#���i��9+&�Erw�%[^���O�u8u�}���QK�VQ�Z�z�h��[�c"��|(��gs�K�rb�X��?�e�����
Y[v�ӧ�]���Kx�V+מ�)��Qd���5[5�4!�v��[l�:Y�M������F|w����@�U�y�㜠jB�6m���fu��U�V�1KƁ����u��u%�qU�z���� �"�ԯ��"EtQ�U"W����m����3���d�{V|�۰�\��}��I[iά���$����<sWo�[�����Z�|��݋m~��H~1�k��	oBF�:�zi���J��/��?��(��Q$��9Z�w� 7��q���H�����W���#���<�ͭ�H�+o����-q��G�������.���}�2�6!��$�]�WQԼ�?|���@�omt�]H�=�yS�aǵ~�8ҩ�ݽ�!w��=d�*:�$�0`$f��w|�����(j �Y~�&�b�K���/�a��QpG?�7���������c^ʎ�^O��%U�����'$�7�Od�C(��=k'�\DŮy���b�#�#�W�5��jb3��5��	-��h�%a-hx����%�B�$���yg��|nr�+$�$!���^��5��tI�x�nd�ܝ'����(��(ڏ���P�=�7L�2��n�<BJ"�J^dC_����o�@�!�z`i�n��1���a�Q��	z��jM|�6^&�u'��A��J�:\x4t=땚*Gs������I�J �@ rMȗ_�P�KA�v��OZ��(_����K2�Ypʂ����fr��JD<p�P����"f5�������=g��NY9x +�Ƽ"���ѿ��/���Jpc�Y����x�����a"؃q�����L>,d	7�~�� �Jv���	�^Butp,{%3��2�u\�I��z0�M��"��F�����%ƈK�㽉Dd�:;1o�'�f�$�~�_��T0�����{�6��+Vfq��n��Wy{瑒/?�q�8-6d�B�cM��K���Y�ʡp�b���d������F�<��bu�5���L���-g�T��ԕ���q���ck��rØ^��.�6h����þ,�D� i��'jd>",�Ž���l:L������D��{�u���r�D�􇙳�8@XӢ��)�Z�Ӣm��YBՂ�P/HRi�h���+���r��T����HM ���gﴄ^�����	'��L�?�bt׾����j�\(h^{)��s\��=4=��x�U�q���i̈́�]�S繿]����	�"�v���J���2�B���G�����rlv�+�Gu"O��ا����C�+��c'@a���6(�r�n���jIɈ��U\Ș�����^z��V�R��(��� ������O?N���F: ���q����{f��?Cel%�0i6��PE���w��CX����0��&�bTQ �8a�ٹFj��V��1��'g��������:�2!���~]���U�"鱽G��SJl�V�/4<i���Ձ5_���7�u����~��R�$E~
��?��%�53IA�٭�!;�#���O٢;��V庋�u/j��i�2Be�%�s�����q5�-Gh��r5��4R���a�X�y��c(WY��������r���g�0}��.ܭ]R��{��M�����B��T7�X���WO��-�p�ѷ�"�����I�T�7(�|�ђ�0���VUմ_B�VqV�0� �ϟgxr��k^����zf��e� ��x� ����۸a-��h~�v���1+�6�G�����`��)9~��QJ�K��@��ph8�o�
2�0gu�>�Jw���!�'VX/��\�S1����C[KާM��ǟb*dpQ����^z���
�j���Ԟ�j�%Ɉ|���r�^\ ���+�<�?0�ʭ<�ཌ�G�j�|�W��g�ɺ�)ݴ6h��
22�u�~����eK8�W����%U4,�s��-u�0G��E��u��7���jcǠc*�!}Ʀ��W������i��M]���>S�$�L�y-	@�3q���F�'�e5c9 �%�Q�~L���Qx��|�@���z�=n�S��j���m�R�D$�r�5d�ϡ�u��h3�L�h�A��qJ�\b
��#%3cmFL������l>A2C��?�Tp�+���Ki���0�f�m� :l�n$�לn`��p*������JG���'���;3j�S�7�0��U�[+|�(ҾȞ�V~[R!#���̉���>ZZ񺑺��MQ��kz�~��c5�
�"�Z�h�֘���i����Cg�|(��X"ĪP�M��W)�e}�W��.�m�]z��
�=�km�Ɗ�)�����Ē��`PUKaR�	��Sn(�����KBItU�L� Z�P�����ƔX�����ZE\��}[��8s5��]��}|�9dѰ!�Q�	z�����F�j� 8)upw�S�So8ɉt��*���xoT�-�����(m��Ak`Npª
��А�7��,��� �D�?W)v	�֔;�e�^����x�i@�)@��P0�K�7���d�<����'凟Ѳ�W���'H�g����<�c��6pǤ��0�1�,>n�r��!��a+��b�m�x�b�+�27��qb�M��Ӹ�ڊ��-�ɝ2<�~XP�`�ga#q�\� 
"���3��*���]� �U�#�O�,�RKn<�[��*m��Å{7�?��E$�
j}D���죌A�2`sf~;�\��^�m!RYo�1�n�2��n0V��j2$�gu�Iq�������d��<(8�O�?j�I��?L.�p3�+�묕������/�6��e�!s�b�Ԫ���ԽND�d痭�6b��r���Rf����i94�'�����W^P���}�kk����`O
?�a�_ ��猧����J�W��D�|���i�In��ZÞ/�;����<K��~�d��Em'<Qt+���	�~<<�	�2�YQzT2a����D&�� WVlɏ	�#4j�u���P�]GC�{�>�;,2�2t��,�mW4��I�2�������x�����#���,���ԥ�Ĝ��ҵu�|D ����F{f���lQ���H��O���%ά4$�2!ӼV=�O��Q��unA��]��!�7W��-1����?ےK�Iq\�x�����=e�l
Y���E{�x"��,�f۞��݄��_t�50�@�l��c��sd��b��~���N5/K=�+zcn���r���%&��i����V�ǭ�j�(a��>L�@�9����L��p�bWO�x>���i~Ѥ���H>��5Ѥk�D��l��WC\4P�Szr���~���g���3n߶
:��Q(��umQ��SuY�����VU���8���4��.��A���zy缼�N����$Z��o�B����I0m6��I�0��_�A^a$?l��Z^G`��i���k�?���;,47�[��G�o��Ҭ�n�5�zH4c�Ce>��
.}�f_���$.�{�x�)�"e����Z~�[,K�n�P���Ȱ��bOv��h�����8�tAwXKn��o��[zm���M$�k��d�ŝ�=��s�U^�3A[;�p�G%QCa�x�v}]��/[��CY��7�t6*`�'�c�L���<���|����׹��o+B-���t'�r�(CT_��2�(h�90�-��aӒ�ԡS�����k�l��xX �����7qV�Ud�&d�9s�6�$�3�i������1�c���5��
E9n�K�G\��5��4�8{���ke?ީ��7��m1�̄�C[�i�Q�Jr:J�)�"r�K����@Y�km{2bf6��'����i��J:[�����.xq6��YX����⎋��!8U5���y\i�f]����i&�Q.����;�eH_/�2�@��/�]��ύl��2K�f-jU�@��>d����xQ*����0�vH�Ħ���A����)%`��s�����V�;A/���0����ׂ��9���r�3��\o����0��P��n�ы��E����5��J�K"�k�`�܍�?��m���3�]ќ��)��np�~�\����fp.Z�e�C��&h�&ČC�@<k�I��ϗ�8l��8Ќ"#����M_�8
]$ձT����(*@~�>wG�Ԗ�֕~5H��o ���O�j�1Ikҝ.Ѭ��r��Q^�m�����ުQh�}��6l�R˯U�4����3-պ�
��7߲˩dO�4Z��t@� =>3J�=ܒX�y<<~��0�n��GX��\������^t餴W�.�ڨ���q����\���W)M}H�aNJT�l1�>:�q���ѱ���72[��Ri�TR�N�uَE��/�/���e�2>�~r��2S��y�R�f7�!�N���.�p�,���J��"�������*4fG��ou㈵�]k�9�&�p��((V��4�l��-�NOxM���L��v�'r��a������]��l:�z�4��>,��f��?����G��}c�;oҁ%b�?H�p� �R�qk9ptt6�JZ-�x?�Q�/����Wx�O(N��EU~h,��\���Hv�])T�Y��.�W�8��b��P�.��{�n��5w�ޣ���V0`�����i� �K�I���t��*' X���7�_�]�'껑5h�	iʷ�m�`6P����� 0c`��+ֲK�+��b�L%/a,jk�p������l�IݹbOI���q/n������=�|��n2�d5�<�4����to&�F�y�`�ǋ-Y���ֶؘ�f;�#�����r�˦��a���4"�Mm �����K�b�ǣ�F�r���<�<7PjS�0]	�UPzM��{����~HcO��ZgWh�d)����������V�wv���uG�����=2^y�=�]g|�����Z�8�s�k�l'M��A��ω�o�=�=�$�_w'�
4�n���#@2�6|{���
�o0�:n�^M��b�+ֆ����7�eI����[��qϱ�a:$F0��M��%����PXp�������m~����I4*�$K�jfd����*nS��#�H�}Ù��P��h���;%��5(�;�����eo���,����9�����H��rt�2�}G���}O{w�A�����x�s�>�4*�BeB��S�*���� -�����\��(���/�3��2%�ُWR%(�5����񠭮��y����k�#��q�:{A���<�W�NV ����>S����f��i�rZ�G��M�!:�QG8����M��-�6B��S:E�����ɭR��j�x%b}!����1���U<L9�N�ˑ��q/_��1���G�Q�Q_X�"L��M'hRL��Z(��s�PYʱYzƞ7�{�H��g`�ɿ�[(��WL�)��Ғ�Q,�3>����!��X�W/�O�_hU�  �"Y��&��Zk.e���=m(b�G��X���8�`ft2�LJ.�*_QtZ��Iq�x���W	�'ִ�P�g�����i8��h�`V#����Љ�f�w'�G����Q��WM��*v�l8�Ә쪫S@).��h1?��2|�A��"x@+�ZF�%<吞�������M�b����X�7�e�GS�+*_54ڧ���|W4,�l����5��5��7a�s�`G���`n�}d^O� ���̙H�K�u���+?�V�	��[�����Cƥ��:1ᓚ��X��8�5p�<���,ε��(�w��V��Ww,U�/�R=�0��\Ua�O+�1ܜ���S��8e�tX{Uf�֎�I B��6��yh}=Qq2%\VL���8H�J��w�JO�Q1D<�_B�H�iEy��G�$�ih�����Wt�Mz���T�]6��2��8�y_/[�o�\>��mL�$o �࡬����)�$ކi�%�H���$p�Xo���V��m�7�T��d�8�s,��m��1�<3�g����t(;q�I�nnz�9X�*�����u��d���2�|@p%���>>X�a���&ԩ����4b�� \���,/�+%@�	�ۯ0��]��"�J��C���vPQִi�ZT���8Qt�"9Cg;׆jR�%��.K	�����#���r�s�U���#h�ݬpofC�D?_	+�e\��D9J݊%j��A�I�O2�DX/s|zЏ9�� �u,6D�I�V�@pn%=Ё�6�7�_��0J�-�
\	Qģ�7ۄ�3ǧ�R���]:����U�$<Bj]G��-��E�Gq�hz�c$��j�A:�"��o�&?_�N�q\�-��Ӹ����d|]�������� X����;�2Y�'�<���͒ ���F�L�����[8�g>鈷W�m����v�Ǥ�M:4��y6�u�At���1SH�ģ1�d�j��;��"al}K�|��"Ug��g䫲�^�6][:�r���|d�
ؠEQ�����݉��Y����"aΉ�I����*h�<D�lҒ��.���P(�U��N.�$�i�)��7f��U���Z��4O�R&�?#��`��tS�KhTx"d:�\,ʱ�٨�_�Fߺ���~X���}5�d�"?G

���,�>r���l�X�oF�E�⨭�.�r�nGՊ�>� !�L�fY쌋�C��W׈j$#)� cxX0�2�Lvel]2�p�S�ap�P"�$7�&!�Pr�q��i�v�{�;!ʖ�H�e��-JI<�1����`�Bl��������ȃ���^���׭�0=��eL�M�ל��AF|
�v�0§nJ�/����zӿa._~��ܽ��B�e��hS� �s��܁��5��{�L�P��?�.����e��M�ꈂuT�^�@����k�׮q>���j��{�_��~��%7�.��H��)��SD�N��g��+b=њ��r�1�ë�++p��H:�Wi���Щ=��F���$���$���j�g�b��M��I�&�+�_c�����ƺ�T0D��Q�ҹrkT_��i8Q..�5V���o����H�9:���t�f.�Y	XH�LN�?,yz��z��&H� .n�ȸȃ���	[���"��{ڜA(�Hk��B"o.�YS�a�n'�}�CU��A��u CN�fsC�gL�=�g���0d�itK ��(�ᣂ�b�e?H�����k
��Kw����a�pOOADӬ3�zQ�;:<\	�H� G=�B�5��nd�;��3D��.M��	Q�CQ*��/���0��$|���j�A��9ȝb�^�'��G�
�����4.�`u&�O��!#�m�{)ȍz:QD�&�x��{|����Ⱦ�'�k���tN*����<ԃ+Bp�CA|�|U�g�[5�ȭ����se;�������e�����3U�H���ж��
�3�t�����D�(T|�+����"��b����0���ܬ�+.��h�&!P~�|ZO�P���V܁��Nx�������d嬉}~����3+@�w~��oX���+�_4����h��:�+a�>oaJF���i����zX`_�����h���f!���ż�B�j8֊�f�` ShR:c���X��}�P�?Rv�2n��9y�T����7HZ{������8�������ZN�H�Z,+��&w�^ʺ���>܄��!��^-Më?��0�:���eO�l����{�--�Y��Tj�\��WZ�����h�5;��B�U6ޡ	���Q����r�sN��Ķ�
�}yJxP�K�]��:A��zk�+��,�B翥��3ՒHp_��vU(R0�g3����e�7������!��y�p2|�Z�UP�LH��8:,��(�#�l�+�Ԛ�v��nqel�T6��6�#2�6��v�#ĉ�*��|��dr�m��q�V�!7���OOz�aj���/�l�̙�YA89C�O�q�>�� ��F�-=��,3�!l"NU#��l$�+�qJ�qa�ұ�v�$�ך��Ku��J��յ����<f6S��>�5���%M��m����?{2и+�Ҧ����i;3Jn�x��*{��A$� lڱ�� Y�A�@�U<��5��$*߯*�l#�9r��ԁ��Ƹu�� ��z/e����^�GM�y\��}��1��]�;J�tsQ�@���(.J��f�ev��>hx�_M��o����]we��2�b���N
����������i��.�nttU!�����s�p�'K��mB�v�!ҭlO���)��PZq$�O�/
���U�a̍
O��2�9&r=�^�4F����F��!�����Ϛ����w��.wz��̄��f�o8���8
i)�{~(��6�ߠ)�����3��tq@��k����P�����	�A�g#��ఴ���ƾ9(�o���Aà�	�J�k	2�Y�A�������fH�Q:X�3�M![�jܥ7lB(��$M:����GA�ڪ���h�Ç/�j�0]��j.=#W��ʾ
�1�q4�X�$v`޼�投���B �.Q�p��<�¸b��vN�Pp�X�aHA�2c�����j�X\Ƥ�#��DM�N�������dV���ea-�9\��J/�O�Pp"�"���欁��SDU�:N�f��jmf}��g�M�����a��=*�9O�޶�7��;a���?d#r�c����"] 20{S�Y�ui�Ϋk09�� Q�i%!�"��bmn���1m��R��cm����<�n��L،���6�$��)Bf���c�b� jsn����פ��/فܪקb�]�Dz�z�;�=�)��R2F
���
N�����	=i�v:���N�2��;T	t�!|�舄U7�qL�n.���W\ɵ6r.=�ƯS$f�J`u>L�%�d����IK��ْ@B�Yk����*��b`���ڥ��AQ���	 uq����is��Ɖ��)�����<�����Oa鵦l�8�����n�� ��P�]�<�ݥ2ז�5�?��u8�a�j�/�����7��1�t��>&�QUy
�U�4c�d�ʃ��3�U��=ƴ�g�QVj3E�f7v+����%�K�v �Q/���Y�y.�:ó4�����5"P�Ã}�1c�2�/k�C�I�y5��U/pp�U@p�����	��8��l데G#�_w���Y�h��ģ��O���ej�.>}�E�Y5�Xy�l���9�;�Yؿt�o�sJ����E;���%���b�TC�&۹�Oq�qmBp�0^�,�_ER�)(�c�n;���$���5L��Z�ZT ? ޅۍ=�'���ŀ���g%G �<��"T�����h' ��
^%5�(����r�s|4_d�������n�w��)�ϋ�9ެ�;O9�Q��s� �D��YP>Z	_���1'�$,�m���J��28.�۫Y��T�S�Oi��KGX�oc�kC;���<�i��
 QT&6]��r`�tl�lm^�Й�w�|�웬��ʶ��B`���6�++������s�i)2��Bt�<wa�g�s�"�~�dck��9���lL���<�p$}��w�j�L�<V;�'EH���L�����;9�`oh��d���@��V)��qRctt��3B?q��9<�8����P,ҚT'UE����;���(�Ra}Mz��q��(�5�����iy$ih$�j$�?�e;���1�4�Yb�R���"fKO�wz��}~"Z܂���^�$Lm����ˢ<Qa3cj�'Q�ޯ�s>��^p�p�Z3J��Q��.�O��og�����:<3:8��nq|&�c�]$.wf@��P҄J�J��eqW�z�P��mK��=fW������w���!�G�9���:�>�l���(k�/��9k:)m!�C�����3_�}�
 �~d��B�'�}*�z�(K��ò�	H؄dV�z(��� �O�-�GJ�{��TJ�Ak(�4Y���0���W�h�L����[j;�_6��~�K$X�m<rMl�95־φ���5��$u�v f�k��.ɥ��%'q���b�<R͇n^mYY����`�QJL��a`N��~�X�U�K��ܯx��zɾ��d�/�lH5�p�tǢL�o�Y�]�D�]	
���Ȣ�GK�tLU�4������"L�
l���?Z��2�J�����]-���Rf�st����4��Y[�ׅ=PɈ=�n
(�prɷV�%�A����v7 �ݜ+98�r�?π�P�\ls��N�֫��N̬ ��\�S�KBe����A��6�. +뎦,	ޒ�h�U����t��鄏mV�4���:R�	����4I�^CP�+� �v�{���������?���(�@��|M?���px��0�)t��R�l�t j�ЁI��s�yj��fyl���rmڈI?�d^Љy�{�^��mp��E�u�n�	g1y۔`�{����3��n�0!xRb�ē;��w��;>�|n9�+�	lע$�7X�g��?��h� ܜV��m�>�I��]�G��)+�~(-�a�j@��ǀ#">b�"o�8��E��v�>ۥ��ʆo�rZB�/�Ⱆ�}	<l�� Rex��!�*k�G��0�Z7��^��xF������@w���G$qYT9U�0`��3mlsc���mn-�Z	֩��nn=�P�-��f������������ޗc�e-��R[��� ���H����\ ���a����ynv�h����%�=#LZ��;`��>Dg��?�(��BP�NM2{܊D����?�u��4X'���B�%_!L~��F��}�R	k<�2���F����1Ī���#���cHi:V^Π�)���sV/h��:*�"��$O���|�'|-q� ��hH?e�,�}�p�9?'��⏐P_$�W)Ȥ;�ry۴sH���>��
�:w&���C�T�>X��>s�C������ޓ�1���S�z�b��aW�@���6���C`d|����N�l�%�+��[�*�˵���܂�mּ��c^ziSO�Mz���ql��d��Du96z�Y���J�oq�7����L�y�eA�����i���_���W�b<lL�ă� `�_|�-�@-	���v��)�J�h��_���6���Ay>�Q^�D���XD"�>�u�s�.�{s�̺(��$T�Iq^ă����+8�T�6�?ո�.�X��9�Éd|�����ib���������\!�.Hqx���J��!rF���x���6���^�v�����V�S���+}7x���#I;+���+�����b����X�ǌTٷ6�X���kp���9�Y <�WP״�)nV9�qLg�v[:�=�B�_g9q����gT��#�%	�Ͽ�fI`q��&�?L*�}+&m`���W�j4�@�rn�W�SQPL��,e�T:�8g8���g!�<�3���*�^�"r,F��7��"��+Kܫ�.R���?��`�H�5	�z�w_��Di��O������̉�ȗ�%�R�(0�Ж�{���)Y�b�x�|��Y�<��<�@��M�ף|�w>O+�X���͵$%��w�J|5R�K��B �����>������u'Гx�������dy��ti^3~���b��=Y}��i��w� ��uT�`ޡ:�������� ��E�NH�LvJ�3�:u6Mh�����T ��jmɼ��]!������us���o��ړ��)�C�N����R�jBc���.�н6Z���ױh�/���9,y�&�O�C�%�ި�J�%������?�A����e,��QzO4�C���s�2��B�����\8-��TC�M��ӑ{��������w��M�(ת�:����;+�9�Z�!v�0ά�L�iא���5%�4�Y��̷
\�;�p `a���2�T}@��H$S�����}�0m%���UG�p�.U8S��Åg����@��$��{�sH��:߳ᘢP=NZcQ��\�.^~��|������a�?Q{)�C���0�Ȁg<�d�������d=J?��m�h�kȳ \ �X�Q���s<ߏ�%�Kګ�:Z��=.������s:���ݡ�$NY{M�S���z�z~w^���өL=z������0�y���u�QF؉#8ƚp�L"qDw��a�8jǋ
��Vz��\+�n�d2�����茶Q2�J���������5:u��48;��!��s�l��N��aj!� CK��z��oAv�JL�e��\�� ��P^.��m�N���.�ç.��Ɏaγ�W�0��%BY!�nҙ���Aqx7�x���p�\z�*3��L��2���L�|$�>j��:=8v/��-��g�iQ ����!�	J���b�ڻ��t.����FdiO�Lɢ�F��̻T��6~��jS`C�2����e�~>u��O�V|�m�{��]����P9�90��.�_��t�1عc �u�,�]����x+ƨ8���F(w��9w�j7��E�w؝6�?1�6�qv(&�"�����s��bZ�v:�����A�Ѡڱ�����	g�iA5t]o�q��;�(W���q<���:�,c�^�!�����N����3�����X콖��|�m��5�e]�t|��5W?F2:��e�"��O�ӗ4���i[R�k�4�k��h�{`�D��f~o��DȦ��?�0�."ǊiS��Ym��^�83��}'�9 a�}��G���l �Vߗ�+ڡ���K� b�4�YÛ�Gׁ�L�4v �z��z��y���2<5�s�a�1N/߫10^ah���u�V�do
`���痤c�r��DZ��:7���:��%��0@�����*G׵�����a��K�|	�<B�J���1��WUA�<=�t��j�"�g�	�$Ɵ(�����g����)p�{ωl��� �̻�OZ�� /s�t�^S�l��
�][s@y�ҹ*�A��'dN�A���8�Xzs�A�H��/Ȝql��\S]pv�����lWX�*`0X4����A��l �A���F�u�0�<^��9/�'N����)$gW�A����p7
���x*��ԙT��jAL����'��2*ր?�
V�x��-��NM�m�ܘ	g4�b����w?H�q�5j_�/��P ��؋+E�-S�9	��d��|c��d�p�%��Avl�PA�l�>�L���H����р~�Ƶe��y��N�Z4|K��-��H�"�`|�gw��͡n��*�z��.�4�-����<�����e�L}�)�t�
�����֖)�?��6�4^Y�-�~A�+&ٝ��1Em�߷�:�)�*�g�xX��z]��8>w�و,��AvO]�V����r���rA��+v��U��e1?|�{���<��R7�}2e�����w��!7Vo!��?�����?V)i�P��Ut1�d�Rg��
E��í�hi��EW�߉�Lqk� 50Q���Vħ�q(ZX��zQ@p�/�j�z*�NНω�7v�����g��e�W�b�.�E�~&�)�iQ�K���?�=�!!��Y�>�_sz�!�*�,�ȸ�|�5�<�d�\��9�+��h(����oƁ+�W�*�����t��R)+�.�ߑ�ȶ�����R�(�X��?�'��sٝ����$��Ξ�?O^���w�"�΁�#���}���RjwEJ�")��� ����E��θK�i� �kh���x�{b1�}���²anXZ��nk���{�z)�S��k���R�A�X���
�4������a����������+�t?ļq�o�/o�$�4q��H:��y] �Oɹ[R"{��g�*Z�n��<�`m��G6ϑ�������e#2��p�.L]:�*�ܵ/Aq�q,����dO#Dal�A-Lϓ��@/���!��3V�� ���)p�%T�\�A�1����H��'�F���oQR�T�0�D���N�i҈�Ӟ�U����gQ����n�x�ɣ��&�g��m!�̊�kzgIm��lMe%ozͥ��c_  ��Und�jV��pYǛo����*iI�!����]ؠ���H����� ��T��C�$xԺ��3@�D�$������� ���tu�$�c��kg���<�NB��]y�v��wT�EL�0Ś�𢤖���ϗ��rwe~�"��)�L��I��1�o� ����{ ]!Ħg�(�b�1���҅��p�k<�b���ѿ�i_��G��Č���r�]�?%�M~\Mȁz��&�0���8V�QM�w�gҦk4�vH����aA��u-BJ�Q�l �A��es9;~����J���7��v��є��lW���Z����%����'xk�ٓG���ƅm�#�"52��D��O�t�`U��ᨩ�/���w���q^�^Am��tS�nt�{Aw�[�JmM���ŀ"�=���G��N��|X�t>�b���*���z�Ջ�s�#�F�)�6ⅸ��b�$�'�:��&x�֪؞�ϙ=&~�rBX)�!���3�8d��T�)M� ��'�!p�����BH��c�G
Uu }�%�L��Y�ٻ���	�$v�pt��cS��{�E�Y2+k�qyq��DS�TĪ�hP���M]�Eq�C��ᚡ��|�.��� -�)2��v�I޻!h�'d�� WQ�6o�c�[�c��V�V��7]�������=:1���ӟF��" ���8h[�V�e��F�%��xW�oOϗ��	����R����+ӈU<�ܐs������H�B�Hk^��uq=!g	�6;���>���=��Z&���:���^�0��P۷X��wc%�*��վiMj��z�f‹I���F�*�9E^�*D�Ԓ@S�Wy�GZ١,���Y&<v�{�i � ��T�؋al;mƯw���Cz,��NԨ(�ԛ��gR��MS�>�^|��U�9y��sGr�$J�: H��0j},�gh�v0���"Q�2�.0󵼣X��1�ѥt��[ϊ�,�JT/�p1������Ē܂�/�n�?ć�^6x���( �����]�Go,r�%�S`�k��3 �����(�M/��F<��DcRm�m�%r�d盵��,�r��!q�<$�]/�;��)�o�mx����m{� W|IO+g?"Qm�����<���M��%�q�@���&6�+d����T׍a�X�fs�ch�-��W6h�i�X~�-Cv���N@>%�'�L͖����̺��Z��2�p�����vc���->5b¡�I�Ɍ�u�ks%�`TguQq�<�r�d<o�������� h�6J�q�P?z+l$~�X`�|�X���࠻����<��;]F�3���]M~cK�R`	�������}�ԁ��B�3(��*�z4z�f�1|$A���;�o'�����9�E(Ui�V����7t�i�~��j�^���)@��b �g�6������81�<����/;$O8�҂��̼���R�	��(���<g�TG�.V>]@�2�*�Ί�ΖK!@�9�7��ܟ��f�B�7�U�jPE�����S�8כ�Leߐ�����p��T)p��0��1�F(С�3NŒ%���G�8�X;�������!J~]m�^ �8����7nvލ�7��F�j�7ך�r���<��F�$͆Ѫ������:c��S�!�;��P�[��֐�M�H`Q�{fC������ ��n���fC�1c�W3�(�0P���Mv�� �Al��O��Pj�7ERx���^r"Dt���#4��N�ۉ���2����/�� �k�#«���t�r�X�	�����X�&f�P\�W��q�(��5��j��p	�o��8�^w4�0tfL3�n?�M�ՙ�0�����IN"�#���4��=5�s����8�
��`|�E�XEX����h����@�p�!7h���l5��NA���?'��H�S�I��#V=!��4-��P�<�yq�k�;[YD�}�^Ɏ�	���V��)
p����Io��Р�,Ɩ���BAyx܁�Rh��O�ֻ�Z{�ԁ��a��Xe���jN��-BS���x��$�q�5��:�&;ca�,L=�_�{���~�y� ��	d�����<o��5�����XvW}y.�q�q�F	,�5&u�1L������@�V�V��ĉS@������V�˸��e�x������)��5�0����n�X��"2�ÖW==%D(R�<?kh��k��v�(|\L���/��G�N����:>�?#�=�e�G~?�E������A�L]���u��܌����5��@#��x2(���k�.��q����/u.�P��O�&��=�_�Dډ:i�:Z�q|�2&�U|���@���MӒ�C��A��+��;�j�U��{d�k-�ˇ9o �1]I��>]�~��J��Y�	��E��gE����� �����>�n�����Ҏw��O9�T��=�]�a���Zf���[#X-��CNH'����`ci�0!�9P{��h�L>ۀ��(k�]Yc3����|
��=��s��qIE��i��W�c�PtŬo=��4`|4�&�a��P�Sι<}{��^`�fA�~m���P����ܞ�k~���ۃ:��}v�G+}O{��X}I~P�@�%y��bHv,��gTo[Ͷz⹾�E^,2ґ���0����OʐET4e?��������i�� ����:���u("z4M[�)�u���������Α �sJ���~U����d���4%#4P��������'q�hf�m9�5��,_�����"w��D��փ
c���d$+��p
�͓��`�;7��C�/�ou/�����I�3N����C�D��`��h�eӻ^�.ja�!�E6�te�u����A!����;� )�',a�������NRKw��/�2�Sھ��v����N��)^PDtł09E~�#J�|JDϼ��[� �]��*�Sj�0��?���5�@,lj4XP�����^POq���y���b�1e^3�G9��2�+)�Zw���*��;2�������\��aiRo<p�n6�&Ї���S��K{�1���jv�kO'C��O���9g�a�C�UM��O'����r��t����Z�O�
9A��τVk�e�z$)x�좗p!Xрy~����b�� �|9�4ݗ����Ѕ�]i�����&#Gm'�����<ѧ���1�\,�'�Y�k�?!-� ���>���	�5U{�k���g��<''��j��a��+rueṆj�9y������(RB�S���o?*$�.� ��M�p�Z��)Z�	�ʭe�ɢ.L��* ��#g�j��:��R���z]��bԚoDT�{�a�b��X�[��&�0����rU2��L��[;�ɏ���J��abO`�	R�z�ߝ�l]"ۙ��L��\����ٖut�4�����ׅw��B�t�P�mRN�}߄�O�b�J�����`� �g���(���U�&�����F���eJ� ���P�+
�D�S	 /��$�f��%��O�����HJVJ�)S�Jk���c\;��K�q#�_IR½\�_�|rӌ#�LK��L��8��X6W�襍
0��u���	�Q�1�,�k�bj�O�`�)ٴ�b�m�|QJ�D�{$��U~��!r���s����3!����rh4�Р��R��<a� �^���p��	�o'��h���g��О�a\KXh������V}���rshF�j��"���0��e�lg_:�x�%��d���� _'���q��u�<�]�8�"b�81j����_lV��ĞF��D�ʃ�Z)�Tϐ�����m�}c����Ob�.�hG`���z���Y�F>�- �ќ���p��UPR�e��X�+&>�y��;ʹ���b���ݥ����]���d�΀�=�+�j����ְІ��K��i�E�Ij�[H�t`6V���|�}���.��V;1}������0a���|G?R���W-M�S�
s!���Zƪ_T��~�@�.�G ׯ���q�V/#7H��_��+Z��K92c��/Fg��.#`̛�c��`f�|9>��rhki}? b�k�w��L�G:~:�Oa�=`t���uu���[r���)t�F��u>���$Ζ�v��O(7�Z���4i)�5X�<@���1��pK���D�����y#��z����hY���H0!����Y�&T[N__��M6ytK'}�9���\*�7���t�b�У�g��H&	?1��	���.�6$�b�ސ�e�H��Ȁ�8qȌ�4U�YY fV�G�e�6ט���Rw��i�ε!�j�A���@j@p!�#32����#τx���O�͉�-Z��S�hW'�"58$~ΰ#�{Ġ�yf`�o��}킈$"f �v��L4����,8��pq?`�Č��)Zi�dvM%TZ�����t��4��&Sm�	[���ُ/����;�|}��vB���x2%8�.�$;���#����Hp��0���,����˓�y����>�C�om3^{��Y�*��
�3�?���	{�ҲO��p�c�st9a�;^f����o�"��w���t�.������:�˖zk��Ʌ�����$Ѷs���ʪA�����;��`༜t$���g��EA#�P�U=L��:����)nSd�m8SW�T͸�:~iI����Ads�;�g?��WR���`�+����ݹ��&�/&���"Шq��P�] Weh�:O��=�d�ēR�DGT�M1Ο�B���\����]u�+� ��C���[)x���M��&@�-�s���h@&O�6j@;榓R4S���9�{�����C�}�Y���S	ʽy��W�7U�n6_���5Ad�ǧ%����lo\�կ�{��A2��[UVEn��?�J� H6���^_l��G�7E�Z�s�I�aH2�B�Jz�C�QPj�Q�0�D;x�������*�,� y��R��|��7�>���3ʤ��1-��E�۱N�0�aIIl�q2Nv� �p�t7�$JaٲԚ��xɶ�/_p
�~#�y�����{���y�����c�"P�t@��8ꊬ#]�z������W!w������X(��������ẕ!�}�P��⌰!�IG=�˧ <��ь<�y0:�2��o6Q��9��5��?��k�}�!�g'l8��yX�0�]��p!ƥ���S�o�!E�xt'v�I�Js]6Uo��&n"�!F���5��XK�JZ+�f͂8�I��Ӡ�B�"#Y�=)�^�
�B�ǁ��nF�y6N�!w�s��
*��/���|�AԜ�!�0� |��*q>�Qى0\T�PcU^���g�w1����E�p�E�\�Yχ[�_v�%7bq��������,���/Z�����՟:"	^K`���h]�:#�d�#HХD�Y�B�b̦��W�2����;����<Eq��gL.�U�"�gZ�	�~j�]�}�\�2<�B\���Z���4ƢI
V�\�u4 ��ڮ�1��d�!��r=Z�K�0Gj*�W;O�ҽM[����*�X��g=��:�b���������R9H�k�<=�?>���]�B��T��L8��k���<�!il� �r���'/!��2��7F�\����C���a�P���^<�Zy�
ɵ*���'�N���1�촥�<@��׾�zַ�{�b�I���@���Wh�.XX0S�o�x^E���_%zg�9�a�o��z{4�������i M�����_�r��t�GR�`M���o���Q�a8U(tW~�1 � 2nj��"����&rz����ܿ��}�8�\;��Pb=νWYt��͡�zp���'0�HP[�4��~���Z�q�2��ɜ�EsϪ���T�B���~@�TwF� ���
�k�_�|츁����ZO��,CP}J�̘N��
�\�(Q/��ђ�E�$9�7c}�r�J,9$�ԩ��0W�78���VX��dP	��>îljՂ�����'��{�8�@�	�?�����ҴH�[+�	����9�3���l�;����͡�?}�����T<<�b�^�DƗ)$C2>�;��v!���)��UrV̸�_(&�1���+�J�v�}��P�0�/��#1I _�0R��\�[3�<�w�cM��m���I;�Ij���^(��\"��,���`|P(���n6�=R�;��+�A.b��8A����쭩��7��e_t��n��6�]ճ��lq���ڠz�A왿�b��7Q���0�"V�=W��AБ������ZF���a%R1=l��f����6���{��Y���Ǧh0�����9����چ9��(a�)�l2i�*���·�/[��g����j;�����ރg�<�!޳6Gxfjd�<B���g�UJf�cv�,e��^��K�<N���GY��A��'0�K&��	�(*�bk�K6iF�J�!�D�_R$1�7_a�����5VRWL稉�bwj�VAL������[���bI<�`ۋAv�'�4klJ`Bv砳��k���}�S�ی�@ p�������u\�x#����¢ܛ΄��=��2;K�/��Xd`���V�7�m�ၖ��Z����[#X��Ga��͡� ҥZ�]�%�]�9�Ç�m$X'�x��e�	/��ޥ�'d�W~\�ڟi\r�1�À�v�����+&��{��z�d$�ҷ
�G�=����5�d��Cr	 L�&��\{5�L�?L�����j�U�Kb�[cL�Ԫ`��z��C6���ԋ�^��>��j�%��9q�r� U�<<]F8G����V��H���Na ��z��B���� �C�n�?���ے7�b�dM���	tp�f�W�$��k���:�D&���4C3*84y��J�X�^
�w��8�)#ܱ.x�\��&�~{�T�L!��
l�ܪ;�׷1���D,j43�L�P)[ܜ��-���B���/A�h��R����^mx��������ڡf���(N�\�}�a� Y��-�����f��&U��L��ԍW�?����[�c�>D3�p�'g{P��(t���;�**�`�qf�h*����*qy�8/�+��!~�]���p�pε�����_���9���-ndzzkGE^:��X'3#�z�"p������'�y<���3��E��//f����f�4~d[(�b���ʫ͏Ƈq6�B��ќǞ���ȉ�ư����Yqe���;w��n
��d͏]���t�6����5aj"���A�u�b�5�\Z�����ֺ��	�Y�>���d���z��k��4��~����֏�m�����r���4i�I�]}��TmlT���۹׶o�
*G�1O�.}͋!YE,��ŕ�滆G�Y�7	,�]A�9��h� #�e ��9��ɞ'5N�&���߮!���ep�-�>ϫm���	-�d�\�0�� ��E���L�|���%��oCK#9Ʌp����+o�>�"~Ɵ__,�0��%��u���YԞJ}�}��x����4ĮQ�`��������� �x��DQ��4�e
g�NN�՚��k�����7G��<�F�39�'�� �wn֏-���I���t���25��=�~����8M3*�
�
�_�"�)Z/�v�bj2:AP�)|/3|���K/�/ޙޗ����3�@lً�,�`ܢ-{��L*L�Qj��b�Қث5�o����8N'�)7�}c�+Ö�M	�W�?��Y�D�O�s�W<ܮ�y�Ć��ڣ��*�u�b��qh �BX�k\��E��`a�^���;Qܕ�y�k1`HKد��� ��(x��zp1�~���9ٌҥ��x�,����}p�q�=�{H�w�+�x��Od����j��b+�h�q��/�c�4�l=�actZdȴҧ(���д�4S\����P���Wە�ސ���������V����Q'>6��:��Ꮳ�F�[:lJ�����!������v���Q��}�;wt�K�,.؃�]q�����F��D�'���7.���_�̙6����G L{�]d�<�T��1E��_��n%3��F��Y�Z7i��.D����ÅT`	W<���?�%Q��犫\��5A�	]G����+�����H>DM�t���D��3ߖ���)EP5�s��X��)m���{N�K�n����>e1oZUL�������q�s�)5H\c����:k�}��Q9��.U�P�Ց�ʣO�U��y���3)x�	ɳj�
��SD��M��~	�JN��A4W+�})oH��*�֘K��ځC��Y]��<{��a<�sh�K>�f��ye��(h�v<�l�w�\yK��6 ��U|ABx�Y����8P5B<�}L\��(ߖ ��d�����(u�����f���4u�9jU�J��F9��2ݿ��	�h��?ɕ�{t� o}�5r*�p:�N7�ڑw:4��zs�hL7�6�t�����O0�UYDoݥ��'d��0]?����U��GD���xI�����PE����CP�2 �\?��C٠2��9�n���p��Y+���]w��+��\Eg��bq4Tp;�X/
�K�:��q��_+b3�S�\>�y� i""�&>@�5��D��d**�z�1|C
��� >u�ߩUXէڛ��4�۔�C��ր����;�"�V{��V��LѬ�����w���b�N�CK~
.۫���*W��m�hQJ�9���ؼ���((NI������sp3����y�O��?��Z� iN~uS8�J�i_b
<tS��~f,�� b�Pl1qq�r��(�Pm�D���Fs\K�q@�N��)�|�� Q>+7V�)��h��>� �e�H��μ�=5�����Hh�M�f(+Z?-�h�Zi��M*�A�&�)�l�P^���3�I>|����p���Ž�b�5;��Z����="A�?���-�Z����ts^PSc��V���Y��u�o�&f���"���q�A�7��>u��b��ь��@Ozai��"D��Ǿ�����ڟ>�~1J*��k�9T@�τ1�D��s|����9��R���(Mk u�{f��+�b�O=BȆ�w5v_��6��8pXB���P�7@P�l|a���L�Q������f��r�X��Y��Y#���T�:���)����D��8w�T�[U����ޖ�7#/wc�g�9(�mǞMj���cum��c�vr���5���U^��Js�oc���� vμ���f��X�8����2���=$�6��d�	;�F�a���XJ�o�7�=>�3���%3t����&��� ��-Լ>vR������S��M�� ��Vb��B��R�^N���/ 
%���u��'�T\��7>�V��R�X�cQMm�D��r-D�D�$���ل�H"^�DN˼��,r���}�[��	2,ݪYv�扇>�����V�2B,k����!T�ۊ�ե ��v�/�P��oD�P��@y��}�����1�C->֫�X|r{hB(�ӂ��?*�O�����ɛ{�^$���C*cݮ3�f���ٞ&F�Z��44�=�pVɭė+7�|�	���͸o�'I��m�.3a��F([XX��{���K�Q��)d���T���m�sd2"�ܿp����Z��d^��o�6�M���k�.�̓�h���yB�>Iʋg9�7��칒Q�ZS���Y�L
a�_�c:�V?��v��l�Y��w���: q�~$(
�\�D�%��¼f7^��N5w��Η���A�N���H�T��P���J����[9ү?&�`��a�(���ʝn����FuT���U��'H�܃��]}?�㪽���M�R���Jz�2��<�	A-�rʦ.w>{���2"�AgHT�JԾ���AҦ�s�Y$k\��>}���r�,$�.��!�w��i.�J�	s9��\B�����a�8З��::��f ����4:�f{ό��a��Bz���%�gkJ6c�!ȅ4+��m�\���xK�D�4s�S����{F�b�7h���-V�0o|�a�'�NI:�Y�f�o�Xa��"�XT��0��X�{�גx���oJ��%��Y�W/���W�iV&�b����m,�b�96��X��"�p$��>��>v���8t^	>�1gZ�x�v�)�y�b�)��E�{D��W>WI� s#�U'�sϟu񩕻��L��q'z���e]A	�]J�DS�z�o��Z@]�?�I�2�#٤F��f J]xQ� ����=v{h����L��@iDu�!�������6�;`DY�����,iF
��ʙN�y� #��x#C�l���0���I.-��T��_ ����pwIF�wq}����J�0������L'���+*����fs
kwaV�����D߱��[�;`��SF�MX�~�ԧ�M�L(�k<��V�\���rɡ�m��Y	fI��o�0�2��J����g�M_�۾9_q�:����"=d7F	��?�e
�l�&c��;6��gSeP+�^�G#e��q�D3��F�l��&x��I�j��g�Z<"�7D ��q/��R�
�ߕ��.o��o:c��`�7|�4���~K���R�`G8�r{�ĄU	��N��}�8��-G��YH�E K.t�nV�^D4=�DS�}dձ,��.z�^6!�uV�"��pZ !8-f���c��y�-hﯥʗ�b�>@[�y/��y�&��+eY:	�<�e/7�:����U�(��/г|�H�
��,�HI�!��qjye1=�f��8
���������5�6�2A��u��� �i{�L�5���h�֮l�jhĿ����|������(Y�gKo�z���]�@z^ �]�ϟ\�H3Mn�o�xR:��V*��צ]QF��"N��xB�����8��K����ҕcO�̧uɢ�?�T��v�C�
�H�b뽋���	F����Y�V���[K'�x����V��<tgsjCd��\=��2��L�8� � ��N�˹c�}nw��AV+�J�8jKz�qg:��cn��&��1f�|�6�%F��|\��mE(1zH
r�Q	nbT�¤H��Р�p�/���g�=D� ��A�(��&��t� K��'��;��V{'�.����JȻ,ϐ�h�n8�N[li.����ί�3F�	�E}B]]��oy7��2yQ(�C�҆<3����I��l�t3AN����V�n������ �թ���1% ���j��N���GR�$>}���<ߺ����o�GP��\l��2��a���h�v2ĝ��f��ߖ�^�ʖ_�(�m�➬�%|y��z�~Fqj����f��'ہ�OE*$��vc��p�E�����B�� ��奴p��tU��s�K����/���/�S���]D���$Ou�1�Au��.�|b ����_/l��wUj���b�u�#��&�2K�	R-u��d}}S��p*%+Eݠo8gm��i#rklr�1�Masb�0˗G2�4�SH�6�-�:u�����%��N�;W����𨅒���`'�9ާV�ޏM2<�ߨ�~Ԍ����4�q+�����j�h�,F�/[a��&��e�{�!��c�8����&hf�g������ӊ�9=^�P��j��� �N ���<�j�yr�݉�Z�4u����NĚ�������"�cތ�Y^dH������W*�g22q�JI$�^�Nt�,5J��㨭���[��LisU��5�� ONX�,�ϩ
��'X~v5o,,EN��
Ƙ�,�0��il�-`��A�U���߽zC,�^8T�|q�i�^�Ϣ/���N�[V���p���l��e��ޕ�?Y!�K%�ɐ���YVB���u��&�I!)���^+8�,z����!p_���?$� �*�wC��jlEL� ~�ި��"C�*H�]~�٠47����jw�WԐ/3�Z�N��/���*��r���"h�A ����w���vS7��5��A�V}��Bh����D�AK�+weS!O�n�	�q� ��:�U�?_���յ�K=��x!AT�2w����=0�aƩw�^�ђ��h=��Y:���U�����n�\���!��:�yۑڞ����e�6"��	������V������8�$9�q 2-�"��pxL�<�)>M�w1+�n|��j^^�e���9�WdCDE�Zz5&wொנ� ��Y�<UDX=�ܥm�,Ou�I*��w��	�0���m��c��I|Uc��VE�'��t1�!*p .�n{�n���c��j��ϰ�Q�"a<T8��}��Y��!�z�k��I�P���v��~D�A����+���Ns��Q����G�(�̎\�լ�����ʃ�hq���ܠ� :9֒g��ͭ�N��^֋/����VS��V�z5����ƿ�ⱥ�����`%�I�P�~�)�Tu�rqY�r��6nύ�=c�4]q!z㈔fn�'D���(X��n[���6TQc���]6׋Z��;�9�6��䬲�E��C���`7����|�__]�̽l}���Pi�u`3L��a�=Ů��I�����K�����=�>�Fg?���-'"��R�c�X7?fXL[ڜ��Oe���F@q�}|�t�k%Z	�਒�>W�C������T9q���9���������v��]f�&�gșL*���Qj C�M��@Bj��_�\�d���t+_MyzK �.�\L�H�h �کU���DZ'B$l{�+&�}�`�C��*"d_6j�Ok^%���%7+0V����w��(�1[����&�f���Kw�'�#8�<��R��W�K�i���>P�?�A�}��F�JN�����-���jߜI.��$W�%4\]���JO��w�Y���T��`�����^k#&�\����v64��"��9b!���iy�����A.�f�+A�f�?���޽&>�΍�X����I�G��Ag������`k��,0隣U�\�ܽ�s~TNSx�X%J�A��~
�]8�g���.�C�-Ѿ݂��3��.�=��ʇr*��i���ץ�޾��~	9d}eU��)z]�d���b`+!9]�<p��(���\�Jċ�������	]�|���\�m���T �s�l�=8�"*w��C8k2���m+{%��l�Y��*�L���db1J�(/DO����/�3I5����~�����Ⱥh�Ѥ�Ǳ���«���M�/��p�7���)�������ѽD��I>[ފU��6f ����6��ՙ�����.V�1K�����8�3�Q�!�
a_��TY�빮`	<(q���C��~"X�5���G/����5�ˑ^�/Q��2��g(��@�~���u6� ��W2m�hʾN�J�@�Ǥs$J;���]][F�97l����W���{��	,3�����C,���
6�I��wn2z����`���X˶��r���܃�jG�'{�Vm5.�0|�KB�?���Tp�&��0�	L�x��gåM�\�i��Lms+�:��n/��unsR�SbUg���	�Ǿ�Q߉u�� ��At��B���TC4����֝�ݭ�����k�(�@�	0E*�s�E�l�ܖuo�5��G�<Za���*ǩT�K�����<���R`׎�X�&T����Z�E�`%[C���1~���|�;���۷�'�{�2�SqF��$����C�D�]��D�>��t)v��(\��U�F�#&��fjbD8��Wh��|��$u�� W�)J�����t���`=_�C?�|�SWG!�`��\���*�/�M���cB>+�K<��%�Y'��%�H�<T��<z'(�ؠ@O D���L9�GH�9�=� �J�?��S�V�:|��}4���P7*IE$4�oG�*���c�	���9�td1jЬ(w4�L��kf�&{�⁲~��C�)��J�B���M�䭮#3��{��?��&\u#�Inh�{Nz�=t%�/��������Q���h���1�tǰ`8{wᠣ�8�7���+�^�Ͳ�f�pC+�hK�Dq��v�Y�ϜVr�8J��B ���I�Јٟ?��]{/�H�	6�Y
�����;��]6
���?�.�����k�8�����ç�+^�#�p��ml�α&���b������^	q��s�avr�~f�)� ��� Dݡ�繃⭆�� qY>'ʿjy�n S�P�*���rET���A[|����A �j��+@�w��z��C*�����)q�-������.�S;f��38�k�Y�hD����&I��� =����t;��c��h�f.ƅ��
��Z�������3u�Y�j��ep�a� R�$9`]''���ؗ.7��̥~���]���!��vdB�CL�Au#q��#ܜ�sf<~-��x�@n�8f�%�S��M�x�0���X��8�L+��Ꚛh��w�M8c��89z�AO�P�bɬO�4.�}��~�%��,�����c��)����]��(;�f\���G!�� ���۟���6 
��~��ٞ�c�ui��U'��|����O8�畂wc�Hr�3���j��
�Hٙ��v^hiQ��}|��E�㤡p��ve{��5-)[�ԉ��o�9� @Cl���aˤSA��N�=
��k�/��hf�X�����= �h��=�cp�<��fU?�-I��=�0���-����x�|Ό���gpȰX`qW�����i�W�u>���"��~�e�ZvuM�M9����qn7�ˬ�f&�uS���Rcv�Z�3
%t�F�8��ӻ@|C�(E�ae̖)�Z⻬�^N��j�\����^��d)sf�V�(�KI�����a��S�p��yMnЩ��t�$�`�L6zR�_#���՛�OޕM-�篭D�V����PG_b��gz^�>hSu�l��[�C:��Xo0���휲&&"��L>�f��0�� �3�mv*&܁P�x�$��b��,P�X�풨'����j����>�2�:�/8��4��0L���ֳ�J�&�-�zf��IXy8p9������/�c����#/�(2QtAQI�k���1,�^�7b�x�"k�֎��T�2(�%9�^j�43�������Y_T�``�u����*4���A��U�gO ���H�:��6#�uP��s8�����Y�B_�K�0���k���\\Z�qh�^0[@4��$�c��z��K�,'�<�b�| ~�KI��k�B�Fdx�^h&�盾>���dmx��?�2�y�T�-�F������O$�%I�y,����M����Ȧ4Q:��wR�qxUt1��_�ފ��4���+rW�G�~�4��Ƒ�H������k���&�G���K��OFuB�"�ȧ;8ȋē�8GC�%ۤ�0m{�ש���T���;�o�������?�Y��v��P���`�R�Kvў���"jEZ<iP��%��2C�R�'s5B����t	�w�.qX瞸�	�JȲ���C�R8fxHD�{�FQ�p������c�2���x�wZWT�(��x���������5h�d�[�rZ��n���q�}��b�$� =�;�{	Q�e�ج�~IE�Q���`h��Զ[�=I�Oͱ�2��/�����^}dR�1�`�m&$6�����@�R,T]�	]��J3�Ȑ������`Gh��]�_Zm���/B���w��<��9�÷)kN�b5?�O����\�J��9���J����Ȇ��oۆ��F!�xB�0+���
�\ϵ�DS~D�[ph�Ճ�`!o[� ��������k��g
�}jm��cv@��1ҐsHF��sB�&�OR*)�N�t�`x]�<�������87�̇�$u��qA�v;�2�U3�O�@�ᮩ��{����X�Z�)0L�tވ֗$���i��'+�Y���W{6��H:� \��L���34`��c�0�¼��w�m#Q_��R��6��9�D{h1�K��>[��a�o�H,\��&�t#uj�dg5.�!��-��U�x�6�d1���*��^�d>�v�E�~�X�*�V��x�!�L�<���*�+���|R��_�Ja��d��Q�����#��,�������v~��[� n�x�8��JB���1���M���	�זFv�ו�6{{y3J���eh ~���{�o��[i��by�����a:�Va����a ���!�s>���-�Y{�R;�I���dj����� ���J#a���OZ~��V�p���U�ccD�����Rtx�fC�yZ�8v���~v�N���� y��r�d����1G�L�oi;F��@PH�T�'�+�(�A�VTs�$1���V���8�����G�v�D0��?�11ւq��mz�Ɠ	�sM��蓬����	\ěB����P� ���~6�!���1��,0�{�u�h�~�R�B��4��E���
���s
z�J�B�y1ɺ�܏��^�@_����|�aP���7;����H�;�����:���PAJx��=��8Mɐ�GM�����F�\�E͇�	�h����v��۶7�����>�(B��/����v�/.ah�0�m��ѝ���H[���]d�9+�#��E�H8�w�=���:v���g�G1��*|�g@7��&��S�� v-Pd�M���c��u�?�w4X�袍Ʒ��^B!ANE�nr]lv�7�F����2�L$�?䔨�)r)��x�ю�hL�Y���Lw>Ɯ�Ztk��pX�(�\�֥=��[�k�PX(�q�7�ޖ��2�>�Z�����d)��H�$����/D��&�������!LGFH"ҺM	���8mU�HP�П�E ��ѱ�>ԩ�y"x�L�9�P�k��v9�)�4Z���N��	a�[X�د�1P|D�[�g	~3�� ����}�* ��4~i���T��l��ӓO�V�������"P����ܳL��>��O렑B�G�R�ڛ� ���̨�e{�1�ʸ>^UIh�,q�AD��:Dvq˰u�2I�YױxU`�"�ݖ��aC��WU����cM�=�F�S�CY��fwGt\7��!?��l �{�����2���7)�F��s�=�n�af2��o`��u�C|�/W�`�;V�J�eG�O�CR*�x=P��M?��\ۆs��R�F�\,,Pl�phF'>	qf�7���!#.hB06_&,9��aC�	��ʡR����㾩�-��@����lqNf��6���d�LOs��9/�(���	���?s����P�.��]�����u(D}��A������w�r,�����y�腭R~���z�q+D��a�,���{xSbX���%�L���̶�vZ�6n�/.%5�v�)1_.�p���E#yN HarS�� e�z$	�/�k�����!`Y�\<n�~�"4,��(Y��'�����A��faǂÝA�3���&���Yxw7�6��ȏ�z� >�D��/���Ex��.��]���Q++�n��H]�K�J�`�;�Q&�݃��� �R�aZ�"�rBD�_�SA��䝬�`���RŤ�� >HG�;g�:Ң_�^T�_��R8�q6J����a%^Go�(8Tx������-�²�ߠ��%1�����������p�F���}������Pw	�-ߖFi�ѬE��ݎp�� Ԓ��PD�@@%pj�P�_3�t�k�zy�L�";0�rA�	-�9d%�H(%���Vckǩ���$����<��uBY����?xյ3�m
�:\��YA�5��= N~i)ti�D�]xt2��d4J���%Z'��ʅ��mr|��g��"�\b��#����(.j�dcK�����-���z����	��_��_j��C����a�����׌+5v��W֬���h����~�#�X�[�����J����y��b����W���a^�AF����D��_�1t��D���|�Y/$��饑���A�D]J0�%�ѾD�ډk��FM�r��QḄZٔ3g�k b5����L�k��͇��gY�ͅ���a�������m\9O����ή��0D�wrf
t��m�����v��U�T�i��Xk����햁G/�'��PkX�b��8���eåبTmI$@8�g-�ŭ��$P�G���dS�@��zA)�\˹Ӎ#�^[ʅ��J���}�`�}9n��u��HJ�bl��Og:�����h֜SEa�b�! w��0bB�_|̥ާw{3��x���!�9MNN�Ya�d� �i��t����w�=G�E��!j�U���� T�M���=1�{��U3��gfm�z F`�	�y� [t M�/��ZeD~G�A{�r1�
���j}?���.xޣp����YY�Ț�t��qp�5'�3"�3D\��r��>|����]X#W.��e��DYnR��ͻ�U��ށ�ap�ѷ'�p�@�Wf�1�iT=)ƨ�6�)��V��6F�ƌZ��$S�6Q�O]*6,�eE��\���p:9i��eA��7���Ch	��?��$˕Zia����i�+�y�#��Ds��c��7�9�?�I@;��VT�(�:5�&�� +,�C�O�I]J�/8�ZCګ�m�|+�9��W���r�WhxDo_��M�����񸇎@G�@��8�@a|��vK`��2v�؈g
��$���3��1f�����������_�-�}BJF?�Ω_���Ut/��� �3_v�k��s�eƞ}�y
#<	�Lz��$鐵�G'ѩ�H�UL���".��)5��|�r���
Ѵ��� ��ֿ��1;;�8�N���x{D͆���YWH�fC ���<1�¥����7d�m��뤃�1/:+���ɩL�������gdR{v���rn�������U����^�o(�ڨ>oY@�L�}�'�ޮft�C�&�hs~fP�l�5͉	x!\ݔ�%Q����2�(FA�ǵ��ү��r����VX2�3����W�Nb�H��^��%����`LL��U,�o����i�gA%|�L���ɮx|�~�s#����ТY�w�釮F�}v�A+��Ib�+pts�=��z|�0����]�^��0_w���A�[��q��Yk4�:��p��8�W�Ѓz�*AX�|�E�Eg� C�%�fc�S@�t������-ˀ-�R�O�"����V9���~������ұM^�_�
v��~LDO�a�T����b%����M
��8�ܥbD�c�@d��`C&'���Mv*�"�K�=O1q�"�4��l�����%D>����-vT6v�V}�L0���n������o�IQBT^��=	D£���'��</�9�ﭱ��׽��_�mkd��b�n���FYڠ�Υa��ͷ�'��8aW]�*�5'�o���dnJ�dH��<�?�P����o����G���_�g�;�(�q"xl�7���I�˖�]���#r���h�.���C�`�����������R�*�@ܡeS�Yu`�\?6����J����]+�QZ��>M�M09~\� f��a8c`$͡�U^0�ghkc���N�c����vN�U�������I���͌��z��Z9��m���\i�#�P%�m0jpp�Llŏ���vv��ߓ�N�`�.
�j^2z��%�.ʍ���Mʇ�$S�M�Y�q[L��{�6Y�y�<�Q�s�g[��윸��� ��_��>�C�H�h����r�塇%�z5Hڭ���HB;����E�,\��q'�?�߇,432ʫ�G��;�;w")�U��lg]��d@���X��B�a���1�S�N���jO}/�^�94�1oq�W����	�7�>���Ǔ����#(��_���#$lx ��M�V�B�|���UO�Q�,+b<ѝ����b%X�XN�ܡ/,?��<�o ���i�O<��EdI+����.�ҋܷ;ꏓů?ش�����هyi�s7��c����ut�'�AȂ��붼��D��Ty�W:Ղ#�)w�H\�PZ�Q��B���j*��(���|m��5�}�e� eJKެ����課�J`�=����h�r5r���	�����)�\�%�<����������d�Hf0"VX�Z(���^��b-+��Ml?A!�c����S;�����cK	#K☱���W�{��v�
��O��V/,�!�a��l����þ�c��_HZ
ׄ|���\ONe�6�Ie���D?��sW��2�v^�o.���ĜPM��Y+��X����?�&�����@���RQB��@!�mr���A��>"b�PL�����؃J.
~�^��7�aܣ@5z�����ܙ+p���1���G_�4��	��ܠE0��+��hO��
�]��,�����볪����8�:�ނ��2,�K�*��������6L�S�G;N>�	��ޒ���@a�T�ԋ�43�RW&{�@b�m%��qyq&�]GvvB-���t�\����;3��x�/##D�P��#�v��:;�dM7i����ȯ�a_�j"�	���^�ؚ�Q#��e���`��T�\%XӬ��A��2mL�pNQ�ǁf&�!�G����s�N����ܔ)BijN�M@��)�`&���ӄ���E�N�O�q<@~�`��C7�O�$9e��������B�Cbwt�h�����Mmg�4=%��@@����jT$I�l�e��R����<X�{C���3����m�c�6\�s,�P�>2*�~�ħj���E��.r2�R�D^Q��M��A:����if�y����f]�!���B�N 6cJ��Y�
/T������F��5-p����z���r)��f�{e"��e�ז�d;����h 	z)Ik��\x�e�90�������x	�m�(n2Lw0%�D������&�k{:�x� �[n�a*����3���Lji��K�>^��S�e���d�h%y
c*&|xl�|x��鲺��EsA�-M0�๗�V}}m��R�.�V�������?8�r���֞������j���H���+M՘U'�^��y'�c��j�����}���9y�aX(�� �0��a++x�ז�������Kn_��5�y�|�EO�"�st�ʼ��)�����k�0�%�Q)*�����X���ĀOJ������R��<���A7�^�i�t>Q���>�v�I�l.��N0
����o4>��r�X�l���-rL�PnGjp9p�Q>#�7F;"#�+�>c���Z�7���?���faT��Ro����L��t�^M�83��B��� ��_I�%D�5�J\w|'V��N��z��8OK�Yz/ǜ)`�����6"����pB�]�ڗdq��f�s�l�|.��+���ѠX��>�<V����R�a���)�V��k���<�=����1��.u�RP��{�NU��MZR�y�E1��%�I��/�UG��ς4�eY/i1}�,���ut��Xt<�C���
�Dh-�c�x8B&�?�����/Z���� ��Y��Z[��h)�*ZX������92r�:H�#F��_��]%��JWe������_�&��Z"�Y�G#_wАG�6dv��4�(u
�xˀV�G��ͯQ�������7��� ���-��?�Jzh�[�\��A��q��R�;d8�f�b���$aV퍧�ޔmi��J����JC����~u�0 �ٓ�t:��fc�-��h���R&�(��O���fl9/
��ߎ�V����J��Ll@�Ơä�p�֝ɤ���i���]m*��!�e�s�������#[A��E��v>�֎��{0Ø�uB��<v��Q�-5�*�����X'��O��b����g&�6,����y��7���F��i�α�(�s����_���y��݌[�i�$u~0~��� ���C���*]D���O�:$C%1=��a��P<�O] fӨL�iA�[sB�8  ��9�������!`R��_���;��-"l�'��@7^�g(��q"s�!�?}Hp}�XErr)�}����>��g�i�ׄ-7�| �0l��d޼r�<��+>�"�sc B��;�
,A[OFZ��'���>�~GWrr}���+�<������K�a���F{>q�5�g���vY�78
E���ʾ{�Jh_�d��#n�@��m��/�&ug>&¯���1p�OZ%���+R�Ԝ�Z���($���W�����R6�YQ��ue�i�O�_Oџ0���2��J<������,�k�O�:�5�}�.��攱�A*Z����MD��Z���Gt���ܢ&�lP���d=�U�"6����������'�Gd,�>aˁ(�z��+�T�\�jt��.<d�Dt/m�;߼VC����-!����'��hV�~�<>6�wv'���9�߃���>�r��4�+\�@�s�����[T�c����E�ε�u�5�� �T%{0~�����*�z��q&��:4+����LVXP��=�K�������r���PN����ok	���R:X����K�/��;}��7�)�l�;v�R	A(�%�k
p�8 ���p��%ΘL��l��+u�e�hh�*��#�W8�)�5��jm��h�t^M<=�T�r,�`0ۉiNV+����� R�|<cR�7Z�z(^�l�����t?n��%y�%�| ����W�k�N
]����3�h�3���J�"7�U\p������/@x�*�o4X�J�	�M�1nL�N$0�&#(ɶ)g���iU�(�v�{-K�6�䜵���X�����ɀIo;,���	{6��(��U��D>&.��֩����gs����^'���%-� �U��m��E��x�}tQ']�5s�FMI����:%���4p8J��� �Xւ���S�h%u��ڸ=��d
+`R,���K�D��zy�K�l<͌�;'4���0II�k��[��Ә��������{�]&x�����i@��,]��~���@���0�ࢼD�^V|~��;�����%W\=�yZ^4�hyܸ��)̹��L�r7Z��x�	��Ы�\��/��cS�����F������F�]�]����1�2A8�Y�x���z=�� g��c ��ݲ{��{W���:��	����\�sr��c#"	ez��E��r��A�׆Mػ�0��m�2rf��"����ln<ۻe�"����x0`�^���, {]ߡf�K�4�r�֜��{ֳ�� EZX]�˵��21�M�*�;��&	ۦ�5���݆$�<��j�$�{Ax����]���
�\JkZC�-��paEKs�?A#� f�U�"�xD�Gؾ�I9�H(UfD]HG	��_�aD�DL8x˽u�pG磯]۩ *B�$:Gg:L��a:���*3h�����B���Fv,�5�A"��KL]a�Jp��dqb=Vu9ΫE��2#�� 
�6={�cCCR7U�nE�ǋ�3���&�X�k*���\�S{��ul�s�����d���ﻀ�U�ٍ��j	wC��{�((��4�$H��/ʽL�kնB�^������ �*I��'1ۡO^B�L���7 f�:KS@� W�^�ӔR���[MxY�Jq@��ɥ�ָpt)/t�e<���W/M���^K#���ܯ�͓��+%��&r5�Yl�����f?ң�c��`Y�,.l&X.����u/�B.��4�W��.�,.�F����c��ܒ��`�-w�n�����2{(8Z�^�_�r���W[�����O �[:C5� ��n�jٻ���R���P���.��2uX�D�Zv��ͫ����������Ix���4�f��񉳳H\���̏��e���-��e:��'�wU���tı":��E-�b��x1������?���<�p�w�j��b-��Il��Q�ͧ��⇛�~v�{���]r�o̧�r�x >D=զ��7�l��� ��y���ަ ƒ���M����O����J�g\��oh-�<#Dr��N��oe/�/�\z͵���-d�%_M��6><��N��x�g-�R'y{r�«�dM�}��ʉ���|C��>���h�B���ȹk�����j�J&OMS�E���1�TB!��6m� ���q_P��t�9�w��Z�q�[�6�ϋ��;���KCv������X���G'��nOq aۦ�pց�8�HP!���<Ec�uG{;�jvw��̝9a2��# ��>w��ZocGV
E��s���#u�f��<�E�$��I�kV\>ܥ�/��қ�)/���o
�t�y�݈b���qT�}Ųmif�d��ȯi��=�8׉X[۟��î�^
߳"á|���䐼�N���$|㍡j�o�p]�A�������m��n�zHA<�N��U; �y��� �y��j2�\���{�q{[Q��GH/�w�e�})D�9o�3�I^�(�;o��@}�4f�2�
NO���$7[�jաFz�"(��"+�>��&So�l�U0#�?-�=y^�®a?z ZiG53=�yꫢCky܈�\d7,T����	O��x�� (�ݠ8�7I �/TKb�UOQ�G�����,�wi�<�;eS���R�(r�ɖ6}v@�Ez�?�N���a�Sh�IB��0�C�oѮ�*�B��(��$]!�\B���)��.��J�=�VI�8�B��X�����۟����\���[����ȭ��4D�7V�AY����Y���ᷰ�����`�j�Nd4���[�eP��g��3�D�N0�1;b	�j��.���P������<����Vwu�`��k����^9�g�)�F���k �L�z@h6����u~+ж+a��s���\���tK�z��[�^~����6�(�+�e�޸��r�G	K(�ۦȣAZ��d#+:,q�?�����sIL#�C����q0�TM]H�%C��8D�ޓٱ�2�Ak�
{��1�"�ڣ��LB�������`e�u��S���������d)�Ŋ]�tɅ��uR
���y7t�)��A���	+�m��$a��V{\����~UNu���
��>n���l�B���c�����2?�JC;6\ԙZe���&#yv�!��0O�`_��I�6y��k�3�uz,��H�>&��N'���H�|ۃ@�-J�����9��7Am�i��m�������8��Eeʱ(I&JE(*}QZ!�a����
���
}�&`����u�V��ynE�����cR��h���6�M�aʵH���R��X��u�Tֲ>�ć8���k@�ȥ*�6�R���~�#T0����Њ�R;��ȸ8yG���k�u˸M�]�!��`��v����>�`4-sU\/{,��f�.1��<p��'����zn���,b��ԁ��{���y?�.{_����	�����M� ��5�RY� �͓��~� =ly�ޘO	H��[�����<�<��ᵪ�-�Ea�8G�&���ޘ̂���¨:4}~;�{T�=˽Х�KR�c��<���+{��o�|W�1��H@K��~��Fך��?���k��]e}6�H
���i�1�~fS��~��n�
�nR����>��q�ĸ�ƹ��
O����&9��@|�N>��9Ӄ�t�x�n`|`���t�<�`�T��*�D���/BN΋��Nt[�.2�N��@u�9�&���Q��oMn�lT�L�{叹Peo,�]��	ԑ1!�T��V�Q�c��*� �mz3k5��Va�">f7��Z�� �ZH���+��$�%)��@&>!�9|@�-���.H���phF��~�	߬|���a��i^N�>K�Qo��0aL���;��@�}�[�B��r2�HBUB[�����e�vQ�u,����p}�9����[ȓk�thp*�CYtʦ͝�LJ99����5��l�
���Z�:�jkr�l�\�\�{=哄Q�]ҹ�Z`�td���&Lfyp�[�4�\��һk�,�S�L^tY�����S�����7bB��N ��zj��3=�ؼ��'� �r�R�!���_�V�eӥn`���4�9��
���H��r�[�%چr�P�/��J؂���R�$G#�h\(M�vTEq�bf��w����d$XN�%LB�*�Z�Sr�{> ~�b^	)1��q�K���lt��V�[��
�Ǧ�,���X��:��M%d�a�PS'o�M�W�*a|G�V�MZ���i���k�dY��yA�+�z$9{G <����?m�0v���ْ��]Su��;	j��\��k'F؟�j��̓8D1�	����8�t�q�گ�H�����R��V7�����'3L���4o��v��V`���>�urŒ��3a���|�܅Ό}s꠸(��\�>c^G�49�iF���nC��( ���#��u�,G阡�Ӕ����ga[�4�ʴT�*�aA��-��`V��H>K.1�1�i5���/�E����tD>2�4 ��ل�JP'Qpw��W�Q<e�)Zu��s�*��H��޵�)kA�ٸ{�t�qS�mk�m1����;xҩ�M�j�$2�]�N��M3
�ˆJo�[*��i3��|�
B���X�=R7���M-~��t�\�"��g�+��8~:��Q=�3-��}I�#1p�u�@M0Q�͍T�5�AUދ�wU��SbM��*�AiGy�}]��i'7�塆�*~�Ȋf<)]��������7�3w�G��Ǖ����R4�8��u7����J��<tEe�)��8Q�?����R +�j�>���ރ�Md�-��8�� �/?L�ߠ�p{�q����W T�z���V��i�)�st�IEP'��߲�R��o}��/#7ѣ[J�YCX���R����π̠��_8)hXx�9���pL���c���u���H�3#�0B����H��24!����$���t�.�/1�<��Q�=�H&5��bE]w�����(�xC�^���
�FW�<>NF��g��U�'�,�IO=�����uc)L*2��������?�4ҥ�m��T���X��_]b?��@T��x�=�Q��]C���n�7`�K��:#T�f�&1��.�0Zm�pD��ږ� �J��S����c�q�b"���L��'��;�X5|��4�l�w�e�3���Nb�Ç�C�C����t��`'�Ǜ��+�����������~�:�;K��o����������4/�������x>u�ÏA����Dn�76�C1���u��:�,���\<�]�:\��a4���v��JׁMu^L%��s匠�)���ɍ�%If�DQ��2k�ܣv�baP�+S����!o�[��W:����,��n��ٶG�M b+�±8�.立_%E�=9�#z_6e�^^�V�y�@�0���܎5��|�.|h�[�	�r���N���ki���;���7�3���f���ΰ�fv�wh1|��`��bR܄o��}g�c�2Ĳ��!>��W7}��g�(S�`;W�J5�[���Q�n�W��7�{Q��(�}UI���%�*����R�NjR9�|ݐ~P5&mǷI�a4��N��9����C/���@u�#����������q���1�n�B*kI&|�;�[�Vr^��c��XCV���]�ݣ@��|�o]��"�c�a��t�DZ�Fi��Б�����u�<�NQD���X���۽�B��("��bX<?��p�����!��p#�q���)��($Q ��q�g�a� Ord{o.,�%mp�j���wxB1�i�*.G�m_�Z��F�k�D�8�ƈ�c�C=�C��) �q?����N~:5��tC�eL�W%��H"!��g�����%@av@;:�4�uQ�KL�M���L�~�r_^cb6���EP�D�_/D%�Hl����*���wPT������j�(uW!�\�I��h��[	=��:|+��ڎõ����T���²_�ŋ|3]t]f 8�����/p�ʶo�������� ��A%�U�݊P�?f����[��L� �52���y'���VX�(9�{X��A��U�4�;� ��@N�s�ho~���-о����pGL��Q��M셁�=3<U�j�@�1����Ɍ.��l,�r7MW�ً��U
��7�q�mD��RLB���y4�D@-N�dWJ�0��X���Ab����'�� �'���cJqF�(X�KFx��<�����@@�H~����߰nڟ���Q\c�z�ʆ�
f4;��]�u�ˍ#���v� #��/&��z�֫��=�g�ۍ��
��Ŋ���ԅC�^e�rE9B�sF>ɌmI�yy��5s���Y�H-|��OK	/	)de��G�sD�r����e��L��(����[��ǞʄE��y*sy��K����y�?�i\|��� �
�F��%j�9���X�}�! �7��c�$F���E���[W�R���|�W}+��S����Ť�Z��vCN���WE��Q>8OPqhV�I(�ɭR;�;���g4�]�5вA4��:���i�o��T2��ds㛰HW� �r��{@�Z�-ѧ���e������\9�Q@�d\[��Fk8� Ϛ^�G7%�[8���ܴ]�+/~#�|+A�5��!��.��7E<Tn���M����Wt���C�{��[��?�\�D @ؕ�|�9Y��_.�wZOk��G� %�f�ۨ��LHt�Fc�������
yri$L
�HP��*H����}ꦈ�)�Ǣ�;QGv�'͛�jnʁ���`�I�1uAԂ��@�g�
��L2=�´��!	?qNI�o ���Y��S���!A+;>���	�����E(���Ʒ��M���X�r83M]�D��B�26�����_l�٢r�UdJs�a��,2X!A8��q�"�M��$��S��P=dp
����!<b���EV�����
K�$
�n����s�@�B)f�X#r����m�}�4'���R~k��1��š����y0;�0e%��y8����e�/:�F`�|	�f�Y_\P�	��"k8q�#o �OK�tn��KH�� #M�8qo�ry�+����(E=�f��g�=�f^�u�K�XHjݢz���'FA��ad����m����D�'7o>����%�{w��u�P�Gq�+#���@o9��5�j�v�-U5,���	�Ҵ�l�JA��6�y s�ua�q�U�Y�<������X��@2q�K����_W������4����J�̮_|�{S�p0\�ӆ���_�>�k~�$R�>�д�Q��˽6�r��ZAo?>���X45~�M��<��P@͙�mI=�npGw�L}oh"�"�㕅�L�z����&k�]�Y $��z1v"�x�&=A}�����
�:=U�]9
�_`ץ]���<Ǜ�Ibj(bv� ����ub�s\������|[��`ט~l���{h�ldiQ�i�������J]��D{oDic��}��sf�9w/'ɼ����[�o��]��:}�,�Ԟ�3��c���C�1)L��QעΒqՁ��	���^wG'�gS�{׫�Y��\Y����
3M�D������23tǌS$b^��x�Q�����|թ�Z���a�c~D�Y�?������gc��f"�	w�&q#�ݤ��7McV��A��J=OI�E��{h#�Y#cA�Lcl &�]|^y�L~H����*������+(���Ք�ㆳ!�`��kw�8s�`/��~sr��쩮���MI�V���yEBT	d�LI7F\�秽.�Z͆3��-[y���6t� eE-G,���3A��>T��J�v��U�� �7Ս�T�p�N
h?$B.͕������:��a̤-��k��P���sG��˸�_4�b
��7�qۤ!(��:�*��E�۽v��z���܅[�Z�!A��!���l]C�u����o�W�g:_zU8����حZq�.��-Ǝ�=�|��G�le���o$��%��EB}0�=_R3t��߾	E�T*^zo� vc'2�=//t#��� ȸ�G�qi��{w����䆞D*2F�/�.�ǔ�|-�K����ʪ�x
YbvwN�����W����1�qw��<�N������ҕצ�_e�5�p.�rצ���)�;S�8�����}�Cgͼot��,�VX*��A�d��]?Zfe^14�"�;'K��ސB�d]h�+mg?�w�����H�Y�l�'�&c�'���?�f� ���MX�tD�@�����~�8�(�n���:���C	n�	սo�#{0	�'`wG*�>��&��>�2I�;��ɢ,C:f�%�g�[�j�哘\�����}�8�N���U���~#���O�h>��/F�ghp79,�gQ&�SH�o;J2�t�@��q����f��<b)�|Ab�}��W4:m�����>��LMX�3>jэ�u8VA�I_Ű���6�""�}G.K�(�6$V8BC*�!(����*�t8k����anS��A5�>5#�o��i\��_-t�L����t��Om�QU�Ne�
��V��L����D&��	�V\�����ڸ�,�F�4,n�����K���I�C��Z�,FX������j�ų�3B�7��� &�/v����cE�e�u� K�$N��W?*�-�K�0u���!u�����8�W-��R��ٿWM�y%���!�.��������a�M����Վ�^��?���fpi������Y�]��7�Ej-;�$���T���$�3��!w`�Ag6_҈q�)h��u�g6��o�;Ɩ�����h�Ma`���>���C2��M�|���erY+��
����feb��Bő
��i]=�����&�+q�bs����C&-цO(�|����!!��]��OT��S!C����1I��m�1#"��!L�m51۫�����Kh�c2�%qV'Zc���!��<ο�iq� �ⴟ��`C�����7[uMb@X��:�;�I�����D#�J �Ԯ>	l���,ĺ�1���M�
>d��0���S3���ȥ��6���Y%�Z��r�u��	�C�%2��In')_��$@+�Q��� ��z)b�/j��e�~�w�nPZg^�c�c׿��e3�l~gŁ�P9�3鮞����49DTD��6�����0mV4J����5�#�+D�"ܳ����K���\ �}­n�)��-����=<�C ���b�:nWsi�0�@HDX�zȅ|��S��JZm�����S��_$��mf�*�>��������6IR�yJ!�r���W�6�y�щt��ڎ�����mT'����w�=�������t��z.���!f:���P!�����%G�@�m�Hp�l,�q�ب�Z�0�i8O���@�I��G�{o���7����V�����&JP����Cl~�k�5�C��� 
�+����WuC�q-Q�_���ܻ������ϴ����P�o8!�������׍*g��A{Ⱦ���em"����̆��u�T�����QO�X��znn�$x�=�z�o]'�wI�C����uξ1<yL�����>~�pr/��B)[�12A��D�^�=*<�����T�l��$�?u�5'On��b�����4�S C2I�T.6w�#���Vc3 kl�j���ޙ��4�:lZǸZ
,�m�3�. *iݚ�0�w��9�`��K9fC��%�D�$���zJ���;���+X6�b,����*�o��3�j����}�l��F؝��6H�~(����u�#~�/�Y)��Le�X�d���򲯝A����՝������bt��-����ҶP��\	��Ҭ��
��@J�5�2>&��$���O0ub��X}��ν]~�l�1���^�d�SLj��`�.�$a� �k��>�FS�(w;��`��7�%��9&T4 �Ҭ+�j�����Д�a�3�;S��{+c;���zN@8���b��E8��%�^>a�}��`<_�ר���%Ԥy��3V1�DCKV�d ��OY~�>Q!cx���.��/+]�G�1@B��������U�SM*V4SU��H� u�|ö)�5i�-��vI(�����}�B�~%�0~G��
��f{�%5^��;����K���k�y�$����5�����rQ,����鸦ng�*��^) E�[ �K=��bPy���دY�P̛�>*?�� Q���x�m�0��.�6/��܎X�`�ԝ���ϱ�QgH�.�)�f4��VW�&�He�̙6c��N�'�m�w�WasU}��O��A�ӻ�}B���4��f��t��0&8�W~�ZVِ7�c�a��&$6�*_9��4_.�o�b.�����r�b��1=u�sK��*�c�&9b�8`�!�w;jY�qS�ͧ9"���~�5��6E?��]�%׶��'F}��U�4��񏌔�p�8����>TJ��F�TL���$�X:�py�)�U�7��|3����->-/+�F~e����l�k�ٹ��Õ;=S�H*�\��Xbm��ag���7�
>S�j������~��<R�UO�J>T����z����~�q���$,m.���l��v[��;�� �����:#�;�"ߗN��sˑ�R��䃿�������aS�9S&������h� U};01�ߡq�˳�oc��R�.��������'[�Q��x¿9Q@��{aﲐ�!��Y����{ֶ�h���Ҵ%�5��q�����9'	"-���ѡ�	X\_v���ؾVK�)\g��i����αy���O^�.M��Ĺ̓�3�J�Av�o�?{�+����J1ؼ���LLb@Rk���Dà��������hԿE���nۖI������1P�kc`$wR����.�3O˺	���Y�'Z���]�f��=c��+?��W��I�͢�^��[T�=�������}y�}=C�ݯ9�����WM?�epm_��3��G-�d��>K�X�֑�?^�
�a�4
.�R�l��uh)���M}(7�O�_!��N�GD���F���	x���j�����B&���=*��R�<���p �=���b7��V�U3%fܦ�X/�i�#�:{�5�Z�� ��G�m������4*�Z����m�ԝ���B��oq��tƕtV�6Zl���EU+����Aԏ'L@��IrO�x~	���]�1���7�ǋS�U�j/�����\��.�"T��2��*��*�&���:
zn7��ձz�������V}C ����^Le����S�к�9D���`��dy�n6���OO������8�t�[���������"�{��{�],�t!����@䲏U�8ޥ5��yV�=8���:a��#$H�O�S�O��Y��(2|2��M�=���ymϳJ���E�Z9�R��H��L`��/�R`w��w�;����v?�&J�r��J��."{F��~
"'�5b��}l��E��N��,�LARo����=���]��ؓ�}
^p�K���p��=~�(p��e:+O��F�?�=�'@/�*�NS�&�G����n�XjC_�~p]���"��͏Wr#x�m�`>�uԈ��A��j\�E�'�c3tΕ�3����M�T^ST�l�*k��u�T��Μ�׿�]��ܬM�@(;QL�[~���l�3��C��hE���{��|�GS��m4�a� (3�V��i��Ѭ��"�"b�0I��|��C�i��ܓ�}ťi�t�A<�گ�CQ���X���ðb�CVi��G��hO��c�}&˾�4�!1��c_��<�Mm�~���?��9���r��mL�~ӕ�b:RQ~�Ui$�n����%�eQRƏ�W7z�}��!s��Y�.�a~�P- þ�L��Q'��?m�f��`I���)�����=��C"v#]v.�e��25��dZ�ѫh�f�łBa ���P��v?,j��p�C���l��QHB=0y
+�?�`��ׄ����pU��+�D�ة�� �/�p�{(+d�}S�Äv�In91=���<�x�brk�I�M���r� &�H�A���(Kp�N�h�������� ���H��Os:��O�2���Џª�����U��8�o�>�����p��~L<ߕ`�_�ZYHî�ۓ� 5��юW�����\�i��K��a�G*td�'e�Xb���,�P�3�K���ഖ`�%*�3(�j���"�<�z37WC����`�I)�[a7��b�ȃ}��a}��s��qߪ��1�Ӿ������g���?��ZX��(����=�
�����B�I�:<Sv��ט����ֻ��l�s\cnR�E���R�$�q �TM����N_#p���b9E�@`DF�,Z��.kEH�P[uA4Z��E	�Q��Ԛ���`<e�տ��'�}��RC9˷��.	ķ��b4�u�� ̲���i�W���`\t���X��B�ѭ�ū|��h�@LI�7P����/����2�3���kx���S�i��5z��_�R�>�z�y(�aO�44�oŝ�|�~pW��x�9���@%�T�'/�b�fbS�Ʌ�܌P�_u��䇒�i��뇊P�w�^���"9�=l5���[�wr��S��I�<
�?���G� Y\U-��p�e�1��?h�K���op��K��qp�(}�
[�z��k�&��m��z�T�]�e��	<�&��uSSG_:�)�b4��x�z[aݒ�u;�����32i�ݹ��%�A�u��_	�dXc�o�f;�T\`�E����qDYVr�v-5�����2�����q�cD�����>�O�za�s�{˙�(�
c�(��]���v1"M�nӨ��ǻS��2Dn�<�V���X�u@JS�YSd��&�>~�����}Z[�%�
��2J=�����(1��>�0�±���9叵*���X&��z'��[��H!E�1䛭�w��kh���{u�v�|q¢�@���Z���G�<�Ӈ���� �� z[*�I�d�\7'mh�Yy�����y����k̃aa��w��e�8�R�(w�28>C�nD��=5�>�}��F����C���R5�ձж�9.
�C�*#��v|��-&���@�m%3.:Dq���Y��ɿ�s�:��Н$�J�v ��i>�0Ny��,6J�6תf	4d!I�N|g<��پ��B�:��P�-.GO>y��ԑ��崙�8��.�}��}V��`�A�80��ˌqیi����&QF�~�49`G?�W5Ies�ɺ�'�_
Mfj��JaYT�� OR<-݋P5�1O�,3�U���BZv��n�N�k0�?u��A٤!Z-�6�R�����S�#�l�`�6�)�GT����g�Gmi$g;/f��@���N�ˇ��X��i���3�k8|��!z�/s��7+e���� ��J\u���?`����ǟg�n��N��@ܸL~�f�M1��ޢ5�k5�Q�^�D0��^��uwj��R���bY9���������4�G�Є8z߄̈���5\��i�;u��ۚ�A���(�f�֤qn�4'���('�0,�@>;�:�?�����f��Ë
/��!�Wf�r�޹�"`/��hh��c��`�f�k��l}�ws�f�h�R|��*2�p�q%�7/�����n�=�	�u����]4�}�DLlܚ����~
-G���6ד/���@��x ��}�)p�Dn������U4�-�4]�{�Kq5�q,f�]+�Z|.��\{~��U�>	�Ƀ:&�1����y��;{m`��������"[l���T��P�>[�<�dl��_<������/!v��<��y���k������HC�JB!��z��Y~2ۃ�b�����blS�(�}r+�ڈ��s#�ѭ���ׯ%2�� >��`8ײT7:���f<�}|<$��Gۋ����]λ\e���8��xn�
��"�^���"я��.X�v��g�)<g�n�`�"��P����'ZPQ0&�kͼU��W\4�����4˃�q1����0A\|ڨ%�ө+���7�g��O8��F�|y�����ȁ��r�(��a�՗��5�Sx4Ck��k?Fc��x�D�W�t[��ț9{h�'�J�VQ���� G��Uq����)�����	0�H���M68ƻC�i�j�$���G�����h��7�c�d�v�m'��>�<39E��a%D�*�:�ǃٍ����h�q���U�BSZ2k��f���6�E���{�**T�Gl-��!HD�z���	'��2��;{hC�ݡ�AU_���{���MzX3��fM�ne�0�����5O�X3eMb�a�	=�$G���o�P�]��.��)����J�a}Q����3�@�	�T��8��Uj;�L�@GaJAq⤱���X |�A�É��Ǹ���\5�c+���wpy
�J,��n��0v/OV�{�=j�u��<�e�䝀%b29�c;���K�Ԩ<�+$�^�#P`�)��/ɍ���lq,��������[��2Q�w��qU11a�s>��h;'�����d� �Ⓓ�'�q���o��X�ֳn0������a�<0�1U�
�,|��L��uv�j�
,���b�%i�nU��Ok�0&"��ػu�A���:ً9Վ�y�A�m��*�=��+��u�T���$�8w���1u� ��q&20���3�ƫ�&��D}Jٟ�a.��� �W+���t����>���伍5��a�y�e�io���.���O-�+
���}����U���]�X`wV��j����?Ji���"|��5y��I���m������������-Ipl!��vj�&�¸�e��[�{�DDM=0y*Y�	��4��ؖUb"x>6�=�G����K!UK����a�/�9,W��S�ٺ��f�F�`:�6���Ra8/�x�}͑�uS�#58H<�����l�9_C�2x��8���[:z7F�x���+Mۙ���*����:w��evc�ͬ<��n�ܓ{����	*#�����Y��+� O�<%�E�D"�
�.O=nƃX���R�M%����ˏ�E"�T�ѯ�@�ܟ ;��F68����7��dvL���.��?,�����YC�{�̆V�G�=-LjB�I��-R{`jZ�R؞/�%�Y�����Z�"��(S�s���C	�����2'��g$uA����;���:偻.rm��K:�N���/�%|��tE�B*޳�.�vf�z#��vb�-z��*+��?��%�D�'D1�t��x���w��AM�Y�pc~�8��ǭT!��ut��B!�˭ę?�x��&�*_�ʡ���h�J�X�%���#g��*Z\�&�.N �; ���u|f񙚩���:����A��i
[AVf��
�V��^b�JA���h_�.�h�ч���!��Tr�̾��g�C)��'���y��L��ߩ�>J��_�G*�Z���跬5z�0x64d�C=��.<2;�M�^k���'Q�g9a`mݎ���5��_�p^��Q{&-�����b�v%���U�N	{׼��+W�r�#n�ɟ��Šg���}�mψ>�@��*���ͮ3�Ǔ	� SwZΜ8��,p�4mPb�	��<�ɇ0���;��=]ԫ*���3OEK��T�g�*�Q��&�JU�e���}M��t}�M��j��i?���Pd ��1��q��D�v�Y�9ޤ��	Q5�/̓m���Xo�E��D�n@��b��~䢉�\ D1�Z��)|S��i��^�ß���2��FJy{��u�2� ����G>0�����".���P��c��@9+6T)���,��M����2Y�l��yP�o%�|u$:�^���x�s$�9��CSBK�T��A�W�[p(4����T�6(���j2�ֹրT�`Z|�94`����N�ۭ�"`�()?|p� ��d�f`nӟ.�S���vy�`��9�?5'6V"el�jG�s{�N� ׈�$�jU����եb��V7p�Q2)��੡���w/�Ǎ{%��JZ��BY{�Ts�`�[���Iz�o���y�0��g�n�|�z�L~_%�~-�J�Y�~$��I��uo#�>�q�W�>��I}

N��VX����4q%OmR���&�p�j��2�(���P�"��T��	��C�y�{�a�q�s��ټV[�{p�S���
�R�$��^7P��������yo�S(?�G�^��s[��r7�I��X�-��i@�i����f!��c��H邚�q��i�d��А'i�BH�� U�wś���$��sbF\7T_NkzZ��b��5�ԒO��.�����Ǡ��Ϲ����
����*�����j��m��||i5����8����
'�*��'�	�	���=����qf�N7��D�o��JԾMl8�Şj7֠C�2�|�r6���$�
���)9Ķ���r����]�2�`lc�u�5ZƋĥ���^_�����9��nc��p(��޾��@{Tte�\n`v�.�l=�{-0���2+����İm`؆U��:��S.���.-���fs��Z�a�D����afy���^!�!>�駝�3(^٤��;���o������ʱ����)�L��K���r)�P�4}-
�d�P���=�>hZ�V3���(�2^�#.��'�����V���~| l5#�e��DQ  �/ ԅE�k�����w>?X'��#�|g��H� ӵ�� wl�%sV�;�T����@S�is�n][&�l�}]Lw�� `�&�,NJtxq��$(_�k�կ�h��']]�Mh�0���J�)��b��R�>��ؙ���c������( f�;�Z�\�R�؃�zjL� �9h=u.���9M���ܢ��
8z�f'}��(Z}��L�{s��@��)�qD������p�v��:N9�W"���o�a"�{�@�L�����V��ç�H���Ml7K�����~h?�&$�۶}�VPm"��5	x����{������������~��r�F��4�%|���&����oSL}yK�e�� ��z�3Ja&|7�����Ag�f񨢒�%��n�3#2si~ES����sP�����\�1N*��`����"6�������L&��QO#���;�>�IB�yW����0�6�z��S��:<-(�̄�hڪ�Y��ϬD�0X��Ծ�y�P\��5�����w��2鶴�`�m�R�akbS�t
���-\�)6���if'�yGZ���;���KY���Ⰵ%E��}r��N�l�D����g "a������^�Ak�_m�^Q!�Q6,��7S��kh���ZDz��0��p=��f��������$I^���I�d���
��[2[٘��dI�;�=ۀ����!��5���Cg��_�HJ�}l-ַ���K# ��3�'���WS�<�%De�Ӓ�%�@�^�!�B,��_.�^)*������wC�TC!���8��=ޅ��طFbA�!U��o�@�p'�D=���o�%��0wO�����`�ģ� 񌏲pK?а9��n2�Yߦ'� 0!}c�hVr鬐w1���xd�(в��~9��L���%�V�+�ŜHN���P
zO-�y��v�M|\��Q�$x+?���ς*p+mC,A"A�ݢo�����epg�yNK���9Ҩ�gDh0�V�������.�`�	��B��8 ���Q���iq}p�!�Xd���wa�G����ގ<q����$
�h" �/�9��!�x6��P�X Ǯ�jE�W��M5�`!�^H~�r��tP��-��6Q������G�����O4��Z�Ს�}���s���*vYH)��<����a�u��C�����$�9�R��_�"s�1���J.��\>׆�����q�V+�B(�v��! �mfu��(�oX"e�RN'jd�ҚCq�eaޟ�����Ռ�lt�9��Z|�g,�����'>��y�I0�p5�Vr2�?��Ho��x�߲�.C1�Fl�_{$@�Pw�����튟VG7O����<��8�:��{��ӗf�-�f��X�?S�����"3#���$Ĵ�q����+�ۙ�W�3�,���/T��jmݭ��(uW����.�T��wJ?O�J��g�Z��^ �i�Uh���chB��Ԉ�0��#M8�Co�sx�yX$�#$L�p�:2�'��6J��ƺ�|�O`��U�K�ΛXؓ�����ᨖ�I��^D�[(�%
iQ�mS���N+��b1Q�QK�0��C@�O�'��b�/8ГzXi0q�>k�g>:&���_4�h�o�dUw8; ��f�d������G�O1io����ڿ=�oP�YXH�C%��r2��__g�uO���wO�7v`�P|T�m�l�1���X(�6b���ku�ͯ�r�X���w.7�x!�;��U�I4���off\SG�=�=�^!(�(�hN_�OYJwZ�JX�u��k;*��՗��{Zp�7��a�Y���k�&�5��0���dD4�����^u���89�@�s\-��I)$I�Sm�\�)=�#�+��Z�w߫��5�I��������+��U�ݎ���n�3
�����fh�B�]o�Rl���S>������	ג���g4k�-��!D_�˜�����)�M7���؁���RJ�4X�2��&9F�c�h�R���/��Q1u4CQq!���"�?�K�͹�`�������zE(ߓ���8.���fr���kH����6d���1��Z�����l�F�W�q�猺SDe�������<�N�`o��ؽ θ2�d1��{��Wڸ}�B�"�~gW=a��.n�&mr�FM;�V�G�����$��|qA��
@S;(�@�.��;�2�s�m���	�^n�@^�R�#?�M?��U�Q���^A<ǯ����.0e��ŕN=���A�0�lQ�=F�$-��E��Fм1���[���c�A<p�LRҾP���+L�1a���|���< ��Q��#���P��H�ʤ�Xw-W!O�*�q���`>V�d�@^�SZ99R[�����]u�<���.��W!F�B�Tp�M.SH����ˑ�o嫎��Ru�a������hh#ݞ^�l�A��fO(�'rW����A��t]z
ܯzQ�n�Zx����Pt0 UDt��V��w]Ϧx #��Ky=�ωK���sTy��3�4W�Ң^u�p��M��s�R������5M:�0o2$Z[b�eXbj��Ə�Tv�F��_!΃��i�C�����t���|�C
>D��8/Ԃ;6]Ȇ����?�妋�|��c���akR4;M�W ��ۍ�"&ɢ�Y�-N�-Q�\oΠ�I��rӯrpM��-7����1������J5\c�+-�p�o��;�k ���a9z�Cv������U�;s(���E��t�A0I���U��qh�ǘgz���������My�e�'����	�$"t5 e/�c`��[��6�����UL{��Y�3옔��l��pHp��v�{�g!O, ULX!��z���>�1�j9�b&o\W
��X��`�t�����!1lI��eZ�� k7��tE2xW׬G�|��>�C0���x1�Z�-/lG�r(=uELJ�5��[�8&��/�k��a�{s.Ѝ��-���g%kd�<k�N-�X_�"���Z��a��L��4a4P���&ӗ�tT��dĖ ���=amtG�G�;o�G>YQar��I,c	���i���5Z�6�������� ����I���a�S M���^4}Ї�����$4��&nm�[�9+�cKc�-�.���c8��y�,t�
�T3�o@XUO�m�b8u9��'�t�$����;O��pp�p` ns�)�ْ�sm\ 21xzدKV��N��@5��oA��y��v$�ŀ)��d̐�Wϲ���h�1�JB�����֍Уb>`�!��1h�%�q*Ӿ��&�&�)�������a�QA�]�u�wW3"X�"���VU�ɥ<i�v�U'Z<���=4�D�#��<��\p� �|�IK}���P[6[S%��ݒC ���S��o�Ʌ뿁\IF���󩬸�PN��Z����mᚹ�,䦑�6�a�,���uw)��;`�rچG)/��VC��
{����q��؟6�4v��u����>v7o/*h�j�7�FH�֞�� �j�+ݖe�ZvYs��(℺O�>_�6Y:~�Q��kf�"+��H\Fۭ�]� @���Mi#��_��j7[PJ��⦸f2�Ϯ���ިZ��2Q4��ת�_���]���ٮ��@��$ￂ]����4�z�(_����R�S�:�l���O+
q��D�g�Y&��O�O"J����L2�5�5d]��~^ �B���D.�	� ��ς)�@��R���)�;�Z"L�a$n����e�5�k�s�&;�֤WL�Z����e3a�/�*�h�4�T�=u까����f�K�	^�@%6��
(�u��h.�F�,�^ܛc��>����]��_C�2i�Z�<o���Ge�?���ǀx�6%�B�t#꜄��4 9�q��~�f�ltgc��d��(��� ��s�8c)��	��l/�;�vu���=sJ����9�\k��L��T���ˇ�'fR��H�~@�ː ٯg#�>B��ޤ����*Tn���|�T�Q��Ci����CF����^����T"thwI�E
�U�0#egB���
,�u�a@P3r�|VT@̍J�Z��
�MD��b�a�9���:�tVO����P�#A��%�*+�F��ݣ#�p��&�&$���41qso���*'���<\�`��eyͺ��Q�&	�y(��t0.k���r!V�r�l�䄟�6i���%K��FCʬ
��,�;:z;X�0�3FG�_*��;p4��W<��)^KjRԹ��^;���F����0@�I��M\��������E3/�qIT�FȨ��7�]�}�u�_���5ɀf���%ߖ�R�Q�m�V8�]HŶX-8��WA�g��{�w�^p.��K�]��>;c�Z��?"���n�*ޓ���}�T8�T(�CEDh�jЛǼu��HBY�H����vb�{b��ߟ�ѥ�� ?R��A�6@�,X��vW�~"�SY�J_��L����R�\5���_xx��'�R.��ޞ<$Ґٽ�{w�X=r�m��N��|#�-ԅ��x��v����Ӱ �� K�L�7^t�v�N?s'Q�}7�3��S�\��۵�i��_��w*8��g�Y?��ۖ7�E���A��Fl-?2�I��q~�斘]�88C��`����R�yٕ�R7��*�K�c��D�E:�D�#m�%yW���R���-0n�F�������&�2���R�n�}�-<�s��������c��j���BLSV.O>��(e.̹�E��9;����{����0��\~F�y7bNng���y��MƼ���C���w� �U*+��#���3};��
z���9�����������V��g���B�O[Y����"{~�H�P�'�3��k|q��nY20�=JQ8x���{������t�ass�K�xX����ȃic��f؈fp�_�$h�D$������J ��DZ��۫AI���y��~���Ț��<SͰQ!��d�(��^�0Q�G{/�&�4b�V`^��
�*���<M���϶iL���h⊛ӫ��V}x��ﳬ\[0���j�/�]�#���jK��cH8�o%خ��ÄnS��������0�j�1�!��v]����B �ۭ��GW�K1b�N����P�_|:82�"��͕L��Cރ3Q[e��G��84��3��W�|�%'N�G9�W��6�b5O~+%Z�@y�����a���%��U����Z��]��ܠҹ���'��v��!����=�rC@�/��.m��c������|�Y~��[t?��SR6���9�xA�I�rk%(�Օ�r�b��Ҭ��7�3�s�]@����Mؑrй�s"y
DK.���1~S��M^��sD7��8��0/�7Ӎ��ea+��b�`�a��~J�
�S���b��8��Ryd(�I�tzE'Q����IG!��HQj1��HR�U(uܪI��0�/��[$�xҲ�/֣�}`�F�@���=���۳,J�s�ԙ���h^��W����� �y-&&��s| �_O�P�w�q��������m]ŇwUG�c[Z�~��G]-K��Lr��W;Y3>IѷQբ�ϦDs�`�v����.��wC6�Z�p�3:_�6�����)��3�����p�V�O��OH
"��R0�h8>x�eO@7����Z��p��f�B���k�>�il�]ZI~�b�NB���u ͠G���p�uw+������;�����C�G'�bf�'�(�ʟ�/���{6�Y�͊���I�A�qWV�}S�����ւ�QX����h�S¨�̳%s5 i�� �¹�0�~zV0"�˹#��ᖚD����v������}�oz6��q'����I�8&��b��S�9C>@���0�U�����ߋ&���D�� ����P2�!�fzY��u��/	k}�Wz`=P준�|X��H�%�����
�|���z��PI5���7+�}�v��!���~Eɟ囱J������bT*3�݆�&H���U��� �˾��f�9���!�!�q��r����:�rS:�N�27�w�8��i 7���Đ�I�I"	!�f�<�H�;EI��7#�i�ן��GxPEG F;1�_�qx��ߐ?��ܻ�z�Μ�
����V7P̣�.~�$��V�TU�0���_H���������8�r�z=�tm��=Q�B�!�1We�X%���ƵF�A�9{�d��T>��Z�'�-�a��,1����`���MG؞�fY�T�N�����ڒ3��?
��pN�ק��<��F�v<@v���s�8/\"T��WU�Ǆ�i���܄G��<:@�C潃s9��2l�I��/���w�3x����r�[��p��xV��������}���h��W�� r�Ӕq!�8��[nn�YUu�C�
!�ᮎ����@�@�L(�g����WO>�ggPb�����6�����4Δm������m�����v���?��]���o�����Ӻ���i�TA�i�l�a�~n{�,I�������m��ĝ��b�H��4�Z&L�	��9�eg{y=N��y�o������)���mRA�\�]����ۨTb&����|�Cg/��?݇OB�<�=���rQ�����٤��s�ij*(a7�}�,�}+�Ʃ�l���8�g��%�1j��}����8M9�W��F�>��iF�>� 4��M|���+PE��r�x�Qs����*mv6x}��6�n�'�'j�ق�Q�}p��|%��4�_osT��wk��K�4��͙����^��
��PE���H��X CCa��|x��aj'젼�̏y��xk 1�e�T2�A	�P�ח��3UԜY&S����۩��Pa����{ ���I�}-�C���0a� �Œ��&� d���-��hMIh�e��D���n��=���/y�1�O�|�0�D�'ի���Ē}�%p��*���@���Ȃ�җqL/��h���]�֬�E#D`�Vd,�&rV?����13�z���-ŉ݀�5zr_t�%e�+o�I*ن1to,��_3��3����4ɩ�M���'X�o��~�n�?WV�;E9�v�@0�~�P�݇�B�a3�;��M����ܜ��OZ޽���<K	٦i	�L���ۺ�Ʈ�V��a_̧�XS��t.�!�y<c��s@�Ó\Cؘ������y����ֲ-�y]<)��?H�Z���B��.^t�}(tN�@f1���Z�3-�rZ�֛o�*X�3я�����$�[�\)K̠N8���CSq��̜���VK<P���D����1�L4�'2Ǵ��G���h4�G��.��#�s`�� �g�5J�cQ'6815��x3Jp+P�g����m/mT�A���&�ʰ�h�K���8���[\�� R�g<��2���(�i�������&�ٴ��ݘ�q: ��|�,�u��u�f�
��@�կ3"�%�;���K��|�G�?Tfif���z��L;8U���E*M]�/e���?�'E���(&I�5d��<uv"�j���=<���(*1�mT�e1���/^m{9��(�rN0��.ZrCuuq;�4��$��W�㷉��8�����H�*T[4�"��?��ok�ڽ��P���N��%�O�|����k�8�z67����%uST([BO����������ф��}S2i����NDh1�M�t=I�z�	�<�4�����O�ĵY���.7XHo'#� ��+wp̻��j2����0���8�j�����<
$ ��{���Z .>s]��v� �WQ�ے��긏$�L]E�0d�>�"|� �i����_h�Oiܳ@'E]��3�Â5*�M��[�����^�*>`[@0�/��ESJs��@���%�H�^�����*��GN"��֩�B���&��1t5}T����z��Ѩz�e���5��k�J]�����Tc1���1vG� L�ؼ���b�X�yǿ��o���@~����N�'���Z*��%���I�)K���w���B�!�9ᬩ�cik��4Oҕ��ޅ&��}�����`D�wP�	�{��3�K�bK@cٶ��
���Ǉ\��|,�C��܋=��U<'��.q�����IW��W�q�w99F��We8Ԗ>�Ic�0�R����`c�ኦ�)���/:�O�LI�ۛ��Haz���ķ:���؛��_���f�������G,W�CI��l[d���Z��6�n������7n�ֺ��S8���43��K'����W���֔��^�M�@7�/<�2C�n/�1�
�*e?�JM�z.Z��Hv�AF�Xqf'VL钲�5��Je�DŚ��]m���x��V���8��)����u�L\؛R:!܄�Zfk͎��/�� 9;Ι��7D �mB�q��4�mO�Lk�1L���f��yn��3���T��H#�Rh��j0�e�t8	�ֳh'P`:ř=BT�X���'e�O�4�OЃ!���슮!���������2�O졕RvL��׆	bk)�#1����z{	��ÒsG�J�dm�|Qٯ�N^�jǢD�����#Ew�Q�+Y�kwN��	���gJW�R,#��L!���tՅ� }%1�>���V�)u��+�J���P����]e��m�[�R�p�����}!'9 �%�.c�b�U��'�����2�<������ci�o ��E� �V_���@���Ս����J��C+}r�Opz3e-����W����0颵����)�0H�A���/�U\z��r���E��⛰a�9\e0Рr T�P�d;
D�~�߳lWG��M^�@S��]ԅkE����N�2kg�=(�zt�n��%s@`��ه�b�޺���V0X�g=�ȔL%�,^���vN��<=
��Ȇᭀ��qaF�qЙ[ �������m�踶&�ݪGE^F"�B�gl�!���M�s"?��@y�
��[����ȅ�h}](���F�W���޺��-��6I����e�9̫.��c���L�B����uh���o�D��5�_�a:���ţy#�W�e�KH	>��ū4���x1����Iq���W%yD�˛��O�O����9C���U(F����������U��6�5�D�4�I����8V1�~u�Sk�+�^�c���u5��r)H�����m����j�z
���%u�"�G[��ߊ�>���`�ӊ��9�ϐ��o9H�Q%3k.R&�s��IA^o����zN���N[�L�K �@}��"+�\���F
����}����փ�i���ɽ`I�T��u��9[�>=�����!�Um�X�ϘY���;������,�@f���US�nХ���ރ���Kj���9�[gu$�]}K� C�}��z�&pkL5%��F���r����dY§�@2����o�t��xMh|��5����3�O,P�3��E�Jϸj��v��E,�}�+��1�r/�	�ͭ"[���@���;��ةq�3w&��oM�&4�ݟ��}���dH��ѭGӐ�H��-���M����/|/VK$G��#l;�.9ڔ��I3BÌ9,��_��ٳiN��qPa��� ��D�pzR��˜io��uk���<�x���:��	�i=�)l��.^�֟�7#���|{@O�`��3X-8�,_�d�B��@�$̎���'�0,S���C�Ky�!��}Y��ģZ�Pg/�b#0 Jd2j�����1�#�] ����+>HU��mn�d�Z��h��|����<�����A��-�mN̯Nd%�����PS��H���e�;��۫	��9��K�#�ӽ��I�dW���S1�Iu���&�t��γhI�C;�f�jV.zeEC1?�3w�C�>+`���v��*xk����(1mX������&��\�2��L2�xp�1��=��j�|�P�>�4.�GB�s�
��0ѡ��;���"�2C�ON�l9d����D n����,F�!{��ó����P"�J.�H:���4Lq�]5�~<$�eԡ  �ضEH�=�&��q.���0bc�a͘�@�����2tq&@�G�H�Ё1+�/�J���%�H�����e.�\�!06���3�-:�5�ם��G��0�^} �����(:���!�����)���7�0D�\�����斿������䡵����>4�C!�%�֛��Vl$>w�i�,�,�7�y�n�g$�:;���j�<�*���[����pNN�.��b.�O�OK�^)pQU۫�I>����0vO�BႯi�fCi�6OR��r���wb�P�dc?�2M\	#��r�7m�zj�`L�,��)�p��R��={䭿���,h]��{�jU�	��;ܯ�5\�a��t��\����E/�V9�Y'���[{���<�[��!;���EYp���}�I��K�i��й@�y�EՇ�R�2|�9��'Òl��pFR�d�����s��+o�g�󝯆�-�o��;Q:ۈ̒�5t]Lc䔸�D�ߍ)�5�mǈ�o8GE�y˵��9�;B �..�½�[��磝�27k���}���'����C�|%B�7�Ѽ�d�����'_�v�E������:I�eƲx�r������_��v��y��|
��B��F/�}�_���#d�a�^�a�ɘ�Ti��c�����#�Ъ����k�?;�bǍ=�9�	N%�+� �@�$���e�{S#�q�����|��?o�Vh J�oa�˟< a �=�ܠ/h��m1�l�Fu�0Gy�{��6�˲6l��H�^�"���hv1"ġS� _��D�8f?������_q&l�jC<L���[�3b
g˖ ı?�\D���h�O��\��<��
f�e��v��}$���3n�%��Ap�}UB���"q�`4TJw@)��]�8��UAA���j��T�(�4�(�\Ww�K�x���MeH�	����O\��뜇��D��'0��n�?!ݿw�Xxa��<S~���њ���bLKx�	?P�eZ8��[��m�ܳli[�mN��	~�X����m�}�pX����:�p)��K^(�� ���m��8p�V�h@q�#�Wm�K[�
� uLf�t����t2�Y�a��2�ۥE�X��J��y��Xh�`�04��3q��|�`M;��(�u�1뇟�h#䚱Ny���c"\Sw�	�5	���I �h�^h�'
�yrFh��>e�be��M�i	0� ��K� &��~H.�������3i���Sf�l�r^��z�;;��eNrO�@��y`������z��X�]���t����D�o�
r����N=�mZ��c�6L�Q�_���1A��\O�1�^�x�#٭	Um�
H����_�>����;Lh����:ǲh4<�tgs�&.ntz�4���˕T0!��?B�r�G��
���+)RQ�p{��?������@��4D�i�p���L�*E����n�v��@��!,+~�g[�-��������씩��xG9��\�L�C&Qa��N
"9J͎
;��R,sz�O�u�*E[ᦢ)iD���: �/�ۛ�J-#�T� ��s�3�˞L6��_;�����G9�R���3���o�<-��9Yg��-5O�i�`�kZd x�ُ���ȡ*�b��l��A��ńBm�z�8��M\k�J�+1#���4�u(u�1d��)]����l�5���6}���j�Y����Bf�}�êT3�/~�֌����x�A���''�n8IkF�f�x�ȴ@M`tM�Y�/׻����9�N��Nc� ����,^��g	�!vJl�5�%�]Z;�#���[�D�,H-�>���«�A�j����IP����*��-@�M�ja��Jo/cM��Q���e��2[���)cF|t���w4K����Q���o0K+UH~���&�sym�a�4��2V�#/�?5�sk���)Nbש=��P�Tx��#�7��&���RE �f~@��.M6���:`l|�yvuI*�CK"eD���XP���ޝ�j��u˹P[g�W[���?�W��-1�AJ��SO�?��/q޿�Fe�X��Ds8������O�>��f��t\�ǋ�hzs�_�١���l�=o��๛1�e�����?g��t�y�	�Y�6\v���YH�喖Xh��@�U���H��{6��u��۽��迨�F�v���7�i��ٌc��~��(d|Ҥ��3�'6
���D^���S���DҴ�|J��g]Fx�8��(��(�Pt[`p�*�!�IB�9�K��1;S�gA�=-F���ӛG$L���F�n���m�i{��:($a�A��C��*���RLcwb�DЉ`MFB�}v"�͜s7l:J����ɫ�7ZLo��v�A��An�5cb�*�lȉ��`D֛��w�K�&���Av�S�\J�VQ�Y��F�\��"%���nH5(���?A��݁>n����c��m�-��l�p�Zc��?����'D�~�WG'�t�/�b!A��YY�E`&��3 \�rl-&@8�мJ��s��yefc��D���/|�SY��7��6��V����n��s�b�('�S���v�j~D�IS�;"N��R�w�Q'���|����`�R�my���R��a!׹0YG.�yz<�"b&���Xz`L�c���,���ZU�gZ������i�3c�
��3��e�'�t<dw�� )c*CX�프�ozɫ��!@M����p+���x�����j΄'�V�
;nu�§yBWBJ�\��]� �TD��䚹�k�x��&*�C����OF��ᴞ��Lc��a���<���ܐ;��.�E�����"*x�99��ٝ����c�����Y�|��'�I+�	�HN�87�B�3L�`�ۉS��,(�ݿ���FU&�pׯH���5m���P�4�V%6��H%\B��w>���H)�L$� ��@���/�;mp��B��0�埿d��� ym��r���@�~/�b8�ٕ�rV��/r��kE���?���V\�{�C��s0&�}��N_�p���F�cP�F�����@䭉��L� �S;������1\�f�C��Q&h��18����4�8����7�t$a$f����Y���)X�Mq'(���#����U�C�m�dy�1x� J�=��������4ߩ��JXO��D譸D��jH�c!)oz.�8ǯ���`�T��n����OZ�@�gMUG��ə�t�|��k;-ʝ�_���S���n�ρ�lx́%k�a�I���'��$䠖�/�u��>�J�s՟�3�u	��-���r6ј���L�Z�_sw���FN����Í)��ؼy$ 
���AL��v����OSϏ*k��] ��,��^��ԣ�����B!H�=H���j��C��x!�݊.S�hF�h%�}�!2�1r���$>-�n���2i���H��Tf�Ǔ���)�zb����.w�"�:�r�"V�|�Q�y��g\��?�`t!�� ����B�¢h߰v>��x[���UX`9ٺ������3�����?w�>Iq�3��Fd�{Z��#��������|NY 0�]��N+GGå��#���c`ֳ?}�94�y0x\�������d�f
R�Ȋ!�1�隔���H���/���	.�E�G�E6�e�=�y����Q,D NM�?i�M!߭C*IO⟅Ļ��C�tX�6�b]���e���]Me����7R�Paq�n�D�H�S��Do�U#������/��vg(E�_�>��3>� ޶*Q6f�ʂ�YJ�9λ���pǢj$����H��{��P�=[�q#s�܇iW.�IW��eB�\tg��W�1��A�aP48�3ٱ��vQ%o�wL�����+/q��y��kAP��o��$p���|�~*�8��5+H�-H��Bn��*���"�jm���v��y#��~��!,���?��@��>\o_���I#F'k�젂�Pj봍E�w�$z�$~i�rR����gfA^�$��Q��h̐'���?���I+ֶ���=��O)��eG�M��:�NX�b`5�bXk�8u��ľ�b��c��S�������Sɑ��xl�����Qro�Eg9}��6i_/HR�9�b=�Q��`yf(p�sϿ� :)e���:4�����ɝJ����ٟ���<�zJ�pyf!�{D�mm^
8t�Ld�P]*�(1@t�ǵ���ʏ��lyZ�$;�dm&3�=bEuΫ�1�����Q��F�-����cz0X�p贼SS��J�ime�����`�V�}�m�Wk�Ou����yPU1-�M;&0YsJ�oP��_K ���̟o])��6lj���<R2���Ր�	<Y����������q�ݓ�|x�Q�_�^�?EI7��������檔�m�\��Л�M�*ds"4��y�\�ɰ�W��wk�'w���Sj�S�W�A`�Ԕ$!����Єb�D���q`h��!J��W>��En���k�P_z-#����U�?K��_m�=T�D ���d����N�,@��x�YI/Ϗet1�ƣ
j_��ς4����=|����saW'5�6�9��أ��#~CbKdFU�.�D��̆R!��+�J��	�E:�zP�Ȗa�Q��xJ��P�<}���l��i�u�RwRۜ�-8&�"o�=Ͽ&>`h^^�`ʫ�U�����?OS}$�q$����~��`q��}���D�]v@R�ì9/%���ۅ7�~A����͒��g��@)�4�5��^��ҿe��kSu/�Eg���g�(�WJz/��t ֵ�Z��H����&V�$��`���;���>������u�6��{�A윷A/��SI��ߎ��/���pC�d(%�`IĄ�X�?p���P;�����o���B�$�����9��ӓ ��	�q��"O��m�����E���#���&E!WFs�ծ��Ԡu7���l�oN
'	�:�0�f^�=��������o�Y�E(�4RC8I(�J���Į�G�}3į&�\� �b����a�J2�ɋ��9 ��_�ɩ�C+y�)������)�~�������W� �)��M�4���"��diX��zHG�|Q:8��8E���cms�ʕd�"l:�l�@U�<��f��_�W8�h�3R���}wD�a.��d��\������"*� �93��n��q����;3���/�=Li�*����Gk�&��9�q�G��/�l���c������I<��1A�7(�&�!��#�a;5)s�Q�L����!t}��9�M��:᥇���Dm$��:��k�*�09�!����.���y�n�qD���R��`�fUR�=�4����ݐ&���iLm�j�	4�G��;��ڂ,��D_���}C��r���`ԙ�|��rf	T+,��k�<�9P�i�H/k�ư�Ho���':�m���ɨO)�^ Eftv�p��ۡ��F����srN�+���j��yV<�&���K�7��B�>ڂ�����U�@���K7���Y��q3��@~Q�Kvv��?����uP���򥗝,���ek�{��P�^�׳�,;|(�:�q�'�e[����O- <z����ʏ҄I-��g� 6�� <��ӑ�d����/q�E���c߰�ea���ԳvB�+_�	odsd�'L^��\����gV��`%Le�Y��n�{ѻ �Yo�wj���,�f.FФ����O���ё�@ǌ�k͔�p�#8��\>�[RLH�����7P�=�x���TΏ�B5�q����Ջ|��Q�z[fV�WGŤ(I~�6�)��-���x��<p�WTK����<�@������/�!���.]U'���m��ka\ΰ{E���[v#}�ccZ8f�FtFh�w.��1�	�-���=Z��B�tv���D��'�!j��>#��o�k�]�����K���	h�9m����p&�b-�	�H*ͥ�������8GrV>c���)����\���t�r:i�j�{3�A"�N*�S��m^�#I�a���4���|�M��pg ��k>#�����"�)����g_�&�K�W�5�f�W��3�r@Z�W��z�wG�:�-���"4�a�1�ӝC�E�I�BPV�gj�0Me�.�t����9����rб��#�[����t0Xw��T���pO�Gr$e%��S�+�S}ɪ�j��ѯ>"�8�9����&څ�zl���u6F		�����ɏ�~�W?�Sz�_�UE^UH�;�*E˕(��'Ҟ�]a����b���ı�zrƻ�NA�qu"��OF��\O~�;K�@x����`}������=��E����凑�(��C>��x,���C��M������#����w'T��"/��F7��QȸKߢi�*�l�I�J��O�QEz�ș3�rai��fGp��Y���.����/G�_�������f��.��4K��i]B��鰆�:.�J6[5���ӿ���PF�Z[��	�����>~���m�c3|\�Ȏ���=;��.I�r4܌��֠#DE	�"�[�/W=�}P��eSJv��4:8Uh��d�|��j?�:m��%� ����}��8)�>�B��i�0�D���-.Igv
�fuU��ȭ���Â?��u�R`a�t��1&���;�FQ+��T=�I��^O�� bW�M�<n��s&����f*I����P����\�C���"��E��a���#v�<����{H?"�_�Hz[�\m�}|7���F����]6���Ċ>I�]���N1|��@�Og�TQ��!�_�OBVu�	�J2f�S�(r���~rJ��+ �inO�0��!��ɯ��=7�󉰲~���%�<�i��
�V��Y/���
q�|0�m�O��n]e�6H�܁op 
�2����e�n�����ֈLt3���h��bH�Z���͈ %�z*>��Dn7��w��Hi�`��;(�blYz{·xr�v��"-�.��~�7q�e���&���S#�|�g�G4�4ko���'mX���r	�uJA| ǁ3���S�fTa�lpus�\M���y���M��<�":� �?������-�h��ϙ�36�� �ӈK�w��������`G�"������.1r�o��mz�ݼJ�%8��u't���.�u�Ф��k���xy.%�o=���i�q�0��d~h��3s�o�R)9(%��P�;��
P9lQ�f��sP|�@۬� ڈ����G#."�̥��4�z;cuR��fa����p�,|e1��|�k�9%���Ҫ��|�EM�Ngץ]�WX�G{�j�&��c��H�~��7+@��zy���u���ޔ*��S$t$Y	Պj6�+�x��`<����'������x!˓o��x�VC,��U�74"�aeRw"џH%ڀ��|;40���\�O�"�e��F���TUÏK��pc�%�2��Q�Y_ߠ�N�f	�*��4���Ms8��S�Q_�U�γ=���+S���=@�U��F��n�u�/P�;č��؃��=��j�V���7k�t���vx1(F5J7W�V�{�9�X_f6^���2�j���w����ԓx�-�M�1�	�ć�(���;����=�aYC\K�%�b���XԠ��ԔY�� Ǚ�G��q�z���<�����WK�Ƴ��'�r���sy`�v��vio���;���a?�Y	��g^���>�]@���p�-��9t�#��&�p��d#z$GX$��ev~��C/�ap�c��	^����7�*��J���/4Zф^зfAGEiv?�X]��<�
�"�S�Os��V��o1>b =�N㖼��YQ;`zY7(�N�.n��&���2�%�uE�%"���m��b$����!���� i�jj��u�{� Q<�u*j@*���`��ֽ%:Y_���K�RD�~:� �g�b���U���/ ϋ;����E�6�>�@���%w,�fG��Њ��fY�H!�+�W�>�	B{w��o>0_G��$�8U��u|w�*�I��������lV-�5p5 �O`����I�/�3ߔrV5�Nj��֏�5�
��K�ŏ����<��p;�����u�@��H��1����-���.�C�w�?0?=��x�p#�ղ���)
$K�&dsO��u50;������ױy�����(��UċӚ�ʡ_� �;�E���W'��s�~�:��$e�J3.��I����-aŔnU�����_��?�(����4~���|�o�Y㨓Bw�W���OT����J'|�^f�ģo�R+#�0���=Is��|�륄����@y���Y�	�3��Q"��M��h��1�)s��W��H������������SF�z��i�=�����^G�9�f���屣��N��,�q��O�A�h�u�+�H$xͤ���{\$S���C�	��+�*���S]�("�m�0�	��f����v;ޑ�/+@���PK�ۋ�T�K����n�^lģ&f��}χ1$V��`/��S�J���R������b�ei�Ӓ�6e�_̛�NC?��//�Y���RNEF��'Q&���*�ߖ��s% PR��.¾�ܚ!�!	:~]E�r�?Ov�b���s��
���76�
��J�*�ؾ�(�Sp�����>��b(�v�ą���CA䯳�����$�c����p�i�si|v㑓!<���N�ӧv.�?�B��b_��P_�T,�8������$>�?�iD`�$��-�a�9��Hj�flA���p�
�ܛ7t (bG���[������E$���q��,�~<�8"�P#�p�Nb�J㠣��V�&.����}��!cF�v�÷�������:��d]�_b`���12��s��>�Z*������� �^߬������y���2����.������)�df���v�x��Ca����)�s�VXϼL��9O�n��<U,FB�/����l�ǆ��c����>q{B�n�J��.�yjs��[��}��g(���H��� ˠ�]���6�F������x�F�+7V?�����ÝD�	=T=�><�7SP��%�M|��R2�ڴ&�(���FQ�W+9E%/Fs��%
�[�.Kl��͝T�ӹ��!L���Ƚ��=>�#�䬢e�Ẏ"�AD��ۇ������ۨr���L=JWR���0/�ݯ��n�?���I�j����mA
�iL��p?��Yò @��m�-IȾo�l̳Qг�3#كn�q]����<a��N�a���Ruf�X��_=�Y��4�[��2l)}M�+فÛaKZ-"hpc�����M/�y���MAAy�r�����z��(���6�:TfB����:DC�����60��9��B��-��A�~GAe�û��j�%��(���<3�I����y��h^ir���OP,������w:�Q,�Y8��o��~wK��֑�	�&w�\���,�{�{��1/����>���W#�d����Y���>�T���0�:�^�$�LJ'����p�K��.<-�6 ��H��wL!����m�3Ŋ �ڥT�RA��^i�2�ȥV���#/"8�{�҇��������[����~����-	a������.m�=���J�\�u�˪{l>4���g����F��;��#C�t�w#m�ɘ/�c���1����������R�kjs�'�Gb��VA��:��{�;�l��31Ρ��'k)��Ŵ�LX���>�V
�g�Z�
��G`�70
��^�u�1��+� ��ׂV{��\|���8�B-Q���&x�ڦ,r-c�@�		!$k;�&��<��Q嫡�g�5z�1�O�K���A�Eu�_p*I����ԋ�����IM�\A�U,^{V�4T�]?yb�@9,W������3�2ke��J_��Be�!�:,ݘ�4��#���I 3�^�e�9�.��.ͻsN1F!4C�6�n� ��4X+�սB���[̾���}z
��W������}���m�$ӗ�7��^)�N��4�Y%Yrh���̵�s?�M9r+�C�0�q�zo�V�%,b�|���җ����/n�	f�f�!H^�j���W�:��<:Mo����M=>��*�'c��'�Oz� 5�R�R[{(��N�sĢ-����eUҐi��Y�i�!�����"�uc\��!���?+��M��.d�40"�W-H�$7C!�/,�YR��ܠ#EL� ":��)�izz���e�h�0}y��<����_�bE���Y�nF����������i��FW�߆y�&odz�thW5)*|X��m��4�sU���5�����X�O��^�Ur&~n.Zే�&�{8+�Z�?�(�	x�.������h�-��Z5�d8���ܟ�N���c���B����9���e�s�L�γ��w4���Y]%��,��6��߁Du0��_R�b�t�E\�<U�M�/o�	M��M���#Se����R�eE��R?������k/XUv\�P�N�3iNwҬ����g��.���r��,��C�½e���v�z7��59����-�
�B���+`�T��\oD��h7?tG�lN-�y8�5�/���<n8L#C���![Gpn|�YX�{�|a�*�s�{�� ~u;Z �YP�'|S�9V�4Za����YBl�(���Q�A\j�M`BG`�~�B���l�Nbـ�J�{bZ[�{�[��:C3E�W8�:���y�&��
.�E�J����c�l��-����	K76�tl2�GX�����Β��:��d���#嫅)h��R�4�-4 H탓�[l6�!�v'�OX~�.rE�sZG{=�	Aɝ��א}��7�9ά���Y�_�䪋>�8\�]/��
�v:�ZV�*�	V�D�Ǐ�Z�Y����}��l��̰R�]o����{�H�33�-B�Z�E��2�5}*�r��i$ wLj��>4|�@�H{7���sCј�ܖ¥�x���EP���lDpq�<�I����2<`��)��ݰ��(du-�l�D-c~ăG�̒nw�YtK��򒓮����P<��/�� L#t)��ȓN�g4+]��"�����ࣜ�3j��ti�RJ�.$.R-B� uĮ!�g�w�?��f�=����G�x���g)�1p�\�<�2�6_��ZVu��*�N8��v�%m��b#,�2trn�F{��]�.e�"�Tj4�>�@���D	}"�IY�@^�i	�%R+��..q욱7�Y"L��)˚�p8�o$��+�_i|Q(mG�T���q}9;]Q�8"�j�}��n��&mk]Ӆ|�M}bS�I��º����F�r�a�@a�
u�r�1��9'�+ƌ(W��ok��s)�%���B�C~����)�ɚ���qߏ� �rl��c~��n�C�t�0�������]�)	�k�2��f��$�x��ȦsD~�+�O�5�� _��T�㮉�?�����?�.(�E���=0�s���5�"�X�T������ة�c��E����X8�ܤ:�N���-PXXN��d��ܚ�����yh���<��Pm���EY/w��r��� &yg�e^e���;�ͭ�Ă��hG��p,L�<.��#�c�*	�T���;污7��Gݭ� ����Si�Ӗ��9���S��VĻ8~h�~;��t����"�?�7��n5��+������n%��Xe�x"��o=N�K��K��L9�М{��
-���E�h�-��+���Q���4��������
)���Z�&�s�T�q7;v�i��/���}ÜE��ص�m����o���{��(�0����_^����W�b_~�D��(�:	 \H��C����b�����_Ə��B���mm���@$h��LtlY�ip�)[nVa��#�HT�D��T��ȉ]��c���C��e�Oy���بWM!4���/}����Tr[�\���(�/&��S�#�.��k�����;M�%��&؝�FV�H ,�7�,�0"FKl`ntR��.Ch*�m���6��Ml=�@ǎ���[�t*����o<H�[,�%_yM��.�m���� �L�Y��s�xfG`�K�V�U�FB�.�\�^8֮��>�UZA��<��rX��|q�B�>�m�w'���*e3��?���D�����!=��ê��Q[�q��ò����`��F<Mrl�u<�.8�2Y���ĝւM��=���o�{s��v����-�<��vBws*��g3���A�óJ0��s8�6��+�&���Ġ����V,�vD�
�������]�� 3�i1C�����뜠�⤦��qN}�NqN�!�X���o�Y����P,�0��_$*��}]��C��'1θ������H���ʞ'���'�H�a�U��ֺ��*��Z�+?����>K�,&z�H1�Z�Ic���^��,��w�w�wl�!2Z41bd��3�6�zj9��?p�D�5�if������$2�$�A���oԊ�L�^�=-X4��©�W��`:k���z妚gJؘ=�U9W����B|/��Kh��I�Sa�`�tLR�dk]�hy�}N���$��[)q*�bP�))q�ZZ�0�����镶4���v�-`1��o��N�TF���}_pf������e�&�k��"b-4�P��8D\���8�c�r&�%��18�[��n'3@�m NΞ��6�Y"<�W�Hs��yk��O곥9f�`挺[̊�bZ��I��0���h������d����T���4�0ԕ�6����y��*T�a^d�R�����I������+RάM}Y'����F*�g��tG��4�pM��N�����"63�Roq4��U��SA�L�b懋��v�cETQ�Z4-̩�7�~D��1[�����¤�u�c#�JGo�-�����ȳ���l���7�|�E�<�Ι,w>S w��Z�;�����k����(�nO �wTY9�9O�U���!T�.s��X�#����Ղ���k�
/׍x�KQ$5:1G$�r㾡k�EQM�^�f�����I�Zp�IJ�y.#1g�</����v�a���t
�@G��m~��鴪�����.+��r�Kf��s\FBu�'͑�4ƺ�8�m��A	O֧�)5��6��7���JN�0b.�R���_�i��-,��(:3k>�"�a���b���Y�G���9P��	��E�
�r�xK<~����F�j3/���v���g�R���[��S�����r���������P�:���!�<	�\��6��Zl�ݳ�(�v��4л���\ �������`��o�����o|��1���ZJ���S�".㿽��YqJ���(P?�ޠ4�+c�D�fH@�D�d�=�7:YF-�̛ϟ��m���1����<��B��L�V��G��sc��!#tO�X/f�[������-���~�� 橉,���7Lz�4�QR�<r%�k���K���^��0�n����w,�Crn;kХ��+�㡳$Y���rv�G�S8��i�F:\U:��lmlڎi3�"8�c�KqL��Yݑ&?v[k�����E���.Jq��jN��i�]T�U>���[��ƾ�-Wu�^=g�Ҙ(��I�W`� ܽ��FH��!��_�m��;���U*B��u����y��,E�fw�(��õ�2{>��@�a��J�!���x��:$�2!E
L�J��n�}Xi�����7H�T ����w��y���H�������o��],0|Z����#}�KML�r8����x~�L}�:ߧ�w��[:�`�m��Q��˺f�U��?).@!u�%8+6�5���A���qo��_i>['	X�4��|��a��|a<��3��v����,&�7*�X�|��ẑ�FL[�k8Ev�����t�ٞ�d��E~��
e����j�@��X'�d_׺^V=�a���. :WL?9t�bs���~�
G�{�ne���0�/6wA)4��b���T��Ǩf��d*�����-��鹃��()ǽu�2!o������o�}2�,]L�po��Eik�sC2r'$&�֦�}+Gvt�H��c�xt�?b�ȶ���t���J��C��زSQ)��j��(DM}�=��MA�����̀	(қ���:H�h&��@��c�B��R���ܗ�,ಈ��k�Z�bOS�v����`�.�a�v2���PЅ`z��J�oMCw����ux{�lW�5qH.T@C 0B�# ~]����r:��,-�>fg�ig(����T�Ь��B�Dhr�+���6����YD%��U%��F�<�W�����_^�A0�H��G[t�<�Bz<�w��gg������L�r��1՘:S{��UK�,��+Z/۱+���:�r.d~dPaW�Q@����)�����#�5�g��b�O܁���#2"���l2sj\O.9mfL�R�MAo�^-!��q���"^�^L�d�X��Y��C~��#�W�&�k�bE�uI|i���U����rU0�����ϼ���[j	��ӗ��V9�9N��Hn�s�{�����x(��i\���s�u��@)�9l��E{�%+.#b*[/�Q��B+\	1��1������z���_2Qhu08�@����4��oi��,���̽(&D�2�9�������q9�� "I��R�(p��j�=��H���H�I�T�����K�fH9���P 2�pX�Cq�!���e�잦�$3'�<蟐dk�忐��'�£l;,5��՞�L�����(X��ǹ�	w��,�"g��<s��4辘4!:h4f% q�n��~�9;����fKF����ͱ)�;=��0�YxY(歍�������Z�t��U�̄,�X�4a"��˚^��I��U.���ߎh�#�x71�R%Z���C����Y`P��{��JqX�U ���ZG����� �g�Թ��H1!?��wޢv�7w�r��Uv���'J�6�����nL���Z$0�>�?�W�/�Yf�8��LX]�KkH�u?q�)v��$JU�-�Y�RP3��>5�% ��!ھ�8�#z���q�� ��y�ᭁ�a [�Ʒ�o���x��oefۘm��R�"����O XV�J�Ӓ���U��!sIu�`��xI�
t5{چ��$���լ� fah*�;Nu$�u�"l!�>)�͖3�Y��)�3��[8��tU�8]�`���,��0~Nf8"����*��?�u?U8=Fֲ�qv�|jYinv�[��r�6�] )(?P��)¬9F��3�@�A�vek�Ʈç4���Œ�<��5�֫?���@�f�x!ś6<�|&:q���*o9�*���Y�p�)f��z�0
��}�[q�f�ʺ��n�ی�j�9U�n�Q��ƫ9����\f�"�ヒ����%�C�J���Ζ�,8٘^R1�1R>S4�1���D�*t{^H!B=^��y��fR�F55$$�$:r�>g��U�E����$�q!�&n��1_�$TGq��g���/g%�. �w���7�ѥ�6~m@�s�M�4���n�?<ew�C������R�JC�\��P�d�S�/��'�RN�佀�0��L���;�?�{='ٱ\�+9$~&T?�Jc{���(�,�dH�|ݦ/$�z��U���O�G��6�sV�8��nF}�>ی�����.x���g�U�8�9M��"m��q�&�x'�Dc�y|1����C2���w�����9�Bg��H�C$ʘzz��/����5���y��T��;��{�J!�=�1�Dށ����x�S�1@�����I����&��*L]�s�;�J��2I3)���s�~������t@�qm����kr��y��t�VU�{�)	Xm�Y�q����9v&8�P��>u*ڲ�bŤ�����܈m�l��Σ�{����|��@Rb@S̹��T(�3��C�S�%	F�t����/�p���̖j��lx�jBQ��og����_�`���[�5�y1:���xjp!.J '=�>�:�����s�ƃsf�Y��ٙڕf@�4i����}-�F��8P�>��,F�H����>��a{��W|�+E���?�Ҿ��6hR,������nq��Elʩ'},�]f��	��+us��(,Qt$P+c���i���5_� ��8,�	#Ҁt���F"lx[�1#�?/\q�ѕu{�e~�w^�P�g�ݍ�]�ЉJ�K"a�5w�8ɬ�qg�l\*��W�9a<.��z!(�J���(���N����Q����}i�Q�W>^�����gf��*�/�������EY��7/BH^�gR�����
�R��R�,��,f�>,�O��lm8��h�g��l���%��]18c���@�B-���~p������,�3�����g.��я����*%v�hڥx�)-m�9vk��E�Np�Ó�Bq5BW�}�Z�H�aӸY6$�����x)Z ��?�b|^e�4}m��=e�/�I��W]uie�!�!
�>k�*��"�'�޻�(R*mC�۔��g裕`.ȯ��l��|��a��ĳ�*ֵ�����Q�E�9w�N����3xY�E��$ǽg�a`��QB��6�,S�&�5�?k��������.:y���	�D�e ٓw��[��66�A&q+(�AU��F����Ś�0��ȷ�#��rPu��K6�K�'.�oF�*sjc��2���X����%%�f[�pu�J'g;���9Nw�
`N:���� J�8\���g�0�ި���L?�A���O�#�=8�/]���Y�bm�IǊ�ax�8���]�]�r�]����WP-�gӷ�\�gr���6p��/+�̳��Wbֻ("ǻ̏��v�[�ۚs��ƈ�#p�v���U79#��g*`��ew٩�ȩ���hk�\�}��)+�}yD�"Y�^�Iż�\��^3 `W��t��IW�F
�~�N/>T�0
��<U%׍Ly����HAP-���R}�Ϣ"��o��H]���x�	�o��$��Y �Lc�
r�A��k�%� �F��Փ"q�
�\��ߚ�\��Ř�3�^t�w4J�q���	�����������6�D~)���������O��kx����w���L'|�fh2�5*;��	����2��No���?�h Xc�4A�����oY���[�rB���=V/�OD#�M$f�\��֪)��<h��9���gU�RK.d��춰.|NR�[��p�5و�w�>���\�i�ۭv;�WR�.�P��_���X�V! <L�u�b��C���bLY�]ZTǩ���|X������k=X����Ш�C�G��M�|0�sV9��˳z6��864#��$����5��)�w2�����.qXx߀y�+��YT@���@l�X!oF��\A�]�����>�sF�1�9�1��9G��b�<`U��d��Y�FL�[���ӧl-ow�ML�t��<�9/_��z(MN���J�1E����T��u1�+5�;�����*����r�25z�)�ݜl��l�盃�D�.r|�ϭ���;Ϟ+	�W�fU�8�%Ͱ<I����5{�jA��H�v�"�[����%[&�DC�����:�b�\=}a88��t��R-��b2�v��7g��du#�/du�I��a���M�̨^5�P�0_�4Y���C��5�K{�ĪQj�ROHg� j�@z;�-)͞�;�U�N8�)�(��o��o�N7�M7��1�{�D/Ne����>v����`���O���s�рs�ݘ�m��m���K�:��u�1����Lz��d��^�ܶ��(�!�N_u�onk�.1A��������F�@��.@�*C���:q0i��D�:�0巓��ps2-���ʖIO桎�:��[���8�����ua�	m2�����ʮŇ��6�P�Ʊ�|ߤ�3��.�An�O�>*�U����Z)o\P�$�.��1Kjvi��9���r�qST�J�I^�GW�C�H�-����!�U��9]z�Z�z�>r�tO\o�r��e)�t,�c�o,[�AXe�9C��]n�1r��Z �H���j��w�����CB{�֣���O)�Y�_�<��m@e�'����.�_�-V^(��O&=���G�?��^U�ct��,{����/�cOw^����]{
#������@N���@a�-�i�0�q�/ >T'�h�2����)^S)��*E��'� VpG 3��a��Wr�-��Īx�4�����
�$b�|�**��xF�K8Ӗ_�^:{.O�#C������}p~p��ϰP��nF����xK���b?���4�tqx����SC���u�h�?=�����j�"�(O��K1zt��M� `܈T���ė¼i��&�U�#{ Qq8L�?x5�o{��Q&��q���N熉Ʃ`�v��&9Rt�l�A	����
K�%*�@:ce�P�7�*
bq�' (�_�ن%���<�-���E���!ޭ?�I"Wzk-'��]�Y����٥�Q?v6�������plz"��K��Q�#�Wɂ�_�y7�V�ۥ�d�}{�m�u0�ܽ�OQA���	�B��s��{,����G(:�ss[ɭ�=�I�>bR�	���y��	o�(vU�]w�QC۟��GPۥϗ.����'��t P�lN�11��q�`��RP�!�� �%��+"���-���%�?#{B�L�di�8�FW�
;����yH��Ø:����?\�)��t��Ӽ���p�YU�"���\��4��L��0v�=ѽ�1��� �z��)�j�Yz1^H$o���-�G�G(Q�B�9@�m�#��A���Ɍ��h�09��}SW�� �j�$��f��꽳��٥E�9��V�k�+}&�4���$�=l�ȷC���Cd�>�ZRL{���}���D�X�f9��BO���䴺-����{\q/�q��Y�u{;35?i�����{7I�n[�o8�)����pذ?E�{��"r�t�#�D�WJ�z��`Y��S7��Wűn �0//����M�kc
;���oI����4{�����M!@��ZX����v7D�֟� ���xVЧS�����a��ߦ�@�Τs C-�ǣ+�AĨ�r}��O���zm��ϼ1����=�'o�_���G.�>T��F��e�x7�+�OqAG�ef�^_�Z��៎�����w4<���c� k���#��h����(M�`��"f ?�!��[�#pD4	�@	}��S4������K��eg$��ņd���"��ׯ�l���b������P$b��&]��eE��h���'�{��ͳ�P��G	$ 8���˔F�0?rW��IP�+χ�56;�=����R��h��{Ͳ:?q�e=��Bv�� �W��b�t���Z1�W`�%謍K���A�?���������D�꜄�>ߛ��^W�_�Y��=X��^l�#3y��)`�͐�6Gr 氒}�Je���bň�~���z�95�������vm�j�����j���
�K�����jO^�nk���NL�?o�xk�_��-�N���	�8x�C���[��5�q*������� �ρ/��z�S���jTK��$�X�:�2hV�K����@k�LO��&&h
E�e7� �+0^˟����@�C�l?�)�N�V7zL#�s�^�o���V5�5�9֘��?u�t�l*մ�P;~��BQL�Qi��+_�~#�9�Q`�!6fi��{[�t����]�V`�ֈrQީ=�1�xm�7G��М��CI81a���ʌ��Θ�����!��"�4��Xɦ��Ij�3F����n�H-��C��=WԽ��^��ﲺ���D�M0�IN�y���:��s_85��������I�/��g���d>\Oi���
�k2�&xd�bb�byH�S\��d"�_����&UP���Z	���'d�(4��1�����9�p(|��G��o�
r��Z�� `B�l-����~�3��_��$_d�I�U��1+��NW�gE��>]�3Ϧ��,̹:���G�l\� )]�v��P,JP ��e^��ū˼Uǜt�`�-4
��7�gp�.��<(�<���/�?��Y�Ks��~�ؖ���pp�rIA4�T�f�&�T��-E�� �J+�[T�U��od�#���,�n����3���E�-� �ָ0���;`�;ɘ�^�B��X�4%�h�P�6�޵�V�
u�Ǆ�b��F���E��Y$#0 ����e��*�nt��˖�ph�WI��(W|;�J�9�K!�tŤ�聉��������8��d0��i�ա�V����!�r6�*�:����X�l&��ߓ~[�*n������3�M�~���T�ȢޢN\���iI�`&��!��"e�lp�xY��s��i^��*��w`���U�磐]B
�6�\�����+�7�Ά^��Fo���F�Z�wF>ȥ}/���7�d#�g�l��Z�����wQ���R�0w׋4��o��t%"Z�A��Vs�B'���a��������0�d� �P�^�,NDp���|<�[���N�e��I��[��	�`���f�Q'U�l�f��,hֵ�*v[�&�2��8��
����Œ��V�.ѳX#g�����5o�㫓��j���0ʩS�h��6���0��n�8}8�@ 5$WI�g����%b[�g�""�X�/����g~�ã2}��c�mQܺ��چ���{���#u����=�3�8���h�AD�U���N�}�H�'���;����%-/q ��T�܍�SG��$�3U�c�TfZ=u#��Od�g*-,rݞڕ�d8��<��U ^�R���Ia�5NQ�!ax6�u��S�:V��K��9R���X��s�������^�\2բ�N x��5�A��Ijx���h�y�B* ����Y�&�[�sO�F�v�_t����qm��������}�{|����-]���S��q ��{�F�'}�a��s�z7����<����j��	 ��J��OP���s�@
�r�1��p��}]&{,���r�W���i�c�����pJ�I�+\�����C^�"n���}FĥF�J�&�®�&/����A�������d�{�a��]���D:0'��Kw��;
@$�.����$F�띕H��^���fzt���!QY�Z@9�W�e�g`���.w8FU^w)|k�$C4�%:���ب+�� ��jTQf�;���5+L��Ü���Zf��AT?�z���""�?��<kKB�����\�M(�)BΑ^��=���ǁ���]����V&hz�Ӟ����D��~����L�:�2%�e��0��s|��'��3%W$�o�n�{���vo#�z��6���H�WQѣ��^�L��]�@���B�M�M�ݙ�ժ��Kn�8g��#��zO"-IX@+U�B���8&t?;	%Jq�_o���G���tT��z��
��gj�����gL�-��<��T)�:C\��n�N�J���%��a;�y��(Bo��(��:����Ë+la�3
�j��,�zfDHL��Rܦ6.�h�_����冾Π��<�J3/A�6��>����s���zS���'�.)zi8�u���!�����"�r��e�[k��0�/"���aM6T��7n�h����-�h�n��|DIZ{	8�(�J�);R!\J�ڐ�+�4�ucM�T⃌`�]�<��B�f2UE�z�:Y�o�^���.���E��z�0�Re�k��i�w�C�vr���%�7!�1��<����?w��<�^ޢ�3˚�������������@�Z��&GIO��v�oQ�n���!lS܌��0pc"};��t�X�%��S޻ha�"������'iA��0�(�<ʹ������,W[�^�w�+��u�1#��F���/Ę|JN�l�Y��9�3���Y�A ;Bk�+Nf�
��������2�A�r\�5G3JKX�z�t a-��Cc�����L�چ`�v]&X��rvb��ox�*��O����K̓8�#ċ�yN���$�{�5��D��4�V��2�ED_��a�s��A�Ap�s��n�s��u���0+b����޾d�����KJ�h�鄏���@�����+���_٦��֋�0����r�״��/r�%�ɤ�Eb-���V��!��=0b8�&�SH�e��ҺF����8�X|3�_L����X�
9vJ��xxǲ1��m�Q$�Q��� ��uل���8z8��=L�?`L�ɣ��~��-�k#M�`�����Z������-��?��Nr�]7߄N�6^�Z�V�X�G��y��Q���@�N�!lF�+���J��ûAP�DDpl�*娾�`�U��x�w�,ז�y���� a�����]���v��z��4ЧMgd"�;�z�d�:�~�S��HS���4�K /Ȝ���#���D���\p��m�:u�����jc`���	��m�N��K3��9�hsi��S���-���U-9!�W����FX��$Zk0�YN(���i�u'�ǜ�ց�^fޥa���}�P��zcIR�}s��+�e�H�(0�ňl��ZM�6����9Ln�"���(���;ߛtͳcCOKCR����4.�&�B�&�2& G�gɧ5�Է8K[�KΠ�D��j&�X^fޏV2���%z��c�T}�����YOJ@�NW��A��fH��ÜjP�H�ㄽ�@Ǯ���:Z�H$<�#p@n� �.N:F(�N�ҷ��4�H3�w>�際g�?X�
r�-��\5JGm������S���j�XO*\K#���������!�e���q�n��exb{�Ζ�&�jl,��F�>���Lf��3 _�F��Q�!w�����Ʌ�s/��m^?U¶,����j��k86��C��3��"x��Q�i�Կ�©��ަ�֯�c�TŶ(��X�۴,�M���E}�;��^�ul�,��0k`�.œA�uo�����X��բiy�"��(��O���E��t'��w�)]�f��V�Q��<��u
�`D��XT2��Q�A@����F�L1H�Wd>'�c/����L�1d�{�kg��G^Q��rJ�
7��Ή�@�_uO��ㅺ�_�ȇN+?;���yt�kp1����X��[�PV�'�6:���]���>wF��'lx��n�E.g��K	���/co�Y��L*��.2)�Q�X�͈%�cӂ��+\�1�K��!v�+��/���E�K]/�v���k�/pI���vv9���+�E-*�������?:V6&(oP���t�i��NN�߹ �Q����f �4ɀ��� �
�~f��rmp�0tk��(z��7EK%����b�^�Tl
�����H��י��[��Qn@���a���Ƅ�审M0�#����clW����quoe��G���p��jx��w`�>�Mr�^�?MĊ�VV2����m�r9%��؎x>�6K��3
�)q*¢~6.����K��"m1A��dȂ�VNb6e+ܚ���(+`H��H9e�1����Hy��I�Ǌ;���xG�V��QW<r��T�kh�W@�xC�����i���p�u���m>�/%��;���F�W�Y��N�vɂ�����FNx�3%m�޷w=	�Fُ�Zk����E��,���v��`;�f��^ӪcA�pdo�/�E�ȭ���)ޕ׊!�B����u���� ��؃���%�e�/�#���v�6M/ +�X -��4�3q��.�5�^��&����ַ��_*�~ʘ�]n��N���|?	�L���4�՟+��ס�ĵɶE_1ɶ	Ӭ7�����~qy��1-]y�##ye5�$mo�v�*8��J�@�6[�E���tſ�I�^̢2	�����\չ]�d4�m����0���b�]�P?��V�B����s3CA+\%K.�m�ҫ�\���P�_��z���Ld��l�w��5�mj*���8K�Æ���=�<�5��Tx;�+#d�����p"�����b�8y6G���xA+���9���j��a�(oly���I�LH��\pnI�tS�77�^ ��D�$��c��H�8�[��&�|�#�6I@�R���A��kV͘����w���x���x:���9dQ3F��ܶȼ4W���ކC�]���1���hJy��Ҵ���hAD�2����v����g�2(�V���td�OW�6��/E��3�J+��tS\�V�M�r��'���ƫ������9}�Z5T��Q9(�XL����0J�J���?x&7\�2�V�66�|�@�)AV���%�2\Y<`�m$��������^� ��r��o3��M�P� #�f�� ����~k~�*�\�i���67�of S1Ť4�qY��E�y��}��X��6�߮Cu�p���J4�"��7�ο�a{�T���O�AF"���,0X <D�)�I>d!��,HB/�s�(��.��9���ӵi2�&�����K�&���֪��_U�_@0Bط�zU�/�-cC�/_�\����4m�F�ɽZ��k�Tcr��B����.ZU'*��r�2狀�H�;���.&��ZK�?�2��sZ@�~CYg��Ӌ7��֙<��t���SQ�7�7k�=\{E�o=U#�k�}IǞRu��L��ci�9�Aa��Q�KEy��?�%�sN��չ6u.eOq�����3)Q0�
��s�sB�� ����7\�2�W]��]�S�rݺ�ͬ1�a:M��T�p�@a�(���j�g���*��������i��|�7`�0���Θ*�/�Te�C��V`C�y����G���Z��a�CV��}��X���3�;e�x�-���F;���墿y��Y�f*	֟.5-n%�r��%�k�o��$���Q��]��y����e��չ��j���mhH�\ؘ�ڸ.��p��u�D�
UA(2��cN�(Gr��9������h����g�1*�Q��k�Gs2�c�2�5�UMo_Z
b�\����UY�_=��pF�{@m��F8H�⟉����d醋Ȁ6d�GYl�޵�ֱ�&���+��qG�����˥KM'v����������d��^�ֶK����J�c=\��)��?��Q�F���8��L�aA�J���$�\y���a�>����Sl�{�T���XoѠ���j�o0g��~K�y 9 LI��d.�ƛ/ﰀ���w����9��La��j�4ģ��G��P�'+�û؉_Jc5�������C�c]�@�Z-�F��nY�=(�G��^A�SE'.�/��n��9��|#\�:��������zE*\�$4p.��Ԇ�*���w����0(�R=�=��t}��] ?���R��#�1�)gy�?�8����k��7�2�\�p觯���jU��L�fA���3��\u�[� #57�*|�랂�l��毱�G8�W����k<���L��ܐ�N��Z�S�~Q�s4͹���*�+����l�x���ˆ���Y�u��7yJ�b�����F�-�G�i���[cy��rG�k�5.1V����IN�a�&��ɱ{�ʱ�:��Kx��ZD�#gn4R��1�B��{�[#��U.�� �D��^��������c��`��3yZ>�6Ы�tF>\f��d�h#H��Ax���}�L����2����řU@����1��z"D�U�����Df6�~j)+�ۀr��C�l���0�%0D�!`�BxS��I�q�����9FR���,�f��s��e����E�7�U��e�|9kh��{Tf!:P��ɛ���l�H4&{4�Ϗ��FCTױ�<�n ����8LQ�.���Z�S��+���z>��Z�ܯl�������Q|�Vo$����d�g���
ùnzP�f�oƵK�Zb"�>����얒�(�x�;�o��v�n��|�ƫ��&E5��*�\��!�1Vg�At�Ej&�7��`�F1���d�@0����(9��}�j��%g]�1�ՔN*Ӥ�t�� ��O�H2�
���RhWF�ͣ�o�3��A�䀂��"�K�uk
��1��v�H�Z��0ys����K<�EFa�m��ՑY! o�|����@����@�D<!: ���.��U�o�O����դC�V�����KY�#�,Y;�r����
�&~����9�@'G����xh�a�EF�S�\(�[{/>(�!���׍�틧d$j����� lld�m��nso��%픆���c	�C��?�x3�����l`�@��fF���QJ)�7�H��F���S�/·Qâ���H�,s�DJ�8;S?�)&�=v)z��8����H�Ֆ-Qz����� 掰�2��Z�F�H�$�wm~�R1O,�}�9�h�'�6���1z���� �W�X���e!�\[0����������5�4�֖�	��U�P
��jĺ�3���f�H�ca�.g�q�8J�{u���&�&�v��hMk�f�hV�Ĥ��$��-4~�+9-{�Bo��h'��/1�C'�{c�/e.S>VBm�� �t%�݀��40����5��F5A������6huh�'����n2�:;g��Os(��B���"/�`��<`jUdt�U.*��Jk��n	Jo�c��	��/����	�)@(*�We�-�a�OX�iZ���D��M��%���HJn-e"E+_j��������A2�E��>�t!\SƼ>bS��x��\�5GV�Bv���^�^�96\��U�7Ra��)�t�ݚ}�,XB>�O^%h,���#R�.��;iI]�p�5H�@�����KҒ�g��-7�=��xy ]7�$PL���H_I��i�m�`���0��~ O,&:�Lz��1fr����ƯVM�T8�M���fûc[�:�y��\R�QSh͞|�	K���@m	���0���9[��?;^�3G�/ǢKbϔ�+q�,����Q�qܭ�M��E���
(*��sbh˪H�����Lʧ�{�Oj�Va���������Ѝ���m��`�~]5�l:`�<p&�KY�B��c�8��v�V�c�b��Q�7۹ �Ǐ���r�-Q����x�R�ŖRќq^Ig��U�vz?^���I����:?qh�Da��W왰i�)��Nx}5K6�G�����&ʄ��%s�[¨����绑#��A��RJ«Pˮ̝�h��:Dآ#AZ�n+	ӍE�V�9�PL�$�mekfBP��\b��Ip.q�x�Ã ��
ɀ�eDJ�j���+|��Vl�!������^��:j�[�=�x�#P-����o�KG}��|�s�&��+7�$�2�e�QvD_d���|xZe���9������"L�~X<R5�p�aBJ,�ö����{|��0uɬ���h69lҞ��@b�W�L{��A`p�AE�\FRP��N}x�����B�����ڔ�zJ��|5��3�3�o}�X���R�/��b�%p�ʼ����i�!�]�5\���h,D�,&���M:�h������n&8���4z���k�BswĬ뻖�ʘP�q�,��Ls÷�%�T4�d*�~gQ,o+V�`@���]��"�����G�0�/��<vu�QŲ���\\���BԦ�� ��Z�-��d+��mD(f��6�Ɇ<s�ב��(P�����ɫ�eA+�:��DuEC�"��"N��-i����%�#�'��)��[�8xJ�te�:�?����� L�u�i���d�����&,�P���a�M��GW����tSr� ֘s���.�o���h��љ/5�zu�r�b�]vm��Q|,@C���n�'�Es����hoꥀA�R$���ﻍ|��:^�6@�&Y��Y4.�P�k��ȿX��C������0�)4!=�o�v_L��/���8K���� $���v1�JgȪw�zr�S�n�N=������4�����
�b]��.�f�߈M��qR�/��v%��n���FU�I��g�I��IM��b����~̕�"���.)P@�OϪDzI^�����Ds�E�T���w�CΑZ�7�wz�U�Hv���a��rX�:�/�֛�t�s��b�R1z	|bFn%"���mDc���r��;�h�bm��>��x0HNo�]$MUq��YՌ ��7��r�/8�
�Z���l��uƎ��~�I~��t�}\H��J�hGᡍuh���+�� �2�0�7R�?o��� ���
֊���f25���[ %�����I%�L+<��#OT��c��䛎db��b��G⑀1a����AyĎ���D�=�ԇ��*�C�u��W��J hht������p}�G���Є�n`���p���K��O��	�`�昚-���S���ס��/���F�[U4O�%ۙwx<�NO�H^*E�/	���`�9��p�^mɘ՚)�B��N��D�w�,QA��V:�v�8P�_����4�{�xjWq���+Q�XN�D�ʠB��
��v��aO"��(�2nɨG����)���8�;#��ftKɄ���4*D=&�=]�F�B�z��CS�����p�q˕�ي���c-��n����h���Ign&'�ќa*^��$,C��Wj8!�V⻴�"�j�/����䨙��w�>!��+W$?�ɴ��i_ە;D�k�V(�iĞ�t�F:b�0Mr6��-��bI�Сt0r�ZhlB�ę�c���n�@Q�
���xMU�W��жO�m|&A��P3���������y��;z��G��rw�i뱔�ņ~����F���j�9Z�G@&x0{K�5��
��"�UN�/��㢇�ڵ���7q�������t�3���2'������#�x��&V��I�LC Qt�0n�����|o0�����E�x-�pRO1ȝ7�4<���{ˠ`E:�v��L!�iOg����>��Lz/�n
_�f5�#�ꦊ��v�'�'������j��8�	�wu��
B� ��'D����r�U|��u�\c�L=w� s4�D)V@PJ��r�p��<��5�w��h#a�]�y�²�0 [��z��lDX��)}hD��\v^���'o�Q�	x��-�|s���;�n�0����T�Et�|w���e�$Ԅ�5mF~������øev	��9���rؙ����N=���D�!x���KW�c�\��^zՌ*	3��We%"��nP*(8^>~PQJJ*~��� V��3Y�����X�I�h1^�t�p+K�p�V�g�ݢ�����{/L��]<�_�@���f�+g̣f��˸��R_�T��֭��{Tf(�f����h]�H	�	8OҺ
���γC��
��)�����D4!�
��Tz2������������|�4Oj�K���0��h�?�-�x�n|���̴���n$0��ؠ��D�E�u���1f�ueZ�a[�%:���9�
��Ǔ�v���L�_��U�l�}eq:}�wT]N؃� �a�8A�CeZc��s�O����mb��nP���z��R�:<���`����
`�����ȩ�Mzc�6�Mz�T��tE�i�ޯ��r��V�B:o�KUO�̽U���C���fٓP�2A������ �a͜��"ب�N
FM�]�F�Rh�[�?[/�ņP�w�Y�Y#��&�}���J�q� ɲ��2A�ju��T�];�a71g��hN���%���9���͠��x�b�����%��������P�<�~q�+'��ͷ]�I����`���+�r��{���eg��-����|��Wת���6���-Lm�lx6>� ��j�h�����04.�M���E!�=�d�ԥ
���	�]���]��_��5$a\�`�U	�4��������"?˽$�6�ZKo�̣�\�3�팹���]G	!���|j���Lj���Jk����,'<*dx/!�
��ί��&m�g> ܱ�>��yi�w��>G@@��OW���cW�.9����*�+}V�>S�%�1%��UR�ٲ�RX�t�Q�uD�&�ӻ�I_�{�K[r;e�ֺZ�d� ��2�g���wCI��%Ծ�Q�I�dO�]��.~r��d����;��e5�8~�rf�V�L
J���u��U%����(}�D�d˜z�u��?�WkN��+GS�Y#������M��k��X�zL�-��mP��֝�?�L%�����jd��Ĉp%���,}=���AP�,�K�g�$����	�m5��YI	V�wY��S@{<�~�+�"����?�=�)m&����q�V:�[Q�7����MQN� �d��!�Fk	b|dup���cu����_.�o:=ܝ��8:J�oM.]�a.��?b���-^��� ����Ώ�v����R�^��,H�׎���2�IF�6�o7WC��������h�qGb����}e�Ku�+�&��퉩\���vN�!"��_�l*w��;Z/gp�,���/������Q�t
�Vl������E�|�h�6�=A-��$*��F��JOw�N����>�Af�|�4ò��[�H� �v�{Bl�/V���CUO��H�^���z�I�?ӆ�v].`�M�3ĮL���m/�:���OxG ���wbPX#y�3;�g��@K�{5c'~�5�9���p����=��Z�S�CP�FϚc.]8��)��I�0���>�Z��`��t-ݮ��",�D���Չ�UȽ�^����ӯ�+%��(���+ٌ(N#ރ�8�D!��1�^6�	���^��G�� xK�D�|�nj�7�1^-XQ��uoe�(�$%��3�E�(GdQТ(Hw7:����2���؎��4��`��ѰFu?��L� ����P�bp��wi6�i�����z�E�k.�Ա��X7��ƙq�N^Ѫ������TZ/k,�Y��>RpS}��2)��i'��V�41�
�T)��-�M2S�ټ�GZ� �pb�`.*8Z�,�dۡ[:���cl)Z�L�a����H�o
��S�4T��8c�S�����UO��D�1�Gu86���|~W¯�k&�(��錞�!#u���Q��b��>�'��[^�=�丝��f�c�K��ST�m�8M�%�Ԝn��W��M� T%���-Ѻ���g_u ��0����{�ގ���Gq�y����`*��t)��U�D��L~t?�P�#�r\U��k������7EiYI�} ��҄3���cl"�r��
%,Ih�M�I�e��Q.&4y��6�Di���|?Լ��zd���U6vw܀0;j��/���$o�s3��5ǂ�i��bz�{��;fAo��>�/��,9����P�L�1��z�E��Jb��z�cЫ������.egܙ2D{���ؒ�%�С ���Nc�`����:��M�}�c�h^]�O>O��[�nd8�R�{;�hR��/�	�A��+o�ny/n�V��覤�b�Y+Es{?� ��	N�ӲR�R.���J����z�mˉ�����>�a�0�A�I���S��%�*&]�)�/t�2�{�+���b���PbD�UO
].
��Jh��T��i�Ҷ\��� ���z/Z�\:j?P#uK]�8�6�*ݴ�$��T@�@�)�}�#����ΖhO"3J�4�C��QT�!�^�@�A��H�2Vc���O�(ŉ �B��E_�Q�+�����g��q��J�4%wq���n\=(�
��2_1��8�T�.9w�W�Q�Z'2 ~@�^'��g���2�6n���1nM�ukŒ�I4Op����js<T0�k�����gĎ�&07��.��d*�B�t���lw$��j�l�z����Y��q��O�P��Qc�^'�J��Kҭ�3�#{� ���)r�gLl���F+w�n\=,�@wv�$��G ��N� ��Vd�=�g�L���*W�?ܤĔ�!.�KZp��LbC���.��wNg�-��BH-�ڄ(;Dt��ĳK�G��t�~�l ���gf.xːI8]]$�?Í�H�t����v���=���1�K��N�A����i>=?��'2�%ɦ���q0ߙ����g�g ^C%�z���1�C��� �Ң�F�b%g{�e7/�587��#'���8o���O�Ll�eº���;�7�[��T�}�ɻ��G�˧9�ݘy�\eL4�l�kX,bX�/Z��e��aZ���=��f���U�h��m�Wѧ�:g��@n��kh�I�V�ߓ؝쾒Ep�B,u*��R�)��M��lɦ�����YyH�7`O<!h�r�Js���r�j��~�����l�aH��`=%� ���7S0��H�=E��*��`"����D��Kc�m��1�c����^�"�K��y�Z�9μ�2Rw�X�[X?qm�H��5�w�bԡ�6E-+���DC�RBػj���3j��<M�c5�]$Q�y4]-�r,8oZ�D� �Dߢ"
_����x�S���4
mM�O�p�x��Xr�b5�w^���"E;�D����?Fr��w팿��re�4 �ݸ���$z�*E'\�aWOq�w[G��>��`�}`[b!Uko��`�DY�}���Ӆ�hwBH� �V/��zN!�Mע�
�.�* �J��M�����q)=��3q,�0�v���*dDT/L���PpxW':�t�gL�R�8SW�(����Ktn�Ȳ�	����������� ��pm�@�l���ƞ���_)0�Ah/ؗ[���Zx��(�.�r��,7�f2W��ɝ��+�J�m4��֍&R�y[�����Qq;��,s`E�IC���䍽@�I޳.&�hu$��
��؎��ե)h �صԧ��){eᎬW��q) @��!�y�g�0��U��"k���t�FԒ%�C����8���;��+�($͚i�rH�S5u��o0[fc��&����{BWF"���qH$�C�m)8mdE�{���ag�F	Wj�K7�ݤ+J��k'��k:��ٿ����U���u��B�����p����Pv<�s}6L��:�z��kfzk���7*�W�����M/�D����Et�k?;����m�F@~�(����7 ��F��  �_H�a�V�n���Y�@�~��A2��a{���S��^+`�ݱ�=�.����l�34�*���[�R�:�,U�#�Yo��0�=S�Y'*��d|���"-�8(֮��)�ҠhmJ<�A��
ǐ�#��$��ӬF4l�^s���i/m�6HX&�������b[�������«���5ڞ��j��0���\Y��)����+�2k�*�0�n��׵�����a��h�����k�qL���e��ߝQ2�z7�tIl-�+�����U��	[O�Y_�_��M����\p��U)���������R\�#��+t�tNӜX�����Z�!	K�"ΓAj���riuIf�]��e�yԽ|��r���$Ih��m���T���,��J�|������2�����-�0Ev���� %:����v���v�\�Q��{�Y���x�E����c"p��T���$9��F�/UWP��� 
���b�m�$��׋�h���j׫�������>�;�H}w�Ԏ�(����Cc8��z�����!�,#Ϲ��X�4 �O ����x��.ts�Α�*�ġ��j:Z�$���4H����)[�c��'�2B��>c�1:���k������%޹�PE��B@�vl�G��-]��/wOi/P/��86ڠ~����:=�"�x�v4�[���Y9��R8)���+K7�I���� ��K��~	���x���Q>���c��ח[��	=����'�7�h,Q��Y,E8���cy7~��9�ݰ�[��@jtb�Q�Wg��i�7��L[�ͧ�
"�d�2(��V�н�r�<�ԭ�%\:�,��zH�M�k��6돇��CQۂ�%T)���Lg���JP�8�h�pU��,s���$?0%5S*� â�UY���7�3�^_�M
L(=�g߹�����I{�N饵s��kRB&�RZ>�:>�A^L�/`h��~��	V�Ӽ����D��-6�#} �- E�6?QZ����A��<�`b�{n�)�F���d�a~́�BJڱȨ��?(�qnc�j�xC�Hؚ�A�  #� ���]	M�Dhn��9̌��c 8�����x9�b��Xa��pD��33�LI�h&E�A�;��x�8�"j�[�v�έ���~��'>�5A� A�#�+|E]�#$���0d%��v��5=X:�/��1�C	�=�.�D
3�������4�ܿ��6=��A�MмN�m V"c�f��j�uo�w"����*�(�́j���a1m�f�1�2�,��a,LWA"<� �:a�X'�k0�{�dl�0	������|o�k��|���j�(}�AFV���&�%_dAYV��G����)�ִ���d�2�_��j�&��Iz�y��M�4��.���BcA�cxMckk�D�W�n��
�_lSM:6�1K;j��Wܫ�nR��G�h a:����`h�ߞ>�ύ��Ġ[T޿�k	���d��	y1��7�;�M��8��s�p�HA!E��ZO�z(݄t4���ҳ�K���Y����Q��ڵ�ܭ��\�a:�ɛ��d �����Z��2��.�����:�s��ڐ��\z��)��P�2��!>���cF\����a��vt�l�ao4�$$�r�D:\a**�O��@Y:n1i�@�RM�����$ٛS\����!���<i\e5_u�r>��V��,@H@��F��'j���,��
�J�`�$2q��u�W��q����7gμd��E"��'�-�$�c�]3ց�����=c7�1�P_h�աe"j�LM鬱$<���w�h�a��i�����Yn� �(�uq[����l�V���R�[P����Ҫ�G�eJ��W��d��N�����ެ�P#v@�s�0� \RuAc���2���c)���A'�t�(�M�����8��q6|�XGj��U��fET݉����xW�(��e�L�W"����.�a�q�7Ɇ��� O�����=e��'��^���c����]�z�;�}�l��<�����<�i��N��ȫ�*�vt�y�T�tt��9�I�J~��b��H� �x��T&�UW����`�z����&����ԟ���Aؘ<�"��.:�S�qŋH�l�EA��E�h�Mxc{jh�v����(4O;���O;o��w>��/N�M�[�(Pn�"6 �
*�4Z8a0j�e��(�b��u��\�E����+O��7�&��������Ycz�p^��k�����h���1��R�DR��	��Z鸹7�%'�����h��B�\|������u����B����MEE9H�0�sRi*,����r<��]/���ѐ)��6Z���չ�n7~���W�D��j�� ~-����}E!9 4i`7c� w�@�$�gX�<�VS~�j9��Π�b����-��(��^���v��P~H��v�AN���<7�%X��1.�{�R���I_v�rV�P=^^I�Ʊѩ�JMe�!| �����ŴE���y�C�iZ�A��It�
oq�E��s����+K�:�Q�|����g�?�0��9\�s?�U��;_5\V��M�ښ���MRW�M�K�[Y���X�ɰ�j�R�5ږ���'ZK�xO�̃?/�_0-�$^�sP��6��z$�qZ���_Qz �����S��8mW?���x�+8#a�y��)?T�D�� �T@����&�T_�[ �zԯc΁H`�%9��]��-[<7W��Q�@���p�F��ߩ!��x�M+T�R:��+�c�-=�����)�=�� g�K��nwԢa�K�V��q�\1I�*����}X�q�[�ir��W>���c��
�:��,q�ͧ��bH32���'Pƺ���=�°h�$���F2ս�أ;x���W�Bb*�%��wuF�ʞ)F2���f��J��:9���tV7�H�]4�ȵ\�d�wՏ�{�I Ѯ����cuc�Ї���Ԑ+şGrt�2k�)��	G{������*l��>]懹��g̎)Ja�%yg���0B>p�4��qL���a�v'�|oM����D�#u��8�A�ē��͍T�
2G*�b��J:���)�v"��W݊f8���5�˙��Auiԍhw$y�i�s�YaSnX��<��������!t��s2�����L�a{�#��ު�#ǳ���(8�C��kxWX��-�ҼR��/�SH�*��刣�mo�v�u���dMq���9�:��өV� ����g��.�wfa'S�J���.S��i��Qd��4���Z�nuk+Kྺ��������)����V�'a�����"FL9���ʮ��
��^��S�[��E�@&����uFN�}:��+�m���k���jY�Q�Y���!Ti����!w����,h��Y�c'	���up����#*����u$!�7?�{dc�����E=g^��	����1A6�Ȑ4ȳQ�7�K��vϨnW�e�Ů��1h����}�T��C�����xd���z��a�lu�;m2][93'����Uǚ�{t�\Q��-�>u�j�{zM�
2�t�1Q7�B����j���|� �/��}d���D	���b���S�6_�aY	rsg�A0
_Ա�B���-J����]g�ŕ�9����wL�;V�A�x'Y�j3B��Umj��mg��:��/[���������N
�Ҿ6ð�Q5<:�T�۠�h���9���.��tG%%��Q�����F�������kԇ������g"���q�\Ze����>�7��Oq�VR�w^ymGIJ�$���S�ބ.�QO3��] T��B��wuZ'��8�xk@��0�����0|i������:@s��j0��������(Ø���Ga}��EM�:�{=5����ym�h�1G��]٠��d�'�y�SSlxW�lR�ȭ���M���_d�$Pl�"��{��+ё�*l/r֛w{J�,f<���$ܘ���4b֙<��^�H�W�;��R�q� ���7AK�u���3
R����>�X�q�22%�	���V��B*�7����whrm�b7��W@c@cP�q]�u�Uo�&/�n-8��t���}��|ʸ�$)���p�kE�No�[��8�.	EiӴ�.U�P��ad,��tQZ���>��}}��c�f-ݘ�ˤ���,�Wj���=3$��ʍ5���I/�Y�K��{�Ҙ���:Q�v�͂>^�?m��0}��/|��:�vy�Rrq��Br/5,���ܜ��U���Y0��c�b�fd��8��>���Z/	�E���C!q$ۊ���h�ְb�0A�ϭ�eu��#F�:p�NÃ!FM���̭� ��?=4%�r��.�h��E���b\���� ���L�f�D [�p����mM�Q�u�j���QEh�8�4
��^VG	�(��'c�VrPE�ƟB^+c�Ȍ��,�	��b�o����/�Z!�:iX�e�ڧ�ʭ2+0s��5(�M����B�A�x�A�ɢ����`�]�5�����8��1�M��"�h��v�ý�� tZ^��F���A�U��کCG��7��1��!S���uz,�wM�}�my��h�Z����5�N,�3 ?^4p����U�|�X
Á����P�/�Rr ��i=ɹ~@W}��UygNR��dM
)'�P���=w��Y�[�g�VL���+�$)��E4�U��3�Ŭ��S�.��H��V~7���r$����d�y���7Jޚ5rAO��6A4����hCO�'��/e�\���zU�7"Y2�g�����'^�<9��P�>��б����"�";�V3�e�X8nĦBN2zFK�>��#�d}#��H�*�KI#*����
P֊���L��>c���rT�'�a�K�/TT�����GY�7@n��:N`TssK�'�E���^<��/�Ae���VL��ˉ�;���Ώ7v,������QW?k�7�7�b��G!�Ϙ+��$���y,��˺���Z����c�1B�6��Et��=~\��?>���ܗ�]P��{[Z���~��v9j@�G�w��`dM�-��U�+��z�R�HO[@(B �\��?����6���V�8Y�%����`��n�y��ma�;jR]�7������Ƣ:�-I���Ν��}+���,�[�$��N肸@���>,�ӌ��/ھJ�fr��,�!d-M8���X���2J����2��e}��<6�:���@3� =��[��#r�tM闛��ܱ瞜��޿���z˷C�j�X�f�i���c���__�n_(X�'�L"�������M|�X�Pn��>j�
[&��4˾Z1�#բd�k*P{2���=޸�A��GM�\����ڵ%L)�Y�T���}�z�x��ߞ@�%����[j�&[b������?�*VAj�ڂ�[E0�z	�΂�V(+�P��17�lV\}kѺ��AQ�"{��yB\⤺B�X�X?��@�wbNTd�>���sW�#��h?1+W�0A�Ix`���`��[����e��|A܀n���;pQ�&��g��;���R����|�¯ڔY~���P�(O>S�<jS����o������q��� Q&zh)Ռ��!���lq�7�!���"N��h����}��t_Hy1W�u�b�d�ꆖ,�\s�/2��������c��=ɒ��ktE*��MK�������$6uU*��Ȥ+������ſ�o��U��Ky?zɺ��uk�3�k#����j�Y[+X��E�,�b��z�\��W�_��P�ý�#@���� ��i���{Иj+�����#u��E�X��x!ڎ��G�ƺzo*������n�F2G�n��Y�v���*1�Uo���#s]&,��q�GE��нx��:�����2�ˤ�҄��>T:s��3KǑ�����8}}3�ꖣ�A���m��^l����L��O2{1Rݐ���G�Ƕ�,[�>$W�<����{6�~G*��Ȅ�=˱ ��`���r�=�!���6�G3�#�Ci������؝}/EyƝL�*Ŵ�A�D[�5�����a������P.:�?fq1�ʦ��I��N�T�<9ٻ����T����	�E:Y>��p��W�}�����X5/sڞi��b����k�����_�BC�0�k1ު5~�[ݪ�)�d~_x2�̊D9�|<NXxMz6J��?�ox_o�%p��si��Mvq���K���6[�?�O�s�,GHn��%n�q��`)��s��yډ����0r~��J2�p�b�)�����F"�D�ef�Wp�qod��H�� XQr��Q��Cn )�7|�䅈�O�+�5�f��Ӿ�B�/�s����^?�3�F�	�N��;�8�9���Pʢ���<N�t��4[dRq0���x�<�W����!c�7`[�����U� ��P*�7���gm*t��sa�*���QS��G��y��	�#��~�*9���H\8;�|��R��1���F�+�#��ϬO�ؕ�ঈB��nape�#���M��M���R?�8O���pf7��A�6]*���"���R���%���x�N�;�lb�\�s�C�z��D�~�u�/��c�-,9X����	���/ޥ�Ĺ(��D�ATBb�3�+�Fʳ�vp����ם���u��~�ٽ|kZ�ڠ��6t����lB�H�1? �(�ov�h�+�
�Y�� �8�7��3~�a75���P��,qcj��`���w.>�/Ɋ�zh�իE!vK�t�TGM��5�w6'E����_��[�N�:����68}�3a�ub�*�N$�5��<�R٭�8T�7A���X|�h̹>詍A�bM���0�1��F�s��w�x/D���K8xm|��n�7�~[ad5jCq#�#R�zsV�Z���������Q����lT��Ҷ��.��R�\Y;�� 7�r��h�!R�ǜ�N��iF���<�L���d�<���e[� ���i;9�P��Bì\����.VA}�{$�t�m��.�f�f�b{������!�EL0�%+��'D�S[��v}MYҫW���p�|4�Ч5���C�t'?5x�݁�|*��y���b�W��0cb�V����s�a�����n��f��*,��Q	A���ߋ2C�8��,U�
�ւ���N�|8�M�*͊���WG$ɗ�po�&/�%S#]dm�Ѡuc���x�r}��c�Tt�����m���"¤��f^�M���@:��R�]ɵx巼l�H�	x��)90��r@dI� ɋ�H�	�7�j�d�tf(4�[$�`�K��P�uB������H$$��8�9~�8g�}�&Ȫ}l]���TϺ���Wh��~�YYZG��g$<dmm�����^��?0��{w\����gM5���D�/[I��q� �wS�%�������lvÌ����/�d��a�H��}�;�x;f�U$��O%kzZ=���M-���,~t�����vI��-�߿L��uEn۔�h�+��cd ��|�j�ʆ��}x���j�/�Rr�	_m�Ib�F���ѩ�b�k�ɽ3�|X+�� 
�PCa�rfTL9�F�r_�a����t90�v�ʳJ�?�4eAP���(��.�cXꬕ<Z�Y-�3��3�lmo�~ӝ��1�Z��4���ab��%��4�>��4E�L@����-P�0���	=�&4�`e�`�!�:�lUw������p�����_�H6�&�H5oj>�5��IT7��3�F�݃�Ú�SO^�܀��L铫߅�d�?�Ț���D��Rݾ϶��P�0w�uDm�c�w�хp�-��=���^ґN��~�����������0䶋�xڑ'?#�����j_'�	�&u �7k���� $0"G���k�kI�0Nmk�(���K��R%]D�z�Rb,9#�[ĕ��EFr{����J����%h7u<�B���T�����o`0��+��<�1_�{`��n�5�B�%�ri�W�
E���t,E>k=�Y{.2�@3�FF"�	���
�'!M(A�*;��>�Z���ʕ�H�����$�byp�q0#���k���qS�D�~���Z�sRfvn�^����������Ey}dz&@���!{�����B��r��3L�nZ�,3��~���q>������K7�B-|(�Nh�g�B��َ������m#s����R��U���#Å�:?���}�^{aI�n�ïoÁ�/2U~U��	�v��� �la�t�£��%)t||I��U�0c#Ŏ­�G[/8���}�]N�y�s{1��V�*%�����;.��V�ԹZڱ,l�-�B���BA�S��W����[F�o��䬃.Xn����+����V�����m��Dx\#-������_���55����q+Hi��(H!_�$��ﷷ?��g�������)����ΝF���:@�����j��dl�3u'���r��*�T7�g��"����g���;�ß�����>C��"�������/m��K(���oA�"�w�wt6ݮ�Bcw�?Ŀ-���1Rc���]$𤤵w��/��ogk�Z�l�zu
:���
}��
Ԑ�+�"���QK4���U�(���ɔ�+۱�����a8�v��	a�OH�F���-�|n7h�z 9�*���V���x-�T�K_��]��W��;Rm��_�}�9���J#t1���	z��UpyP�å�Vf*�0��.��P���c�da?72+�j����7�Y�3j�$4�.�!��$��
�R`�m��m)ī��5��a��0�M�e�o�v���8�*���&M�J�� �����f7P������[E?A�`�����I�#B�;�|��:�p�?/�x�nב��u���7��s<jj��	���,�u�2�C&Y�d�Z9�^ߎ��U���u��s"�jV+]�)�Y��
���I�a��Q.#-�8,�d�Vȭ�U�����E�B��9�L!6��j��#{�WkX!���L��Npo�N�V�M��9����^ ��h/�8 �=O�A�DL����{���J��L�؋�>�gX(mZ�z�G�:M2������x����+�N��Z�����D§�{|��@!�4i��N�?��#ֽIpR�������9+<b2�a�����F�z�8��tp(�����So�om��'~p��=�pm�e��w6����1�b��J9�Vo���<�� �G��eǡ��p�u�qK�$�u��w�j7��zu��ۢ�nA�pq���ݿ9��cH�\��zF��]Fj���.���D�;oi����d�Ѷ�s�A+׺�Ԇ���������4'-'��0�f�u;0|�(_X�:���G����S�Q��7�P���Ԫ�P@} T��rN~�H[.��{�s���39���2j�̛ȷ��z���|�m����ʾ����x)^�~��i/���Q�&W�I9 ,m����N��&��Nd���Ϧ+��m��@x]}7�P��5сC�c K0�o�i�>�bw�:�0�M�-C�d��Sy�HKi����ʠuu��Yp@H�W�3�:�[���&�7ML������>B���p�m�ˤ�P���=��8��ܒ����*!觊�MI$�|��29NTO���.Y<�����hp��]n��+� ���@u�w״CX�������*��`%ݛ���%�1�;y�������'N!#%��m'+E4 ��(r��T7��W��8�m��)���AABwp˗J��??��LYj�����w�N4�E��}\�Fs;��塂����%��$5G�'q�ӌ������ � ��1n�b�si��������
F����^��aΠ^��J��{q4� �X�]'M���*%��N��i��	�aIuh2My��7}��W_���巩F��ʌ�q�������j?TJ� ��\��?PJ!��Rs�+�Q��[B�;ZNMq@����f9�M�= K�G��b�Jժ�����1���1���x:3�K"��e�I@N�~;2�T��m����\eMb;��Ү3s�+�{����y�fش��߯�`�o��}���|��Q!b���g�h�:,�yR��STg<������*��T���2]	J�4��F�Z���'��kB���oDd|hMf�~]�����ž��իzy��r���2/��Q?C�&QNԮ:/�wk�A�H�t+��$�����v�Y��I���,���B*{0���]���m�'GX�}�0g�P�{��n����Х�4�U�q����>���
C�K�q�[gP�m!��?m!��I��C�m<��w��G4�j��[�F��
����`�s2l�#������w���K���/ާe&��a<H�}B�T���s��-`T���7��:�j��9�>�|jYOw3{���ڶ A��wc����2]i�ʥȉH=��'�ը�F�6���A�,���3:��D��C�l���4�FA���̶bȑ��r�~l0i:7�Tp/���PY%�y�HA0R�Rޔ��r�B$�I��hM-C<8���yyy�4���=ޚU?�|1�n1kP���R�k��4M�fM�br�u&h��S���������d�J'�|��.�W�CԤ�T��V3_���t���gݶ�YH��y0(z��neO�e��
���]�Acn��b!�3>-�ݶ�Qp�p�5����'��zhLV���C�C�a7BV|���Q�䋫o9��q����y�8y�y��JCSQ(b�&�T��
��a�-�<xo?����_+�2eفh(\N뢒A�[��7"�J��PjuC8'�TD�#(�ǌId�ӓ(��pT������x��q�KD��l����%�c��<~�^*!΅�L#�4����������w���������{k���?�Q-D���4E�t�c/[�ͭ���I�^��A-��-�P#*z�}?��e���!#���⻿	�Y6����O�t�s�'�"'��m����ȭ������뗊l��H��!��UQ�Ǆ�hN0&�x)��� ��_��Dy~�ʖ�}Ȃv.�1?�f]��v2�̌��	�)æ�����H�|T�+߽��e~Ո�����Zxh�4#� /E�YQ'�ҲC$w��|"n�{��ُ�O��I�q{H���hG��P�&P�b��u��or0M�%<��XT�I�c���ZP�WX�x@;�SSp�}
��	������^#�9�d�c�u��)�0�k�{Tc�)�$Y�o�L��6��8ĲK�lP���V/��Wĭo� z>��n�����"���C���DE����2.X��m�w�z�M������U0�y�HT�:�E���6$�u���NޱWaGC��F�F�9��G(�n�[���|�)$ ց���H;U��9��G�KN>�j��,t�b�R�I;̋_c�:�!m(`�M4���Z4�^��p�1!�АH�8]�rTQB� ���&��ۀ�@�f��-��vO�ꏈ==Ը���zh{���t��.4��H@�}�9����x����Z�Wt����a|ŉ�F��_v���F:ޞ�u�/@��4I9���ہP�[���.�(�|)���k�,�� �0��J�p�1y�`I	�( +��בG-�v���j��a�}(��pD-��/'�ΕqC��N*���pw#���	z�h�<���2;|�F�Mѥ��3#���{�)���e_��#"�`�k&x��
mO���%�uA*_"�����Ǿ�g��s
�y=�,c<�W<eJ����.��/LFH}���O�-W��T݁=`�Ie?�&|��IY(����Ű!C�c���ގ��񓫢(
�t�R��`+���5Z�@�|�F?%b�t�Wx%�C�^���"5U�ak8��=���a&61���T��B�t5����G'Q�?Qߙ�P��7�{���9��L#�e�����HX����ʴH:qbZ�Z�g��GC�B�kQ�j*�����H
Ν����������`�8����ni� ���+�y�s�Z��=]"�6TĹ[qO�^9�/���͢�M �q{��d�ӥ@l'��ң݈�X���=�H�y��Y��� �E��Ko=��0u���(���e����h�l&���K����������.�
w :�J�� X�ɋ��Kϟ�q�q^�Ǫty��̀����^AF$�w�XH~�/������a%Ԩt�ܫ��ۙ�G��A�
��V�n�_'�V�\�]�����E_�4���!<�M =�{��Su1ݨS�� a��2�dxX7�I9�	@r���8��M��G�>,�ѵ��[�G�F��tAZ���HG�`��S���Yj��˺��6�+O��Cj�IM̯}@���?���&�lY���~1��e�l����-B�Mq'L���k`hf9sGX�
o3-yL����˴�F[hӮ�2KYQؾag;�.�v��3#t��pjw�*�7�B��E-&����R�;}n?R��f3��P`mb��gH�-8����K�$t�d�M�ŭ%�	W�ݵ{�^:$hg%���_�jӕ3aґ?s�G|d�,8ѻ-��؇��y�{�e�O
*����-�� ����g5@6�*Y"䧭@"�l�uuUS�O,��;�A�����	ŧ�6QC�iG�Ncћ=#���n��4��]�+��Z�!~Cm��-(%k^W����D �Ei eۨC�B'�/~˺`�?�(��J�%���:���l��'B�d�̋�}��)M�>B��������B��ɴclCQYq+�R���1�xU���z����8YG_���sb)�3t��Y�vT-�'o�Ur����0[�K6{9KzX�QlrP3P N�) JbР���.M��Lj-��ƦM��CH �8x��J5�0p`s���l�x����'�_�.3���NtC7G����W��$��h(�[�h[�����?	���g޹��
��eb��:n7n���U81
�k���V�L��v��VL0x�
��uh� I�0j
��F:���V�pzr�]ȋ�:y88����mE����g<k߂��a�/�c.gqD���7�J��\���j`~��
�����[���
	�K���饍K�kY�$���?CϹ9�%�%>�~RR�9E��B4��n�k���#c���ú��}9W�6��D~��$�A"y4VN� .ק��P`�9����q#������x�}u�哉r�J�h��t�i�#�оd�)�s����<ܴٶ�c��ͳX,�~�f��pY�u��/߄�^u�7��Ja�P���@��	ӄzЭ�^�q4�Ֆ����X���B3�����UOf���tr���f�_��m��E~��9���ϐ	pG��fbc3j���Q���*�03[��#��7J�ؕ�oq-��8��7�o�[�_�<���9�O�`�?+�`�~8r�dJkz �o�#*��E�E��r5��
���8��CvQtf��jSG.7�2B�Qou�֬��;5M�֘ L�8��j <� ��:�J�7�dϏx��&h���l�7�� ���ٕ��ԯ��(��J�U����3��2e��L��:�u�jm;Ŝ�����T߄V ��`�L"���ѭ�#�V�q�?�`&9AC�C�:�!t	��T���)��A%���4�$��q�$�L߷�\*A�9�j���P����C��sQ��\���C�M���f�]$��N�r<����8�)�լI�
h	�Zb�����;�y�[��_c	��1:yS��jE�@2�<�2��<.��(��)~������}�~*B)e8ʷ� #�7p�1�֟�9}C�����G[*=�Y��g�v��%�L <����bH؏)��E1o����?a=y!�B�l�v����{� ��5�+���%l���4���ˎ1 k�*�����sl��E���Sd3b;
�櫈*�<R�BGN���j�_J��J��X~�+e��_fwJ,.$�p��r��+4�,�f4�������fP������W��[�	�vl�q�<��V�A����	�Bt�i�΄G��Ų���!��xF�a��y?�s��lty�̺N�a��|��FR9RSu�2�D��,��ʵN3Ⱥd7�[F��x��8����@�0��������X�n�c�-�г(zo�OJ �g�1PH��c��R͠=����8N�w��|�U�|Ѭ�a�ێ�W�mЛ��_%b$$�s�f���X���u��_�@�LK��5u�-P���@0=����w/KG �ӍO�ؐ4�z��(�D5T$�2��M1�̫m֞?�r�v%s�"�����֥��%�$^��$�l�2�)M�>��~̂5��R2�V�N	ީ�`e�7Ry�]�V>r}h���i�:a��7�{���E��e���w� �-� "v��=E�[х;3zG�D���;����ճ��
BqO���#��3X�O��8@g�N�js(ʟ�JC�1Z�	�7;寰@�ɱ���XʽB�iD�݄h}���9�åSF�4��Ⅼ\��#�@Y/���z�3�����8f:H��ϡ�!��~ʂ�u_��"F�M'f>��؎b��i�g?n���� #g	�Cu_�N�"�rJ\~ �=*~��w��97���z��6�ZB���۟u�r��$�U�:��3Jփ.W�3�\�2���,��2�+/��
��Ąd���T�Յ_5�AF �ٳ��ͺ�7hu%<U�ی=����ir��jU��!��K��@<$"�q���� �Ӵg-�c�d�b�G��b��+�]j}��+dc���L�[�dx@��쾂���P��X� �G��S���$1�佇�����\���}�������3����_1�"��6�P�L�����`�E�<���e��ڸ�7�4բ\JODe���iu렸��&�b� e�1��ka�nA�|�&?T;Vׄ
@��<M��K`Ҕov�L�&jy��4�����nk��C#�k�h__����ƾ��m�p^�����׍�Ҵ{x,��ֳ�Q�h�ʎ��-�����d�1�X�j�Z�������N�'�A}��&�ec.W||>w3�R�}���zg����;Lˬ����M�II����Ey�� ��D�~Ą��k��z,fJ��t�F��}mcه'".35��2=Ői��Jݭ�Ü(iƣcz�j^9R���"W��g��7n�C!?�|X��˪ ��:���"�)a=584�Z��6�LR��;���nU:�B���J^PRu� �W�0��f�)e�Q�0����Wl���ӍPE_L
�e����3X ?�!�_un�X?���҂�VG(�_t�3�R9�x>ue��Pb�!�Xp����3���� ��n�k�ۙ$�aWE�=B�R-J.!�IFꦖ��{.�&�D��3��C~��}�b��c�4Kf�:z�u�;^]g�|�ڣ��~']�L|��H����ɉ�C�I۱��)(ׯ ɵjҤ{�^4�9�J�򳣥�!������Z$_2���@�)P��������|�Z]�������{p����ϯq�Ŗ�M�b���O�I��5�T��F�H�^(q���ϥ>+yM5p���f�:�	%WZO\�]a�MR	��(U�	�U�5�p�
9���3�	���q��|��:�+K4�	[cO#@3xG�w�t�=m��\w3_خ�Gܗ���t�k����c�pYb�����i/�y�g��#�x��z�<��K�]��03%�r�'R�be�p�g�M�8{S���'����9%�M��fH�� �֒��.���ᖏ�n(~s��@B����ъ�P!�00�;����Ba	<匛R��b��x�M�T:q9�ܢ��I&���/?�K���<(_�-C�Fn�� �������4!�$t�sȆ �wn�
R9l<+Y�9P�Pf�����nY9vP'k�n��k�cy�в�s��h!��&�ə�L~��n+#G�WЈv�>�����G�v%8��P���w��|���W��8�)>�k
ڒ�1KP��ת��z�um��s"�g��RZܿ�J��=d8}Y�lz�`�=-@��hT���H��c�"<�&A����/S�Ks�$�.�C�B;�ck�՜�����JѪG҇ɶ�(�Y¹��K}r�!X��+������$�Iԩ[{��>��5.m��.�c�����١�����|r��$b�/�WˬYU��w���1�f��|%RQ�{I��K����EJ^�*�uȹ�#�� m̽��1��u;)9���
�{2�/X��m<�h!w�����+�C���s���*0%�&�̪EQu�ν��3����M�	/���}��j$��1ra���Nao[.���M�������PhS+�Q��*��F�^k!p�	�A��Bt�)d���e��2(>�/�-2u��9_(�<{���Q��YLp;���D?�j��zt���=��������b%eD^�c�����a�w�{�<���_#���[�xl��=]�v�p����+�V�䜊a��9r��g+�7�ZO��_��*Up�~9q�M_�B���ݓd�D�Kv��e�"i\st�&)����V=C��=�m�0:�4��.N�_�X;��8�f����R���[�
(v�L��]�p��L��
�x�~�N��Z�&UGb�E.$>,����sv0n%m-gm��@⓺,����4���3�1&-�H)<:&P]F{�E+��yN-D�S�K�r��!�T��4,l�u����Mj��uҼ��L��b,=�CM #�W�p�ę��-D>�9V�H��M�s�g8�V�)���A�0�r9Ѝ<\"��2��O��2�M�kG�f=쒢?8����yn�9*�@t�n��<���1��~��&'���fʹc����Yp[G¡�j<}�眜H�e��.!��ImeºU�V(I<�C�����D�c�vU����8K��uF�6�������i�x�^���
c2�U:e7�*���f�
�ڙg�����!�Q��v0:Ğ��s��f$���@��w�3�/$� ���˘�G�oZH���'�V���H���d�?���`|��@�)��aд.��Ǟ�&�R�*c�������M�b���i=K��ms�V�2$o����跑f0i��1$E3s8Ĺ���=�Ť'�kJ�!+��G�k�&�;~���]T������\��a�m��F(B\��8�\71�%�yF�-P����?�DG�dO��Z��-��#����1UЪ;��zm��Pqu)�����<�hD.5%�h�t!!{�Se9Xq�iYj�ゝED�80�c�6:�0ig\���nYJ��`B�ƭ���9�y������k���u�(��°R-��zU������
[��0��Yփ@9JT��p��R�J��H}F��������[��m�����bg�6��C\���%�D��4S�CE^���|s��Z�@+�<<��8(�}u੣+@{v"��,z������)t���$�~F���2���{߻���t�8D�� y�y�$6�nW�_�}f��*F�7� A���z�^����9��"��ܔN��g�F����x����gω���9`�b~�h(�m��ܠ��	�3��tB  ¦��=^�-�Ń>�s������sw��}l:�\,�{E^@��T��2��v��1^��o������U�U��zg:x��z郑�����RQO��-|Zòln�b��o��U�3��/��D=g�*§\"�)z!�N�}@;(y��LH=�8Gg^c��[)>��M�JL�Z��`y�R_j#J8c��/�-a���6g�\���kj8:�&�y����?�+5���W~X=�l�,�}�
�*u�*��n�Jz���[�$�`o��]#����\*0V8OFnx��>0�K��'o�����pZ�n��8�~D~i�I]^��/0j'>XhʔP=�w*!(B�q���y��J�,-9�WI��;$��_�M���ڊi7k=s�P56i�~w��HKŁ.$�a�E�P[ p(��j8gM����c.kCk$)�E����#��K�biB7�m|J��|��W5�:���C��5;YG�=��g��ʢ���Ý��"'Y�UӨ+1�o���ln_��F���`��q�,~��F��56�EĔ�*	J�����f�A��^?�GH�XC?�ܢ욭#��� ��u{�7���04v������۸ˡ0ë-���ڱ�����u���ǀ����w��qh�b(\�q��q&[�j��-�I����D�3?X��Jl[R&��|,�ss1�ÐKG�9�8�ٓA����{��.��ߔ^��jo��)H�| p���`���a*����2����h�b?��=R�,`��֌�B^��̤r���I�|�f:�%룂����L��z�g�Nq�:X��4��g�(�s�TqWN���<���ܲ-d#� "���広I���je�>���|Q� �l��q���yQ������c��\� �V�,�8ƴ��e�U�E WtOC��0��_ '�N�F����@Ё��B��s�n�)�%yT��q��9�Y��= D5�]�'g��6�� ���
��X�E沉h�������1���fPe���� �.���;�	�ު��O�њ�6+�P�����
Na�OJ<EB��<U����C��	(�:���z����a��/۪Lhi`u�l/��n�2�π }e[J�JKk�h�G'�.�Yu~Kie6ӵ��M�� �["	�ݩӫQ��qKu �H��A��K�%��"ړ�]N�Y"�?�U~mz8~�	�mS�Pއ�P}-�r��Թu�{m(^�	��:�6������5#�S�Y2Dh+
�]��.�ԉ95��c�]Y`o	Mt�4�pk�?����L�a�no���,0%�f��Î�(nC.dm^7ј��g�����g��F���7eP�}b-}Ry{t��*V�2	���J�+�n�m{#"^IU9����BbD�H!�$���]x��x�bx��̇*Ο�4܂}�։\��n?���@N�uQÇ!f�[�A�Oݠ���p������˴�WTU�l���8��bɻ"*�dd>-P����[�#܁���$���k�<?��
v��<��g��3�kӷ��R7?.ei�F��f�QSpj4"X²�R�+�����_�����pU^�U�ImT��8��o�]�Z*�㚅�~d�y��Ae�.����BE�OX�G	�/�{�Ml3���Ni���T,�JDРP��MOv �nG>�y����4h᠉�R�1�@vǳ��U��C�Tu��RZ����3ĊN��� :a}��������$��r�1�8�߾��L	|��k�'���$I�>�N��ƣ& ���D��bב�W��~!�o}pk���/ȇ<
�|D��	�n��Ý8ۻ�\첊�8�&g�h�*>�Z�����ްʢ�PM�&�,O����y��v�hn�Y�?���%���������'���3�U*��!6�A
J:�M��E~@`�8�s�KJ�GtT e���i�N!�L0?q�Q{P�GN��D�cRr�^I�@����<7�^4��X��]�BD,�Q^)�((������0|Ϥو��O��'s�7�E�)%=���"�2�i?�r$��<���@rW͚u�Y���V$k���l�  hd�O���D�2�:����4g��{�s�&�ðظfngqc���ry�]�It[�����ޕ�  h�~�rW�2��HzFz
A&@������|M�I$���� �(�]�پ�H���%�if���&���v4�|��`��u9ڇ,2>�j.aKm�FEJ�8\ӒΜ &���s鲿� uJi]��W��+�b�;&ߊtPY�����!g��|g3O%����Ɲ8'!����,�$�m�D��o��������� �T�w@���(ҭv��>c i��7����1
ӫC3HՐuNxW�@�S��FC�u���&�����vh��Dm��U�=!�OW�%4�(~������Z"��h CK��d�����t�?����ZMK�����f�q����q�T��b1���ӑ��Z4���4aC�i9-����-P�q_y-�͏D�p�c��Hb��ì�\<+�����4)�D���^�cRf !t�hn�u���Dƥ�\]I�A����jY�%~WSm�9�t#��D�4�+.�|$��N�+8�	�������wor?����cc�3�'̌��:�b�ꔋmPy7'D���
�.��l����&b�0]�g$�k��}\���c��R�P�xPzӊ���aq�Q�6l�܃o�؂@֚`�[5�e6Ҩ��^!E �M^�+�^Z1�c_�J���{�/��Ž���"�&��2 ��S��j wx��w��N�A�~�&&v 5��� �����RL��;r�5V4���@9k+��V�)CUE{����b}�s�I��G��#�
y���2��!EH��E��m'ζߧ?ʀ���>Ĭj3/�{��μ���׷t+	Z��xxZ���p��[�a�hݤ޹��F�;�+>��;u�m��zJ<��Ir.���׉��oɜ�&0�~^�Ke�B2�+��{$�ޚ�ls�	HHS*o��Z��j5�h�[)�;�Et�����t�һ$��X�̣*�!�̨��3.q�n�1�kB��҄=�۞V����r񤅔��=K�u�B����`�'F�r&�
C��.Zk���.K҇�^��j��"�ץ�y�@8Ch:�3�G��������^���}��ۃ�����5��n?�J�/Ŏ�<ރ�m)����k<�o��߄����-�弤^�ؿ�U��!Fz��������Fj��T@�NI�}X_(*���"i ��v�� taD����?�������z*g������ӗpv�-�I�P6_�Ð�9�2�|���?�|j����n��}���[W��x��L���� f=x�����O��Mb�}�B&7�ZD�@�-tA�M���� >���fl�Xң<��Y-�ȉ�f��=o�����9V<��/�g�
~'Lnj�}N2hD�.�#�YjkX��,�ӈ9����~L歖���O R�P~��4�a|�VV/�<��A(���6�fr{�V/�@v!�p������?8��F󡁃�K���jq�8-E��-���;�K�G�K#MW�c�(w�&i��#ɥ#�;����;��?s�gZ�0�H=m�z9GF��ͅ��޴8���w-Bj����U�Y0):���a�`��3��<�`� ��gܑl��F�|��A�j��L�����5l��㸒aۿ������}x�b�@U�[�7�ֶHlLy�c��	�7<�a�G��,��C<��fgjJ�:C���ť��n��.@�lJ��Y芷� ��1�lxV��X���}�	��("�i8~��u�`��}���z3������\�?��N���V��V����"���k�����ܳZ��؅J�L�:�l���*7d���H�}�P���@��8��n?s�H�(;"��;�:
A R^�6u�"��	�̅����&���8���ʉ%A)S�<u}MT&�ɗ����
�bq��j"'H��=�W����͡�����Y����x�V@R���|�	�X�r�~8V������,6����T�!�x�V��(>�dO:b�w�"��R��j��8;L�����4��.w|>�[�U�����eG�������D�<{��m z.>�Uf�Ҭ�1_��TJ��\�ʶ!��H_�C�z�!�]YY��O�
�j�����·��R�+�<���
�Tci�p[��aCe\�����������2��� ?�Y��U|���<�����x�Qu� ��p�f�g��@�l`iǲiS2f鈃�R���u�"��3�	�����Y��r�Ҵ���R7�x��-D	D�k���2��#yWG'���q�LrJ%�����T&���~R��9�-�����y��G�='6f�/��3s��,/��N�T|�-Y���6��c�o��E��ˇ����\�XL��+��T�,���0�l�?I[�3 t1� i��\ci@��@�
!�=P�] G_3.��-Ҷ��?���s�97�׀m�o?��wъ�r��$�A1�?z���/\6��c��3����/�k�`n��g���R{|9r2yw5�F�(97��2���n5ok�хu9KqҎ-�}���s9�\�+��ңj��/�9#��vwO�:;���]�,4��9���)LkAL.U��i�y�Xz9~0+����MDs+����L���#�j����q�E�M�i�#�q�Y	��=��iu��i���e�Q ��R�Mh�݇a�d�U��'~1,�[�ؓ���'V1(���׹	�(I��e�i���ɔꩈXi����\J���9���v߶�k�ь����Z��{��q<�-�+�T�@��/� �h���C�"���K��!��Ky���F��%���1�ᑖ�'.�,�� �Nv�+U��ԥ���^�?���:0�90<����7aP� ;z=
^��p��4�M�:�#Aĝ�>6������	�����g����z��N�b!Q�P%1���[�j��xk����~4N��r]/miv��&����V�n�>7�W?x���/�A��]��R=���R�V2���44�Vt��հ

�Fd����E�a(��Y�»�F�=����K|�z�=�|��ɶ�i���ǹ�w�T�;?��9�\��̿^*:[��g�)D2���ovh�;�͡�v��V�n���K��$�;;�,�n(Ti�E�߮�����/�O���]M����j��^
V� ���^���ۻ#�l�$��Y���_�t6F��2BN��m���@*w"�]<6�ސS���J�,K'`�?"�mM>v��q���ǰ���L�]I�=���
|����U�Q���-�t{lx�d�#�[�+cO+�[�.�2ߡdiv�76uɊ#g�/�l�7���m���E��:�d�	n����\#�8�|5���^8sL�ʡj�x���l ��8�u[[��Wx!�,*?�s��@đN2UK�Zq�Z�/��OPq��u�	��:��(Y����&��]R��/�q+өc�8�Ot�Y�SUyi)s���+�z+��������+�����!��˗�U��g��`�i������9Mѿ�EI��n��^���@uAY?PA�q�rOE�n;j�}�a![�q`'}�s�[�Ȩȭ���v�:k�H=�-�݌��C�G^��x���u#H�r�;�I~�[#:J���ٹ�G�~Yb�om�h���6�)�9?��C	����U���;��ܜ����o����(v�(��U� ^h�Q��Y;
>5q��^R�e���uO[>��Z`��x#�e-R�WQ�k���S�vΊ5:?;�xq�&�u��f��9D���õQ�0d~ةI�d6Q�IJ��[����H�3���-AIN��րP��>,�2��s_a��Zy]4�Ү9c��������kE��:\�r����|H��)f��C�k\v9Dɢ�2��^�p0���w�1���-,n �f�+������:�%żs�Z����i���D�S�!��~�����ew!q�,���x
�lLkQ�ʈKQf�?���n�2��.}f��'&UE��gb'm\�DFC�cG��ů�l��r���_�R`���~��Q�!�0ﻇʐ��1�*��A�O��B� �9$���z&E���W�Y�~�,�������˛V3�)���!k�Nt9�`��mu��XQ�7�jj7t\����b}vZ�Qٗ�+E��lپ�he� �(�V��H� p�+�
�GZ�5g��YMu߈x �v����s�t�b&��8z����4b�I���ݬ��Ņ7�)�VK�k?}��H��i�=PH�+�z��M�&7��߁䬼�.9Ǔ��D���[B ���e�NuR�3�}<Yޞ���mۖ��Ul�5p�*�-I��A�sp�]*�K�4�A��, s�Ͷ�k,�d�Q�4��;���m�s�%@.��% �#���N�S�ݟ5�QNr�%����^�W.��Ā3�+�XAE�a;ɛ"��W�n,�qG��/q[lL榖�k��1D#,�uV���0n�kVUx꿲��e��)�`���<�
Q7����E���l�o?��(�:��z4�h#{��L�M�{|���]*^�A���s~y�x@x�'��h��[Vrr���`�e�rd�v -������""�`�L��x+��I�snPN�Z��w�a����y�5"�0�,<C<��S���t��\�I����I(���[�FF�Q�.3�H���1����[�3���c�B�kA�Cn�o�=�\�E��=a�%�`7������dc��f��}ٽ�>,�&����G�V.t�t:�vݔ�j�����hs���Go����9��?m������t-.n��;�-�7�'�@:��Y�4�Ci!�ŬdOHBg�)������&�uNI��&�j��0���a�.M�	P�CB�j7�]�}�?2�l�%K�D�#N�VTqw ��.@�n[9��0����5����b��
ۤ�X7��(��r�Y �Ůl��'���ҹ�,J�"
N���R����f���FIK�$ލ����q��p���pn�N	� �����8p��HQ��� q5��GpEfX�����!C����c<?�C?��+���v@S&0O.���N+�s�/z�
�	{SI�"�B�,h!w����s��mj*׶{�etX� ���;�B#2Zɼ�Γ�;Ͳɚ�P~�)gS�Lj��|ֱ c|�R����U� )l��0�A��V�f-���[�m59�5|�yQ��JJ���Z:���J\�G#Fb�xY����#��ۡ��Wď�P	Vc,� οrW�(�Z�ԕ\���{Ű��5��ٯ�YItA	�4r��2��ȁ�(�u�p`ey����mu]�8�,F���d��u/�����I��|Q@�l���Vz;����Nv:���`�=j��Fbxs1%x`�D�e=�����Z�fz��!�6�"�����*5��J�����^�3£ƌ!3���cwi�T��v5 թ�+�I�J>y�*3GcV��(�����ѻ���Xh��D�^@��/fK��t>��(b��m
\~�?'WtmSn��`럎�� P���C�?�e��>S��,���W</�I�V������
Ѳ&��(k� �w�͗=:E(�Ȓq��Y��p��k��H����9�l�;�Y��l���'�Ɍn��)��x�� ob�w��c�:z�e�06O��<v�fL(}����c�2ކ0x`���sL�½�a^�P��"�p�5H�_z��]�9����4�ё)�q��k#����
CN0s������wHq)"��ɭ���T�<���h�fl�BoX�ȑXe�wT]b�D�V�
���-T��6� H91_��N�b=�`���}�gK;�?�;���(�W n�!k�֌q�#*��;S��؉{����w�_����\{0�ԟ��yE~�i�ke
ְRsZ��z��뭃���������}�12AﰽB#����^�l_#Z;w�����g ź�P�s�O��i[n�����۸�~��ͭMDB�?{��&�z:�}S"J�^B�8�9P��]�G�Rr�=�����y1"�5���?��*A6ןK��#�
4�K_X��J.�ˈ\�`R��J��������Pb�s��ɩ�)����?�Gj�����a�\�T�@�I}z�i���]����;��"3�n_N<c���:�(61�!��R:<�g.��n��c��]-g/�W�;<4���,�U%��9aϰ(���84L�sV��m��/�[E�H(���g>�CC�;�!������#u�O�F#B5L�^9$��:Cx5����1�����L�+�^���m'��FE_q�l�w���I�An�U��O	I
8��l�� ���L�1�v�m�H�J0WF�Y�݂5�1{�g�
l����=Ί�fm�w|z�qZpG�ɍl����Q��(��i3$fH���e� <�x �1)	���3,�p�E�z��4� \�A�L瓏�g��yM��\�!��{�~ÆU�_�LeBh��.ѱ|HP�%#�W�Ap�TL�`����	���s�!�k���2���'�^j$gO���l�S$��;L�i9cimf�#J�G��*��tPv�K���U/��hb����t��l�q�ˏ�1� +��g��	-`PPՌ/;�P�^c�pz4�~H;^��!�q�y_��w�JJ1�d�v�j.��}8��y��	��%d��;��hy�*�x�Ե�,��'@TQr��_�W�֣BE(��,�S s�|�L�Y,R�V��[��x���I�;:�B����5U����?b�W^f��%S5�$)�jIN�RE~�$���G#_s�s��
Ő6�H;��[�~!Wn�n�+桩�*�ׄ�ģd>��ʗ��_��JY���9_>���F4�n���:+�k@�O�bA��˚?�̳*�ID?=��&���mQ(C���2�+�����)�>oc˵$��
�Q�C��������M���Ib���^F��m��y�)�j5�-��D���B[="a	���  �[f���������j �,�Lq?����&�����pu]Zy�7_������q |���-���&H���,�=�wx{0�%�?�Fʵ��O�Y�zJ�0��F��ԄKАs��h�ʖ(::���s�B�Ush�d*�˧�o� �Iq��5�|,��XG���qd�NgK��O��3k��G:���{�hP��b"m"��Б��V2hJ�
��4�K�x�	��wmX�������+mYa:<JJ<V��E}|r���\Ӳ7���ӆ�o6�(+��?5�Nc�$�e.�ON!S~Q�VŷS-=��E��Ԙ햹3%��r�2[ѓ�ȓu��-�k�'�t�5����:�L�~�Q%�9"#~3E�6-���t]�:YT��$"��K��2-�~�'�����O��c�V����x��$�'�
�u��B��|a>�\Qu�*�2�ɩ6Z�[-}��� 6��|��r�u�=�C�1]v�Jw�v��G6Z��Q�Y���H��c�����#ݛ`Mx��L��8�n5�nD}i�c�?�ȑwj��-�\�#�;9�F��`���Y���TSmG���+�؈N�R�{Su�P2��*.��m>��ݒ�
h�©�F?S�2xS9��u��)A+�G)v�$M�H�/�'�ESL�d�r���Dyt�4>�]�˲s��W�t�o�2b��}�������H����lѐ���0��n���d24�g�

(�A"�"ĩ[��Ո:Х�r������ǈ%�������P���8y���Nv7"uao��ÿ����N&<��JY���e�3�z	W؈�4 �L�*Z��u��V���v���2��`_sۙs
U|�+Y�������Qd-J���*��iU�󝓖��d� ��?t�i�/r����b�Hp�6P��9�6�9(Q��sv�"����fxQ*��u�>*��L�`X���1bd8��k��8��+�ǀ=*��+��T�?8!μUQ����~V�����c�?b\D|�l�:fq���\��W�IsF�\rn����"���h�u
��h�<F��/��5ˡ��=6�W����6���Y�L:H0Y����6��/\RHf(O�6}��d�Z��U�l2���f�GNk�4��n4��X��!I��d7z��!�胫��Z��P.Ɗ��&�ĺ���ɭ�)Ih�V}���� ���K�h+�����<WN4G���^�]<Ĺ濿kU)oJf���
�Vu �k��<�U�e������8��	_8*|��J�7?����7�.�̮�`^�C�w� �-�$\�_�e?��񵀘��\���Yv�yR�.��3Գ�w��C�14`�6��In}�N�DD�S#�"9P$D�e���|1"��2帚��+��n��k�G$/z��9�
	�AP���mϓ+��64��e<L�\�/���/�jI�-'~�J�ꕡU�,4C�(��uV�E�����L������tdG	n����{�:|
��] (G�ߚLU��4d��BE~$�ԯQ�.�9�ke-���B�9I��~�0N�rX)��S��L�;�/���X@��T)�C����:�������s�|�z��|� =��9�m ��@9�7:��嶉-_�7��2�@R�e��W���Z�W>�Y:��@����J-��Q��/��'U���@G3HU-���$������	n��7�i]ԃDZ<p᭥l�텚uo �y��g��nFd7�AT���,���mkL`Dr��Drj���"��A-�v�r�
L��a^b`���?,�߯�ʴ' |�ޗ<��vj����n����rj�*|�f�>�;�B�_GHk�T��\i'�<c���_d̈�m{���<���	�"Pi��b��y�� J`䲬�K@^��.Dh�)�Rm��H�Zf�(*��_�%�������[��`�&���EYJ��wY�<��t�
.�"�兹�>o��wc�9�	a��.�yu����*�|�0֋�k�􅄾2E����2��h:� ���E'�J�k����KC���Q�Ax�ϕ^-��c�(F)����� E����7y�F
mJv��|�B�Z��aq�(�匳�����B�N/�C��k�P��ٖ}3#҅A��Mh�$!�A�E|s?�Mv�����N����@�nfnis�)FYB�]ySLeHԬi�!��緙�J��2!"���J�~��~o�r�J�^�̞��Ω?����R�6[)��������a�M8�!�t'/U;k`�/��~J� �`���Q3@��LG/ªf:��f�x� B=�.Ntlx#Z�ތe��r�)��1z�w�}�Ӫ�{ekpǓ��oƨ��bf��A؆������{0���Z��l�Q-����W^��\�τ��S<��oΕ*q�o��`�n�%T�-(�>�}��a�z��e��;�	���I@��~A��!�G�p��tB�õ:�j����F���q�7r��'�����9}@>a��2'�%�K�����ڤ�uڽ:Z�x���GX�9Q��Oe�ڮ�C�����j�,��v�z��a$%�>H}�|S�%�::�nQ�V��[��I	504�٘��l��7���4o�I:��NǙ0 &�s?�O`��G���?`W�����@c�E[=i�#� �d@�j��G��KX� (�mv�x�9�n�Y��).�I��2��;xoK4G�j[�:�zdcc��U(��L�7��
���Z������Ǫ�57��|mQ(�jge�g�!_��{L��#�}�ԡG#��8�m%(cL"e�i��>T��,�ڸ��L'�(N�s�}�Lu��!�z�ղ/���^O�����
j$\|��^���P[����KG����ن����4� ��	�C�=q��f~9H��5H(�jn�$Ѱ&�X���26f^{�K��Cy��L�^���F����3��G=��53���`��g̲O��_��H��q�zJ�j�ˈ���C���A#H2���}��*�F��6��E`����Z��tݰ+�/���Ȝ�ȷ$�u�7�R(Ě�zO���ڋ���c*i��g�x�?��a�^����3#�lc%�����[_�Ȝp%��| j��+�����!��ўB�
4�n��3��E@�V��Ty�!��Dl޷�d���=�y`j�ٞ�մ2r���䝈'v�>C�L��jT΁�	\�C��A,�Y�:/�g�M-�CI:�Z�a �b����O}�pТ+��asj	���%u�(�'�p�.�V�A�	~���^���������L��хa�d$�%s[���]U�.6W�������{
�׸j�ŏc77�D��7q9U׺�QOi�ds>��޵t��q�@��F�RQ3���ր=��q��<�$3���о�E��EA\9,u���E�%G���M��k2��[b���^2���I$�I�H?����H¢5:��3d�6��d�,��q�C׫�g���4���X�o^�@�3#�ߪs���׻`AP�š0�6I�+�]��� E�� �	DU�SV�f��4C�w�zw�{/_�o���&�S�`�|.=1���c��O��<��+H��']��W�Οsؚ��J4�؛�G=���I����)��@
�kU��sA�?O�\-�:񭆓���m�=��1��',R�;)=���K5�R���O���O�G���V�Q�^�R���|B�K�ݦ?��3��گI�ZMZzڃ��,x�ظ��]ZH	�oV&�J+�j�T[	�U�1�3Koh��L��-`L���\#���dO�+x:����䌮��_l�ꉀB�7�3���ή��{���OS�V��C�C��*P�m|������G�wJ������7=\y�����r�5�Ct��u����ض��\-H���8e�*�ar���M�>>߿Q�זiP�W��|�A�@7����_C� ���n�]��gnM=8����[3�è貪������ -�ĩZ����.���ҵ��vg�|��̺~�,�q��/{��4�F���A��2b��dm!�jOz��lZ���,�����,����u���������|�쇘��g�%i���Gg/�l	���e��ͼ_�����5�s?8�\�Ƈ�ݙ��݁\�RZ��a`�댂�MM-.��"��N���TiF�+gS��T]��&�m��?bI�X�{�QN9s����(��3��l�q�~`�C�W���ЧL���m��S4S'E�l&��h���q����s�ip�o�����Kt��:'���a|3�y4�2�:�� �1	>t�EZ��6�����M�<+�Kq��!c�FԽ#&����ᴟD ��
�G�fJlxLS\�+~xK���xo�p��H���QD6��]��R�����U�Zp�|6�;�K���⴦�.�~��:����\��;!Q���w��WV��x,u�(@��IKk9�W��M�<�m�*�0�l@���H�׎eZAG7�^q�p֐)SP�kH�'[^���aJ��$V+���X��S��*qD��P�~g$7�Jk�b%�dan@֟�h��u�]�Z)k7 nڝ��J��u|@h�`�t�4͔���8	��</a���ԁ�H5i	�mwl���6r)y�aR;pp�����B�硏�U������6��zd|���,e���O���كݤ�uy��nk�$Z��@8��2���a�}}�ԧ(c����U��\�$��q�9�?rv0K��K�c�B#�k�^i��쭻*�2�y��9I��v��:2o��q\�Z���d^�m��T>5TF������S6>���b8J2l76���q	%��*ժP����ҢL�`SW$����$���mj�~���N�vK�p\�."P	N͢d;�ۍ�w�|�_7����%ښ!��&�D��f� ��\���I�����K䴽����R��l;��f*� ��gtҾ����[vvݚh� �+�y���qY9����%�;����Q�;���}ѭ9��;�=rt�S��'8�?�r�3��0�K�f�n��׃�דe�iXa� �F5[�<�$�h�S��}�'���`epG��d//4��G�N)��F�Ǻ�� :es���VKT󼀛�U�p��4?�_�6����k��A�3�sv�0�z����Х��_�
<��xc�v�ϡ�d!+(S��[��^�y���B��v�ɐ=����7�0��~�pHf�V`����V���k�)+gs:%N��z��E�[5��9I	mH���[��"������&�LSF�N�A2��pc ��1��vd�j���L@�@��z������=,B8��Y��_�P�C#(o^��#y�-��l��Xy��$
Ʊ���A��UR�2G����3��xs/�m��З��D'��ƀ��)��5���5���9����3�_���B��*�c�o��~��z�t�	����O�X�Ă�c1Y� O�h�����TI�	��h�������S�!V���MH��i�����?�U��?Ŝ�$�=��P �sPl�V1�ekUI�Al�E!��$K^��p�Zn���jE�ri� �y��f��2(� K�\��x<�"z��.결��hQ]O�2���a ��������F0�!A�a]�˦
�)�I#9����}�]�aE������/�����y��Pr=�"i�M�'ֲ���jЦ�/���˘�</�p���Qaz�ܲ'��lSzk�
U��r�Q�R�NCU^�SԺ�RE;:<�􆪭J֔��Xp\U�J���\),a-�߿�Z��u��c���2E,J�2�Pn�����k���E�T]���@l�����#<z��V���y���k�*��<�qEoS�,nU�^=��
��
 s���E��#l�z6�1X����Į�]�l��ϕ�1
&Q V�}A$��U�^����A4-���\��u�5�L��zԱ7��ƻ��p�5����6�Q���f>b޸�$����GR�l��3����	��'R�_�1�
*2T?�4e��3c\\��R���t��(��ɇP+Mu���/k�I.�+�<�%Ѧ"�^2��uJ�&�r��?��Ř�(ʲS`ۡ{Ta�i{�:��sp�Q�|�L|b�%��ٟ��� �����m�@E��<��Նxҕ�����:w[{Xv�{ȴ��l9�jwAHƲ�- I��&9N�=@�g�]��>��I��Xl��0=�������i��*f&�Q0"
�s�x��;���8��$��M/�Y�&�Y��婔l�.Y  M��v!��N��r����=#���?,o�q���A�������A�� m������^�ѻ6����M�[���+5��r��_2�>ժ��vp��H����A���Fʔ���,�]u�T�H)10Q��q��������Xq�NGgd+qt&:��{|�&�-R9nKM��Ma���O�q7W�����5n���"7�1DSu(�f q	���f�;\O�Ds�X������jr-�L�4�֓��|�g3Eg!����"�>S�F���_~��CQ�~	�9�~�Q�!��Vc�OY �k��dY�"8G���Hf5|��4���gר��J^��#p��4n=
jC6�P4"��i6ᕻ$�6�l��fy��#_��a��'�>5�^�u��%���5�KRU٧���S�$��b;I�_Q��������iн�nH�x�x6[$��s�[~�ԋDG��G��R�3o�z�`~t$�'4$�8ѓ�dߖ��á"��Ⴎϰ{��;�+x�c%u�J�(z�t�^al��m�¨0��K���!�(b�<��e���O�]�oM��"+���x�"16�֟���6{��/.�3�h��|{K�O��\C�at�������H���j��F�ᾘ?���8�	YN4Ů�*�VW8��'��4B
�D���Y��U��8[��%�����S�����Ǧ��H�Y8��U�}��i�$��6o|���V�yv���_7���b{��Z�l���q�����?UA�}r D��_S�#�Fv�*�����x�_�}ST6 ��pH�z�bG��j��4T��U����r{i��:�	9Y�tK'�󭈲��Kub�!�{$,��m�����ēx���Y��W q�1@=ݟ����7�0�-hx�W�`x������ ��]�����F�Y�/
` ��{j�I��%�$h�$v,Y`<�i鈲*-�`�����U��k5�)��PC�����#Wnbgٝ˟8%�KE�G9�[]ڒ>+���MP�h���ݪv�z�|�7{�)K�9-�)
B�I��mJ�ƫ���A��,�o?�F�b� �8��%�vN|?<N+3�B��i�mE�ex)�w�9������"_�nΠ� �AXc�H�����S���;�9Q$y�?��m�w���D:tg�Uܹ��w�.�Y��@{���4{!�*�I�ܟ���ŷ���0��A�NQ�� #[�/
E��ho�|#9^�T1I������l��IS˅T�S�h�%_�l���w�cǧ;�3��!�M��&����W7WZ�=�s�ES�5\f�^�����[]B؆�ց�vwB7P,yk	i$��=��v�5�@RثR�itf�z�C� ��F���/��᭢Ⱦ�5$%�dF ��5_-�o��_4�I���4/6��B2Q�2��ϥ*��j��Ux.��!N��Y-0o���������`]U�_)#ȫM��y�T*&�L�4l�vؚ� ��v�Ny���x{a`��x}��Jg�+��;m�o���/����,췃�*0�}ߖ>"����q��`��V�����������UfY^&8�*l�~WV�#	������+��dN!(*v�M��� ����3��u�b/� �P�Z����ǘtu��jx���*�F��J>8V:��F��{^��h���Ս��h�S��.�|0w��*�U�R��f��l�^�ߟ�,.<�m�6��ƴ�3���������Ò�;c7��1S����h�i�TL�S��7����6����0vR�0o�JIr�6r�F�.9,�.�%\f�������*\pࣼ��K2p�D���i)A����y�/����p����}�Vp�=���0�S�p�>KE���0�]��6��*���Ȫ��ȭ_�����AGhNO.��I�nk�$[AI�ᮿ$4'��v��Gon��08���24�Y��cμ�XEǤ�����w���E�2��J�b�hz�\Ӎfc}ΝJt+�]����w)�?�y5�I�%Al恮DC.���!J$��"���!�`�T`Z�b<qE2��B�n,��H޵톧dO�w@�B�ǩ����Z"�i�s%�+�؁O<ܬ�ש4�8&m><��������gסp/��0�?���\i�{�u��ڈCu��*�P
���SŌ�aHI$��cӲ���͙��� �+�)��Z�1�mT�Vn�*�yX9Z�|o�SV��ȳ�lP{�KJ������+��=�/qMp�栳�YU������:ƾ!=�	�����HpeH�VP�j̬1�U&KaK�z��_u ��t�?�z۰Gm� ������k�>��EбG`��/��_?��a@�t�'�܌#[����X��)5���0�"���D����q�U���R��k���^�ەM��-7���<�0��6_U�ɸ$mf���U�a�/���
��*�S�V��)��@�K�g�f�H�7�B�p�.����!�ʷ�԰��`=8aϨ������[з��ٜ`(�)p���A��c/���8d'�i���R�w��U�"ba�k{�b�Q-�f3N��Ni>~��#Y�T�O��.�R0�u�`I��˃y��%
+ ����ւ� ;��r^��Oh<:v�E4W�o��Y�^��3?��m��;�������j�r@���j�<ƫ#H0x�ܨ��}�O��|� ����F#�gh��1�`���R�ӿP^ҐvT�v:����z"�	�LTƾ��0���1��u@��Fs>Ǹds���bE����X
#O�� u���+�߿a���B�_զ��D��_���M��C��S����E�6����}�W��U��Tβ��MKK�;� ��3�������a�]ӕ�:P�^kǷA"������ $G�K�&W�9��@8�~���dO�԰����;�%5s�2����M�;k��e�������N�����E�U�^qpH��[(��;���	� oQ`�&���%����>r���,yY4�������*u���S��o�C����L�î ��@��j�}���)4]�b�� Y�<���+}	:���cg>!<��d��w���j�i�5�t$t�D��L����ܐE�����4�#U������>���v��t[�e8�,��cs�f����:=#Hz��pa�s��+�d$�zddl��.��kN`�X��-z�A�}����0\LD���F��`���rh� g �A�k�����ε/�#��.�06#��/��P6,Lں眂 G�~�_�YʮӪlC6Pb�[z]>�A�X,͙��K���c��-���h_Z���%L��E��?(�y�8r��i���y6ͱ�r�N�'w�g
�@$d㯉�lY\O�o^έ�);�����8#ƶy��ڟdM���P�������;��D6��J �'���1����fc�\@T�(ybt|�B�$�~c7m ��r���Y��c�!ZLd$��a�)6iC"|�a6�d�S<u	�� �y���6he��f�A&ހ�V/��Zg� ���S1��h$��hE5���PsS&�ʔ��x08�b�e�ڤ��mZm)A�&�A���9ُ�z6Pn��J�.^��{y��r�P4N�,���;�����0YD @�����]��n��'��DQS�㒠�@��k~&��/͒o��j�;Dk���s���SB�t��i�;��/�3o܊H*^��Dߖ�./����9�Ͷ�^¨ k0oǬ�p�jt�0����ݙT]B�$"�Ux��v��Q��`Pǁ���8��,�MR�>���{�6�Y½��F����� G��9�# Ho<�������SP�$��s��j\�[�,�Bo;?*H�1UE��!U� �1�L$��:����~�
4g�!c��h�b�+o�T���S%;%W� �8�0���*`�S��%�D��I�T=l0��Sp�s"��;���ӖkEk�o�Æ��C6y��pJ��F��w}�Hֆ��L�����]�����S��֪�2���
�N)�O���ߎO���qw��5�G8�tV�7�w=H��|O����>��v4vPK 5�N��8����b�+����U���)w� e��8�ܗ���С��Pp!4ݚ�%���A���Am������o�tm�0��RSݭD���PZ��J�c�w.�Fy��@J���B��9˴���	�#n��I�Q�w�҆R��[����u��i2D���w8[�Y��'�4n
�HK�Q�X�h��㩩3iFo�����W��BJx'��ӹ��)��0�$=۠+��S��">V+��_;��N,[(�5�"�D>5@B��Z�.��T����s��,��O�ly��k�9ڭOLS�=e�T���|�*�GϔD������^+oe�H(��T�b�
�~7��H��<{��e�/���F$�w��^�=s�W	��2��>��]�-�)�il�b�N�X	��1%�N{�\�T�<�r�_l�׃�WЛe�Y<���	�|�цJN�]-='��w�ArҞ��íϿ��l� ��{��L�$ÄJ����{A���ox���f*-8�,۷z6�\U��)�M�$�@rx{�ǉ(�^^�X!��X�hT6��Gz��s1�u�Vu\�V^�߯�d�n�к�'y�R,���k��*
��)��XK�y>���Pǎzy��4+�겹��%� �薉��C���$� /t[�����j+>A��$���cA�;Gl�rz!OS�2�P�
�S�##����[C�f,$�o���׾�Dk"g��C/4+Bqe��oo��A�_���h�����(�60��e#�n3臽��  mѪK�:����E����a���ż>�n��q$���]�'��ԫ���5����H�ϲ8�h���NBu ��RO��9�&dY�䕉!�E�l��B���6Bb!	B�ɤ�'��P�ۡ3��N}?�Es�"`͂ F$��=i(d�1�X�A�>:Ԍ�M�������R�~L�� ��E���J��7�U�z��r�i�,�����we�`=1e��	��������o�@�Ç� ����"���׋�_�E�µ���I��N:��Q�	������ݒ[����49��X��5�u\�9gM�F���ڂoW����큔�G�*.��_*F�@�q76���w�l��ݻp�-�(�NF\��_f��O�R�<Nf㏾��Ru���;�0�v[7��] ��eO�D��"�����v}��͟8�tH�L��&�L���YG��ݏ>�'�#F��*]��*d�9Ɛp�.5�K�j�Vwћ[��T���1�4)�Z��(��$m���̼�z�L���y���V��I��6�Ra��P��+�3 �Y�����f���A���Q��YD�z��v�̣�4o�W�'K��o�d�.��_�l��vFh0�/�WD��m9&Ю���,D}���3̝���~-^�I�U��WD�؉��+��������o�*KR�c�lV|tFpqW�\[F�mM%a��a�jU������,i���j2�7)�k✼�@���������b�P��z��ݳ������,�#[�R���̇��d���<�rk�:�4c@A��?!��Y�Rabe�1 5�A�ܷ�I�����+�	�J�����jl!�<��I�,�U�$6���� *�j�߀UP����P����q.��rh�<e�@(�2X&�i��GgV㍒�3@����Q�e�9[Üڶ�Duyܫ.ڡr�$��~^�g����Y���ǖ|�A�W���j����;���.o�Y��p���~��$E�/d�PN�q3�;��؊t#s�J_��������i�=W�㱍���Wl�M���B��>?}X��..ʞ��N�sk�;�j\��PG��]�_�_/��������,��h%x,@?�u$��am����,'\��:k���=�a@��EM�(�ܔK�sR7�=�^���߱ݷ@]�Ȍ={�Z�J!86�Ȼ��=0�!�=��ӏ��K�����V�*�7���ܰs�!`F?pO�������!ʑ�R�ZX|%��g�x$�`�����S��:"����	0^�;���)�*�B�Ճ�sR��t��<���βx�a�P���_��r�]�e�����d��q��c����,f�а�c$I�=�����=ې$��x�G����P�m?VJ�լ'mHH��fA�A�,h�|$~sz�1��h��1-;���'��$��*��\/� uX$G�¯������H�[������ׇ����u֮�I<�|���j[ao�����봕�|�*�Y���s�[�-	�L~i���sO8ў�{d.jg��VVG�/<��uh��"���]U^�[�)���?��v�_M��!���`!"Z��c7�p�.#BFrzal2M����3U��=������F;p��m��U�Ȏ��:䫗�FJUmD#�C�_��[�8��G�n��˹��2�[r���qg�lJ�U� ��i���o�'��ș����_;�??l�c��(*�<�|PO|�ԍ�sf���=���BW�~�}Y����h��x������iQE?�T*2DE������J��3C�~�����cS䝶ɬ���/��S%��ԗc�Md�_HkX1�-��`Ģ&����:zŝ����;�]�����>:������I�Ũ�~�zH#l�<�v0n0����l�o��1B�:����nǵ)��]���Ƶ��Rj�w����'�hҗXZޱ�u�J^�4�~o��bl�+��]�Ow\�7?�##���1�Z�A�]��5� kM��V��i(�˲:�`P�&HK�m�^уȪ}�L��;5􏠶��h���~�:��r�T��̘&o�x)���p�ϻ��s��_& ��:����$CSfc'������-V4�f���Z�#o�E��&#�{7o�(lr#�h������Ǥx&`V����a��7�J�b8H4�d�z���)���I�e��YLLGA2JK����P拺XHU}���N+�wPVC.�[̈k��2�L�c���
͡�m-5o*[����>>u<���ɩ���E��%?���|�On�z@�Kl5;A�M�d�ZA��e�i�Kl��o��uP�q����}z��(��b�%@z^"�g9v��dF��'�ĉW�0�2h2\R�I��R�=�L8�h���	&��H�_�;T��LF4۱�nU��>^�m#����tH�ɵ_\������7HL���Ȭ�����(-+��~q�^��hM~lȃchѩ���76�g�,*�R��e��ez�K���P^�t�¥Ɉ,���k��򝵐�*�y�*��I�����\m��w��X�*$E�w�#_[���1C���ae1��h �R�/1;�s�7��b7��"�/�V�ͯB�s����S�	v5t%�Md6���j%�nvZ�(LM�~%�Df��	К����B��:O�}��K:��;=�/��c�:.��T� �9sRn��5��O��-D�z'b+k���>pI����@�d֛4x-f-c��{Ǆ�U��e��L��b|�*�A��X��}@J�Y\�xf���&��l¾�Ѩ"U����_�pPQ��o���r�=MH�L��N�!Q��I(RW�s�f���`��j��;��� ���SW)��"�	,���*gʘUΥ��fíc��#|�G	�z��V$N����-\��9.��L*�3��Jo*��(���H�K"D_�{���k7��<7"9E��ti�D���ɃG.b���	y>����?vN��)9H�������F3u���k	�xLf4J^�p�~l��o�e�)�פȫ	}���|A�=�V4� �G�����ᡜZ?9&��2;������:�&��cd�mS�F ��%{2zC��ZF���f��Ū���j�ᢟ����)���.!��(A���@0��|�#[��ջ"��9G&!�u���9����R�ũ���x��+�m�x��~GA��R��R�L{��}�2���G��GZyj�������qf��S�����fAE'<�{�Pv��<ڦ���A���v����=�	�?���KXsaAM��8�;�@�+=U�٭��	x�QnӰT�j�{3^h�:��	�yܞ�+8mE�	�:�*�Z}O��%/aS.Nz�L1O�3�n��ܤ�j����;���~���P�vl��т��d ��ķ�z�9֫�z�i�{���9������;+"�pX�Č�͝�O��1�3����	C
��"p-N'v��<���O4)͟��8���x1o}���A#���qt���dMi4^#s���l;q�Zfy�s� l�@@)KL�$��#J����V&�q�ԂK�c�G��Bo~���Gԇ�2,<><��,��.�l�q�@.L��i�	�b!Jˇ��B�)Pc顋�qi@��޳�Ƭ�_�]���l^_^��i�CCN�6�[65ʬmWI<�6%Tq��ӮC�(�rJL�7k�å)����C�����BA����VV��L�x�o\xh�+҄b�!�-�n�xF>m�����/u��.�\�4Ͳ~��Hh�\/K.7+R!�V`ⳇ�i�_���m�<+`��rV�'2=��4�:QB'W����K��!���	f����a�f\8b�	L;�vSY�Gb&q�ՠ�"������X`m�1eF|Pϵփ��&e�~Z���l轁`9LI擋	���-��_ �o?�޿�<r�TYOܿ6��$Y��!��Ov�'�u�����@�>��b���J�$�"Ĵ���e��{VQ�&t��"*���;1��TD�V�U����!u�:�AiӸS�a��~�o[�e{�oJ/طc�O��
�x4�!͸��?:9��G\hD��J;��XLr���� j4x�Z̀���[{� ���=�%���"���ܖ3_8p ��7���E%��S�{��$/�+#�?XLk�f��T����0n�,%��,�s�U���.��Χl���d@2�C�t�ӥ��$��f�I�tn�T`3z�\�R񍟎�7��w�W�O�]KF����j~R��~��a׶ ���퀞��O���2q/SKltנ�$x��{a0r�S�7QuL��Ǳ�ЗbT2;�� ����s���=i���9I.�7����C�YW���*m�ʩ �k�I_���L����h@��i���u� ���t��o%z˂8�58��D�w#n �]x�
X3������N��v�7I��2rR��ǥ>�j�q�;s��8	����K0��j�)�t��S?�٬�K�
58"^������{G�k�X���9�����~��X��ƕJ��[����C�̏��FP�jY�ɇó0ҫ���O�n����;�{�;�S�Ͻ��5nG��׶�㺽º�(s��dq_ �&rM"o�9�/�o��.P���E�1���Eq�C�T.IC��n^�t�`C��h{p.�dYَ1~�do��
�7i��Jb_��`��Z�Ըm����lt�צ�.�-B)���Ud�^T�	��b�-7�32���1t����˭ȅcG��}�H�=������D8J܉�ֺ������XS&�Y��BɌt{�TV��,�F���f���8�+�O�+M����f�Dٯz.�p�N0JCκV�ݜF���un�V��n������zd!�8����N�\ײpÐC���|r�A�X���X���Uf��"�EJ�n�Z��7����Y��c@[��n��z ������t�L0��L�ڳ�}P�����݃$hZ�AvF���]���
�ġXG
3�@Σ�x]7����Z��6�ѕW(�����
���E�Y�n��N_�p��H��8ˏ�YotQ�� S���p��x������D�����m��fG{�%���^%����3[�	vIq�ob>� h����DU�i�����$��G��Ֆ�����}z�����7c��oQ͈z���)�ق����_*�v�(i|�ՠ����4Wqw��%Mei��懲7ޣ��
��u�xK��<�����j@!�<�����9Em����GgϹ����` �q�\ VC:�γ5t�N($���*�)D����4ߠ,J#�����kW�`U�k��dƽ�$v�$�b2�7!��jR���u9�����;#'���A�*��s��	�$��l���A!�I1�^y���k��t9�̙P�lI+���F�NQ%�X�x"�e�V��x���kh����KEw��,j��݇Wp�H6�Y��$E���e�Q=���l*6є��\��kJJve�t�����0j��V� !�r�������v����/��.a���c����|K��J>� ��3 �	9Y^1�����3j?��}��dU��M]c\�]I߂�܁�##D �l�_~q��@������Zc
5&��\�:����T����Ȫ "�ŝ��J���_L�^4)S���[��q�@�В��:��1Z|���V�v�A�oWd]��lS�MiԷ �[��L�B�:���Cب�v��O��ʕv�Fm��y-�c6��z���k�~��g�"d�����?pj<��N�:/!Ģ,oP@���� ��Wn5e��%H��D���
����=6�}��>X�<w8=XБ9��.��`�Ex�U�LA�����B�J{D�Ly�
�Hu'�r������A>#YP��4	���w(*�	»�&�,��,����Tg\�v��Ur�D���{�U����~����诰���XA�|,��;��ɞ�Yo5N���^�b���7N��4Z ���ᝋK>�\���y�lGg�K���۱
�:S]������F��q�	�T��(K	b��n(v�F�z>��ω%A;۫�#���?�2��M� 5e�wx�]_A�_c�ymF��T�C|��A���9N��4�L���Wn?�`�ߧG䙜R��h$�Te�~��P��.���	́�?�s��l��}��o�r��9�Q� =̺�<%�c�%�{��D�hiL_��C�:�b�6�V ���[_�����H��W��<"��\c�d+w�f���&Ɛ�[v��K����=�*��6K6&鳜��eӝ`��N*���2${�;���t���ſl���[���;��/�f��0��ޭ��F�g�y���wH�*��D�]�%c.�������ZO���0��ec^���Cն��L�*���O�1����S�v&9��y�n����d΅���Ipr,<���X��k)Ts6~"�'��fc�zk� ��,�wn�)���`
`���kR�/2���V	a�ʉܻ�.��$��_����`�r��UV!�YC}ɑ�P@��~V�7�Oq����i�I���|�)���-�f�ѻ8u��H���R�+�������&`�_{��H�&�4�����:Z��o�<�%�����<�'_��޷YL��=�Ve���t���ۿ���������B�_�B�A/�9�TTN`���J�/kYg�MRC
��P�6�Z��qW:�\�o�4�<�P�hm�ڤ��CT.��z1�]�ެ�l��R�7���>(��oD��1*�U�'h������_�������ꆄ�g����k}����֫n�꬟��t���㯾���TӠA -H�l���Fܽf�s������n�����SO+a~/傢GqBQX``�
���c	Q �����ao(Dp���|4Y��
�b�06��W����;��K`�h�-=W�_ ����=���x��q��2��'y�=�n�($����_��{ .����Q����t��ώε6A.����� ڴ�O�3�j{��'�{�K�����H<�49j?��	��O���'4D��R$�^0�E�X��7M�f��P���y�aJ�J疕H�8�
�����"_��%_O���sDQ�^�xz�Rc��jT�U��Zf��k�� �s�"�Y/!�R�[xԫ��&��T�����Phm5����X$�]h���+O��O �l~@!vq�W���L����7I��M֡`}L��i�o%:p�	�~M�cH�
�T~p�ў={����_HY�E��đYôt\slq��_��.��`X�b]&P��|>�n7d� �RD�����6se��3�D�]@ ڡ\�]S�,l|sD��$]�R�,INU�a�u+9�~������rQ�@2��� SC�*#]��o�k�U!l��4O�Qc�Kͦ���\֛}`��
s�a]>�<�.��Ђg,�9 �S{�ՙe$�p
ݐ2NXު�N�%�wnd��eHp_�Yy��0��e)�y���)�����oE��dox�!������`h���~�9����b���Ǘ�fi.?!�c��"j��o���	��j���=��1^!��z����I�G���A�74�a�.HVjI���N">X7�pS����-1z���?�jp �Ǜ��H�m5���D�y� ���������0�,��EwN��X����q|��0�W��������v��(��ں�-�%�BB@VD��H)\�g	�S�Y�T<O��2����O1���#2�Ѐ:�d��Om�}��8����<���	ޠ���hns��9�.s��ȶ���rG�X��Ӈc�	���͟\�ik���Uݶ]����fV���YCpC5�H���FS�k�U��f�^a�͐�D��d0�������4�T�cr�E�4I|�Ԇ��;���?���_���7�!�[��V�m3��/���ӥ���v���`�����*f�w�uL�h鯓������%n����T�W��-�wߚ'�@�Nt�1�]&uqtcU+�Fp�@sM�1��̹��f�IC2�r+�RǑ"�k�K���C0O��j$�%�D��~� W|d�j�wq	�ɪ{OR)�ݖ�4�������MX��&�f�;`���K׹�}���ލ����y�k�����cG
?A��bˏU���4�C���^��;��@âs)����׵O���G�
%�`M�Bl?%�׵�훛�y��?�����O⦠�����9Le��~�oJ��ңS*C�v
����˨ 
�{ޛ�Ĺk5���;��ޯ���dp��k��� tP�F/� 򯷳�}r���k)����/d���k��>���v��P��޵���9��wo�Q���u�%H�Q�Mh��T�U<<[��|���֕#m�9O��r
�*.e���?�1T^��.Ĉ�S~N}V8OC]�=������+�J��Y�P��/\�Pm ���s���c_ﴵ�h_*����t��Ue�_z���N|��F����iaCr�Y���A^��0
U�5A Y��j�#LJ��A����/d����[��i�,�����>�Jc:����[0󀴳����$���mQ������5^\%�G�Z�r��Q�)^���ޘ����E!�u�����Eyk%�VV�+4��y��a�>��b�HZA��asq�)�K��R�\�~�>�>XL�[�ߣ��r�̨��]�I��Ov��P��"��@9OJ:����d�H��Å&�$��h�$�JYК�->�ء�vň�����F���X�T�$�\�,'#��W7�y4fq���u�83O�a�,)�����=��^�˂�4����)����Id�fЏߨ�~���k�]X�|�Rb��C!zI�]�a�z.⚖a�0�CC�H�f��\\V�:vz�Y��:>���奀�r���Kiȃ���lFß.�K�3>�2�k��t���S�6���X�R�P��t���r�'��p�������T������]tP-�6P�h�1�7q�9�l�I�(����h:�o��1W�4�dmUX�k��������m��U�U�h�N/5i�����ϏZ	ieK֔��qΞ����T|��&�E#D�5�K�B� �������5J�ܨ�c(��s�����T���}9|r�tZMg���B�W��\۷T��n��u�޽q����U�]�T=� $�h�TL���D1I�7�̲��g�=��qN����;]*��,i%�~X���_�I�Yy98�.�FZE���c`%S(�T��Χ}0���_�Y�p�7f���r"&��珦٢Z�ꫭ��\�à�ҥ�1l~���d+W�p4B\�{P/�����Q�����(���3�̥A
�;[�{���EN<�/��?�jv����1`r�Ɯ��ŵ�F��Z���Z��/�MN��g0��y��jjO={��IcC��hWR9���G�H�ê�٨��:��b~�NJ�o���3X�����2�����x;W���cz�}��2_����ǧ+^R�q?K��HA���7 m�z/���BKY(E�@j�����:�[!U����W�]�i�Ov���$�th./e�d!B�����G!�Y��<[�\ݓ�FI;����#�l�N>{�Z�� �(O��֍X��||x����q-D��=�ӡl����!e8(��C
z���������LM��� fUV��XT���@�e�n�j��2f���*��6*�t��3�J����~a��̪�J�����y�XG$G�KI��y�1Ie�e�X/��8�ԊTtCF��n�^ݢ�����ln\�5�vC���cQ��X���*��Iud�ଌ����҆)��Y�>CJ���$#�{�~�hِ(2cP�r�Ғ�ѧ��n��B�nl���,� 9�.�@=p���/7��!��P�9ō���۰����n��c~S��9ֲy��re�m�*�O~��ƽ�,�S�YN=PN��J�
��ᩁ��b<�Jn�{���n�e�|hR�%^ږ���	GƇh����o�)��Ƴ��kk��& �l�(2�֬�UK���������?+EL��Ϙ6,�>��iR]��T*�����|XOL�3f{�Rpá�^5#Ww'�YQ$�L?� P?�r��5$^���7r���>�^~�3"x,����'[�o�X�$8ʝ;<�
z��~�`��W^��H����G9H`�j2U�j�z�o|Kl/���|L�5��K,��I���7��/���m"E���?�s�+���^:vrq���qϚ��W�I��� �K>��s��;�d�LZ�f3Ի�@�����g�zwYK�O# ���P{;�c��j(�[Z�
x�����$Gi����N�yAk���Ř��]Tю��]�"U�+Q�w*Yғ/����u1s�	� �����M�:���;�������Ko]�>��$�2ɡҗ}���^��ܱRt3�lRѤ2��.T)R}w��TjK۩g���z�g�B9��"�R�l=�s�%܈�ݥ�	����E�Og��>K��?<�U?}a�}Vɺ�������v�8��tu]J�5Htl�|�Ņ
5���Ga���jq�0OXY��Z�bo֝���gX@VzY�������؄Y$��N����z`�u[KH̀���'���� (���i�m�����]2ޖ&���*n���]�?9B�_����P;</�X�ٵ�t��M��
�Gs�D�LV�u|�$4��H?V�\M���3ۭ^y1;�^�h�"�K�Z�����<]�:C�� �_�_2��'pʦBO��3�7��a�����>	 �J{ft�'��8��h<G��(���� L���+�����n�>����vO�jE��
-�d�u�"G{�mLU��M�3�N���Ɠ���dj\�
���	-*�>��n�#<0*i�-�S�����M�� �P[�=?��(R��ೊ�!K۪����Хfg{$��b�,���j�	-�3�
˝0���4��4�����렯`ԾC!�$�u@�V�h ��e��y`S��*B �:���Qks�ށ��:bC���.T�L�ؿ_�Ȕ���l���/�)����s�7yf����6��}�Oe�3�zHs�(�@��N����%��/ѱ�po]'%�'w�g��ANf���{\�����"�CMM� t�ޮ<�hdE�Le׺�1VYE|�|/�z����>䤛{�I���W`f<	g����к^V#mJ���;��]?|#����tY6�wF�ǚ��ċ�>غ��.ʸg9�h�?�u��z��/k���w|�~ڠ�dYi(���Z5��tg�57�H+�B��j�G����S��q�HSCm���Rx�(W���R})��{���J�nyV����=�@x��0�d����x�`��ɞn�v�G�O�I�?� X�w������Ɣz�G�/:$�V�`��Ϗ��`x��FN1�Q��U�2�DGb��5��0��|�9�(T%0���:�MC��V:<�g�1�2�l����}�<�`���a"��/�ζ����!<F��f,k޷�K�\:�cJ��T��YX����F�.���9l��)�Bm�
�q��tD��FLg%+^Rp��'p��3�4Ypf�&P���)��0>�����K�z�i�$H�h{R�o�aH;�cH�WLJA��+���i�H, S)��g��#���|j�Hx��g�H(.�+Ov��
�&^}x-"��kٍ~���\�\Ec��0���=���1E�>$&�
������5�|~� -��/*Cp*h��(�^:� �>,Bmٳ/���}:ʾ�*�J|�Q��uQ��ɵ�	p��,0�违|Q�i_��`X���4�	1��Iy����h�u��,L2����_T}>,q߆[�vř��~�և��cʝ�(�!n�Z�~��l1{��"��p�q���*���t�I��}Q�u��K̜������Q�{�"0�ZqS{\�g����PןYe�OeӁ�wM������=��z�V�9�����MX_��ί�@�Z�;�\; �Cߞ��ը�=�U�vZ�����q��{�r� ��n9U]�t�����VA�@�t͉� �Oԣ]�f	�e��2�ߕ5�@O��8�V�t;�O��/=�
���s;�����x'�3]F���u���8=�`��n��r�//��b�~��Z	�jt;PS�u8���&K�4�ռ;�r�����>���߫�Y�sf���{3;���qc�p_�*�es�����*�	���?�rzn$$��h,���fo̍	�8�㏚��F�a̶�6���Z�Q��|���v��]Pzd탡�oCY��P��c��>�%�����ۧ�&@�#�w�D�0f>��{�.0*�n�<�~f�0?i%N�n�JS{�sF:���2������!*�xKY�=�.����?pⳞ�U�J�*~j���x`A3doWv����#� m��%�$�#<���� �`qa�cM'��Y����s�Z�/&sU��)5�=%�M8$�]�I�D����ő^�lN��f���+r�\�v�̭�ZN
k�U-���Y���a�ĵ�j��
l��t�V�;��?���kiY����"�.�?�M�}�k�b�b�1/�唔��O}_?��ķ{���9�uq��n�1M/�0��L�ᓮȑ+6��}��� եLsq��$Y�e���<;�����2�v>٠���xZ L��ʸ�BҜq� �J���9�7�hr]�7q�O�n��j�W����� ��@��1ӿ��c;�ֶ�m,�a��TcyM�t��{E�]�@Y_k2n�&���n�����zQiP�ݾ���;�T���x&��/��031��		��F�.���c2�z�xY�K�(C��1ƪ܄{P/hNE��
H���$V�C`���9y�����߷��QڟJ\�斔(��s�@�B��J�Dn<��,�8BW��ejv ��xa����et���!�׾Ű!+E���;�u��\4�_��v�s���^ڹ����m�sWR������ގ'�pY���H�5����"����Ǆ�n����%�G.��X�,��{����I�ԅ�W�
m�h��sͤ�]��o���� =����&�Y�X1Ò��8�L�ǋ��3�{�BqQu�ЃP7U��?�m&������š��Y�� �Ck����n4VH�ǚ�/���H|�"-ڇ9P�ׂ;�962R̔��W���j!�تQ�er����l��ȱDU��m��F��1k�B�}1�L����3�LK�� �_7_�_Xp^]_��Q�$����z����(VC� ���_6�:�-��sv��T���Lb;��;L=�KD�:��2�o+K�B�5h�c�\�U�r{�&�>4����@�W�ú���~@�v�Y~eǇ�K���^d�F����_��SU�Z,<)�C��D	^bvjmu�1�x&V�؏�1�l�C̹��i���ʋA��[��a��,$
SH�E��e���N����r4V�!���Ub���(�d���è��
�a[����N�n�PO#�tKJ�v�H����lH� ���{D�������#�E�&՘� 
?�s�O._����d�i��GeL͠E�/�+����3�PF8Џ��T���#��|fťgX�jѫ��g��$�t�Bgz?��^��}�{GN	-�$3s�E���a6CQ唼0��1x��B�ud��,��Zh5۸Hv���X��
��0k��SD'�&���윪����d.L�*�X7z�Ip����cj|��T@�%r i;P-�m��g���iyAX���)�t�.�ULP�i�@��x��R���=#��B���t`Pgd5S.����`l�����r��*IQ��+./�ox��(����hF��aQ+^���N_����m�Pǳ��|�,�
�^1��.����gt�X�6V����0�b/H�֛��L1~�| �_h��9�rN%�b��_�_��q!�,�4|��UJo���0�ӡ�IAD<�D�U�\��t�Z:	�"�(��@��&�a��JT[Nm���V����e�������>|��C�ɆZ-� ����Ի�ݼ�V�b!%a�\�:��v.𱸄ۚ;4I�3Z�g��3$b#����p�G��'l�Z�����H?��k*C_#ʶ�5�g��]��cq�O���j�%��e}�3�X�C1�fb�d�i:)r}���N;�K3~,��l��Pǭ��b���/D���L
�_1�6��H�O�?�f��С��:���C�H��w�Z��W죝v�lN�PL 4�r@���k�j� 7��C\A�>���aQTN����!��a�nGN,�)	�%�X+�Fs���bh]��x�������x/���xP ��E<���&mfl$��d�ofl�k(����B}O\����H�����PUM��gTC�PxGXRN�q����W���`rfI����L��p�����y�xx�D%oeCS��M�w�&<Hn��wFIM��U�T�~��y�Vh]n�4�H���=y����o̷>U��Dw�����l��V�v@��a�����=���Ȯ���#.,H�:�S�G���3m��X|��lԤ��u)�A�'J�;���f���n���@��'u�c~% �oE�q���[,�N=P����8���<K��֨6̐��ڪ���L�NI�'}{�O�j��{4��@p�E�-��MA��.f��[T�<�=?a���dc.O��d�"-�'�Nˑ>?�t�ZL�u]��2�V�h�&wۛ2�zx^�z�m �.��l�5�V�f|`�U��#�	y��+J�<�T8/�o4[�E�d��y�_�B�Z�����w.�����^��9� ����{J)'3h���j6y�.@[Ʀ��V��z�I>�����P�+�s{�v���'��Rc���ݪv}R��8lM	o��9�{"m�Sꉶ�vƙ���M$G����*����9兕xX�"^B?o�B%��M�#OWm����%�����Q��ŶBn]3����#�%gX��s%�1^��v69�SkU�0�J�/�Z���Y���N��i6fSZ�4'vN�Bj��vf'���PL��a���+E^�SCM�.��R6^��x_�ٮ#?���������S�'ʲ(G˲�B�q,�Y��Og� @��ɵԑ����5C3��b��/�E�Ԑ~�O$���NA���aJ�;�)nR��~eH��קZ���OW�@Nn�	���̣��
v_<ݣ���%6�)u�7�R*��3�fLƑz��<�6�t���X�1�����vVڬ�q �yZx;ry�[r��`,E3��
���/j�P�����l���<�Y n���C��UY(�$��fQs�QzmѢ]�I�>�������!�G�+�#2n���;�<`2Y��b+�����Hs6Ts�r1�ڑ��{��`z���zz����x`��9w{Wh9�|���uQD2�jG���VN��L����U]����Rh���?��JZD`Q�:��%|�B^azs���j��H�6�]��ܠ��x
�qr�3>va�+���]�8? @��<|�M�ݧH1��:_j	G�>��k�$��?2��SN)�lsQ���-�NУ�<�s	z�q���Q�ym�Z�����H��J!�&(~Q)ѫ����o�A�H�g�n�v�&}�o�띹 �%��mI�����Ru$	*z[�
oKE.�D0ծ�Z��,�~;�����g�ƙ�����F�q�\��C�%\k�5F�[ǹz93b�B@S�3�h��}.y���*Ga�5�~�FF��؝5��`�Q���2ۼ��U���2�SR�>E=>](3�P�k���
��y->���8+u�	�B��JO�@���u��ƺ&r��|�Yl'����o�`&0�D������&��0vL��e�