��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�۫k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��5K�z��!��[��S}Σ{$Gx^����c��Ʊ�U�I��^��m ���"�7���4N�*"����=j�� Ơ��� 4�4�?k?��칹E�u�ѓ�K8����>�E�VN`�j\ �W��K����<t��M �L��«$e�r�8�����gT������,�Rr��׭��)O����EI���>��uG�db���4E��E�c�����HZL��DMo�vQ�A|]S0��y�z��*-���	mVgyj��c��l�`ʞ���)�/�*\�k魉��NbR[=�jd���/���g���=��|�|e,&n�v>�*��o^ϸ�p2�|���4L2YPUm��Ax�jS6eC��?'/��hN������	<��,rǱf(Y�����0c��s Gc�k-��a(��~���`:?XL5bF�T�X�Vm��F��nR	���}1u��;���ر$��ޠYcj��g�$	\�d�������=��wh��o�Q�d���-e��P�1Տ>�����Z'փS�;Ó3��%�L��Z|��T�w��?r)��� ���ؼ�����%@�L�x�d�Z!�n��?S�:fVE�8�a���-t`��'@�hF@(p��+
��R��%ֳ���w�,4����ꀆ�L~<)���v�\�����j&��syų����K�� Չ���RQV�U��I�e�d��G�D�nIRJI�P�U����}�$]л���H�0��h7���,��ᰭ��>뫫���kEF͞�إ� ��ǂIF���66H�m����&��RNSF��fLe� ���cP�i�^�4&���K�ϱ7ߡ㼀��sK��56��9�!��'��/����L+v�xw�����X�<w���gytI�`f�6�pr�xy��=���Xf&�����%��1�N��ѿh�8��幽��ѯσbń�:c�2m�hm����I}�!#_)B�%��^�H0����5���$J�i�ߝA ��^����G�7��Rx!��ztj�w,�	Ƙ_R������y���݈�"vǯ�&ע�[ͽʠ�DFY��z���St���D�B'�*˫�;���V�-�d_����|ˇ���	@K�y�m�Ut׬G�|2�*l����+sTĩy*(C��X�y�8L�oň�,8�.gnh�H^�e
���Z�:<���p�R�y�<�9��#�d�>�gd�*��,�E�	���C�xۆ��Q�Q��yT�滿�I���Mb~x��Mt_�GF�ɶ}�,,	C1���n.���+��<�Z"��z�n��m��zޞ)e�O�@G +�����x�<�o.Q:�kQ!������GQ�1Ɂ�v�y�j�ܶ�4nq�Oɐx�ϘtD�ϛ�zq�B�����q�l���pLM±�:Z��z�d�P�S��w�]��� P1�e_j��W�����g��r�ۋv���e� ?)�� Pt�-��R'