��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,��.��̡�+P�FuX��d-��N��$%�I߽7>wN����u�]��j��ܹ�Ucל�|�=í[~��k�5�P�ؐ��T�5�����#�p"&�l�z�Fr&b6��,���Fԟx�ɅT2n�x��p����Xh	H���9�Ҿ�z�1�� dT�h6��[I�����B�?Oq�_2�9Ӑ@�p���G:26�[�6T%,&'�#JeR�+񸊎2�Դ��E�Jc�������5N�{�����Jz����+�:��G˦�<�_�	�'��k�Ov-��5l��|~+��,�Z��r(?�! WD_����J���K���םcE4��%2���qb�B^���p�G�A�tR+�)«��jF��s������F��[X����e�Ԁ2�F1C0q,ΣTDt�P�!lȏ���$k�4	�O�F��/"�k�F���@ͤ����mj]���A��'26���y�Y���.�NE�L�*$��ǚ!(+U�=�5��8s�H��9�y/M��>�W~0�����bW�L�hA-�������a(�����ya�[�|�%I�%&��S��]�q��ͫ��H�JZ��v�8�K�cdV�.��\	�`�9���Y����ìA�ܮ�$��a�����0�U��N�1�N�QĮh[�<.�=�=��M�܏_���aJA���F;��Źє����q���j�
�3m,M_o���@Er���k.$�hP��ɝ z(�O��
Gc��y5۲&�j�6��������F�	���T�lNu�h�@��Un�����z6;�[2(N��j�V#v�� rܦֆq+�PI��n-����S��	k��ʞ�<�F�YN��S�I�M�i��h��yq$��I{,y `�����i�LC�:��׹�y/ԋ��@gktq-�:�
��r���s<�6������>�|��Ycw�f �������,�Į��YXR@	r�&w�Ԕ�� vdݕ���}��m��p�`17>���$���ul���Bb��!��i����Sp�D�ڡ_�����*����Z�@y,-rB6)vY���$pB~���/�B
��C�ʗ���\�_�l`��!��4�H�T?�*�A��zBsm���L@��X|vD��K���3��P��b+�b!l#��]v5��{�*/s�׷��� pI�Xl1h]��'�NȂ6n�����sg)�gS�ts�I�.�|R�0��� XVǹT"o�)F�t�('�{p����ё�¨&�\Sٻ�OF���/Z'��!���p��L�o,_n��#���^���}���5��E��ЧFI��P�p�H�G���0�����>�iG�P6p|��S�'���t ~�8B3E�L���G-cy/?��?([��=���(7��^<%܇�����s����t�J�:�y��l�*_����4
�1]z�yZ�M�w�=��7��E`m*���Rų��;=R78�J&W��2x�)~�����4�}fT�/�\���UdJ}_0���@�n�@俟�����I�M��4}%�C����gmؗ%V����%�93�I��IϭՆ+�����',i��JP�7��v�sL�Q	/�l����՛��Aziᡸ�#i�QFMe��ӽ�pܼ�������Q=L��z�����]!��˲��^����ț�'#��Y����vZd�"����#9E��`�7���o?��&�Q9��b����L��E�B��{9�Momx��ݲ
n�[� �y�Cg��[��7e���{p�B��K#��c���L�֋�����(B���9C6�G�D}B<X��Bz���ȗ��ld��!��|i���o@�*���Fv~(�>錍��bZ���h��=$���f��"�����[�~�1A�R�R/=Kl;$g��os��å}�K�/G��Q7��d�y{|�c�*ۑH���1�RT��#K,�j��[����V�1�=| �c�#R#Ws��AjE&�=$"��d��D$Φ�C���~��y�=�_�P<s�)9�D]!.Xل���v<7]���ʼ��v����VX�r�#����76/�U����C����tm�ڄ/�D4�^���7��KS�D6ao��]�J�*aW"�2�jÞY9��G@lE�ç�~T���+�A�s�C��-,�K��]>Y�p!���-H9�]�$�Yk�u���x��/���X�]���d�{̎JB��N�Gss�`�v������O
���N=|)��+`6���P@��H���ʊ������c`���E^L����t9/'^e��H¬�T��pb#�t[��y�Dc��@5��|�<���*�jT�Ա3h�SA���t�K�z��Kt��Q7�L�d�Ȫ���;��%\��Ae����F��˼B���&���s����rIp=��!$Wp��M^�g7T�����9��-�E�E���Y�B�^��ְu�J�Z �m�[og,}&�f����i��
��7(�