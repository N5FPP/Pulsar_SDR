��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VYab~'	G�S���n�?�zBnJ�g��|�4@���L6�¾��������S�df��oST��N�i��%@�Uv �+�p�)ҧML�+����d�}��xd�Ua�y��%,?���b�τ��0Dl�_�x�Zjn�T�`���7�B$G��T����<ŉ4\�4M)�D��Eb��nt�Nӏ`SH�1�q��L�,!����{��K�OLu�r�]M�kpmض=f8���֍c�a�:�pT����܋��WS%�+J�!��݄t��$O~�[SOx����c�#TP���SL��[(����jy�{2��(���t٪uر�mȾڨ���{4��E��K�#�~�T����]h���������� J��ڭE��c�}8��V��#7�	'\Sn���/���=4��R2o�Byk�#��uNE8�I��SEtl����gn����9�ä����V�n���?��].��'���"|��|�j�_n���dX�X�O<RO�gw8)��5/��P("�#=�Tg�-��N�kf�����j�L^Vn�g���U
��J����&.FP0o\�t5+)H����,3�������x��R�o���m� ��\h�X;�+3�O�b��N��X�$zOO;��\X�{���|c��8�� �4��9�����'/΅6������AE���\i���d;l|���ڿ��\`oQ�����9!#M�3{i`vR�!q��@�q-{�2�47�6^�e����������q���
\S���\�?ޘ���]�$����܋F���ispSN�r6�Z;6~��{�:Ѽ��0�����b�Zx3G	��5��((
�}�.���GK�#l+�d~X��"�|f�rC�J"z���w[o�&9���t<�:��o�N�)0R[�����{//z��_a,��x�����Z!3�#U������,]��N<l7�@�-L?�X��/H�8 ή��OΠV�c������`e�,'C������A0oR6CJ����/|9gosނd,e���m��o��L���S"���Z��Gʆ�W�QV9Z��W�i(��F��\�8�w�5�hP�=h�>�c�V�U�^"/�MUB�ʟ�h\ߥ�����z٫������@����J4#�u�����+��:�QB���l�yH�9婻+*�����N.tZ��o�+	��'���z��l�a)=Z��ު����,Ӓu�[l#y�ۗc�����G�A3�G[N��� �p⟌G\6ۄ�0��^(Xj�}Q�߁=W�n������[aʮ�T��f�,�2M��f�z�+r"9Q}�p��Z�TfT��T#�}���~)w�d+��`�a�n �l�:�S���8�Yp�Z&Vk�'z����g�Y��B!�w�h��%�i{b� i|(6,������v��6! �b���#��ɡ�V?�Q��Հ�.� ㆾ͒�,% g0I�'_�̅{��%w=D`ڇz��z��qiBZp7n�hG�+��T��UQ�������]�.��w�f�/��F��*��O�8c����6�<X@�	�k>!=���E}r��d���ED	��N��F��(�^/>7�<h����(W�O�T��1��9+�b��ȍ�ҁ�yͣ0N�8��:.9i����]���XH�n)
l���K<-�[��4�7m�Uܘ�m.�?^9��A�r}a�!�a����f�zq��������Cb(L���`0��\a\�����������H/�eZ�NP��=�r�]#3B� ����oѨ�u�Оc�Y�ޛ���Q$fM]���h��^�j�#��w�� s��g�I��R��w��f����ʍ���Qm��,�9�}��?D=��c��z��[:���wϬ�����A
3z��p�,=�G�za:��D��V�GgR�l��Lސ��+9�J�k�|�jKk�ς������~���T���o��'t�E�U���.�apE)g<�0_��nO}!S��H���E���۱ϿT��Cv�R������f�:�<�Zt���|�Mdv�J Q����Qr��;�dP���7���E�G�CJ,,U�3��=�I�_�Ge�_���]M���-jr���T�w��뽑�>G]�X��j�`QSk��Ʌb5c��94�գ�V�`���P��*���g�`���
���;x.�У�h��]h���.���/@��\B����[����C@ے�>}���(ظ��]���k�e�q��D��w�z�e�6'�i���kGY��Ȼ�����E	�8Je�,�*����Ψ����8��)����>�xS�zf�aWo���X���
�ITٗ�-^��G�ٔ/�n���sQ5��0��.�R�S�i���MaC�3��ZJYtb�a�uVM�׎�0�.��,n')ܬ��V.�#�#���eTh�9M����e��sld�M̘4�l�v��A��,�S������U��.E���Y���S��L�Mt�c�.�%nz�xHGtr�`���� ��������8��3��H��.<�f�9w�_�������,v��	�P~I��s��z�i׋���kN�F��i��E��T�A�l�i��+�
i��q�*T�~A=�#�|��MU?�v�,�oI:o�5[*�ʊ{�h~��S���߹����C�I�+hK�&ɞp�=ۢ#i��^��IsM[�zD/t���j#њ�<K�y�%������W3�ڻ�L��ҍ���%�v�V��$e����K2�J�}A���pV�Pۮ���9��[�;��h^𚃃(����	�G!D)�H��7��%����qχ+��N�H�Ԡ�pt$z������L�@6� 2iGn�1��1V�mt�Jə��C�6%++��,�wcYG�+�~e����gfG�@���{[a�&��yi����ͺ��\�+���:^�?�2ʈ�jZi���׃��ˑF�Zvu\�JK�Xځ��b/�o|#O�DkDұs1>ڷ&�'og���H�cC%�
B���g��q�J�ɼ1������
fT�Jh��G}�Gil\��p$�������ĵ�zdk#��"�|2���5�N�:���)���l
]�u�͗@�x�1؋f ;v�q�Tm\�`����{aF|��mիo\�+�ůԕ��E���Pt����[�����G<����ǔ�Pv��cJ+_?O2�C-��V����?X�u�>b�c6��v"k?����w���J�v�ޏ`گa�!RqƤ?/�����&��%�ȯC'��B�_0��m��o�хD�Sz���� �HI�A��&6`����n�<�e�E3JtUĪ��S1?�Q�{>4�7����Na&-�/:�#���e�3��H��Ny"����y�Y�]����̘O��*�[,��)"tM�%�Ed�����VN����o�q˟�w��!
9����z'D'O�PqX$�w[6'L���bo_h�Y�ܜ8P�պ��'��h��}�cu�$.�]�&��S��g������,2�<��z!߯8뤝d1N����ܺW��B��^A�[z� ���=^��R����dh�D��@njR�E5�Gc�Fl>8ڂN&�'J���QV�.;<��5Ӱ�J�sϪ}CY������k�?F*C���l_�QY0�Q��0���A���<�ޤ��h�F��y��,"O��5�a��S�W$sx{�; [�L�Ν�vE�LӤ�~����<0��"	s��=��7����ۀxHq5������Q�(���&�?����.酀�%�m��7��m��&�0�yh��4QQ���Х1��w�ы�</���c���uX��֖����jRO�m��oi��ӹ�LB������H惢��q)xg:>1����Sj�O{:D[ -��e!O�Zl��jP���6��w���h,ww��3k	R�����x�f*狞�Ϋ^����+�y�^9plw��*�.�(JqcO�%Z�u�Zz�i�l<��;H�KG(h�Cv"����sh�I�-nŻ˭�rw"��9��|���x�28�Cb�m�8�aPˇOJ@}km2�W�,x�;a���P�Ә��
j�(!a>>�ـ���`����>q����%�aeܜ4���!~�J�A�OY�[�I�R��(fǸ0�7�h����U�8R�<�H�@㦄rJ�)�v��):��7vO?�A�waG�r�"��0��8s^0pë������h�A8_h �r	�f�V- >�L���N�1<A�������Y��aA����"��y�`�X0ɺHM������f�\'����!�csh'a�Ř���\o��h.
S~�,]W�*�6����=Dc�B�B��8T��N�G�����F݆��uEugB�����{")���,ދӭ���Z�|��͑~�ژdv�6�x�oc.)H�FV&�?γ._�mC�ے#����ǃ�N�����ˉY��FF ��xe`��4����I[%9�Y��쮏HG���+E�V�C�ГK�d :J)��ͫ#�����8k;��5�Y��&5N�H�P��]�g���TԚ�x�6a����1x����of�3&xF�?�6����G��б�>�b�ЭZ��ڑ_˽��K�(�-���l���Uz]=���Z��f�|����#��+��\U3O2R<E�uP�Owz�xye���{vC}�L�L����Ǻ����"#���C�����|�%%��ә�M�JQ�d����l��T�lj�*�ZJ��(7��ޱT`�+&ުC{$�"�7�^��[�d�#Q��{Z�k�b�~
�|�HGQ}����r���)x.��eq8��_��)\���̀�22u�Y,�c�71��R%nYC<�����<"��q9�1'�h�����j�dի'�F���!o�ь_>.Qm7�\� �bA�2#���aK�>�e)��آ˱�~9�Pʝ=ȶ[��OC%<�����H���UQ%��ޗ������]�/�jV�:ft��êO|�S���]�CS��9����������D�����n㥁��9�?j{>K�lݝ��L�j�\�P�5q/�#|$��1>��ٻ�:>��0a�4)8��&8 m�W�w����
Y�2i�P��z�&WikN�T��풔�f�Z˷k�b�c������yc��"�ִ�7_�N$w���E�
C��ɫ[*@�n����|$�3�8-�X�5F����6ʯ��2���|�p;pP)�kY[�o�}���j��=U��"���J��j��.��o*�4���_?��K͌�X�K�)`�d^��-=k	�jB���!K̦]Ұ}�
\�F5�_�e�!dMm���Q@ʙ^�T2�~�q�-�<���bs�X��ڻ�Ћ���qƢ�ǡ{�0ôy��xtB�e�!G�������^D�p+��zZ�\����a���&KԤ��8=��&V8 3��t�6?��T�Z@�	�������
?�($�nP%�6Y)5��|�&@������ki���nP���=H����ncB��Z%�J<���<�W�YC����}����ٶP��D��hlG0�҅��I��p_-�4텶�R���}Sr�1E�|Jň	�I$V��D">y|���DN?�ce����n)l�E[u+ɹb�[�w��u��ԕ�����5�'��:AS�~���S�U��'�b68�����ʄn��\tbyE V"a	�׎��&��?\K�g�w��	�P�.���<i��m�I޲ȕ�T6sos]g1���J��!0�����5��e�'�ng�drʭo�oZ�b8����_�	TN�C��W�$��Ԛ7tKJ����p�-�	���8忝�Cr�tw$Uo ]�1Fj!���M�&�'�K�9d��]��w�U�e)���R�IY7 u��i_���tb��K�iE}]�g=CL��(�A#Sb]��w.p@厌O"$�_ m�t��RK� ��g�ˎT��^��y�Z��shN3�!J��yt�-�O� @���[ρ�Rf��p>��o��8���0�}n���\=��+�Td���`�"s�����O,���q�����Y��b2�3��W��6Ͻz�9��\��perQ����Bҥmc{+Ç��b��g���n�23g���`*C�V�����`�f[�b��/�I�f�5�*�d�����7����=-��1����5�}+'뎯������f��BN�U:�����zH��P�I��^YT�)��@�#YMA?�W����/�WT�M�x�;yC������U�8�E � ����e`��n������/3�B�W����4�Zc��Hw�v�?��S�g�VɈ5'F³AY_b������>T�����L%���b��5L�d�EC9*{K]B��V暱V<O�M���r���O���_�Z�)y�=x"�"�/�G���d �j��g7��N�?��/��2��g�(hnh$�I��}���;;\�Q�?A%r9u�_F{v��@J�*��gd~���5�������Ӳ��&��`)^h��_�3��df!w$`��u��������ܡ��%�1$R`����g�8���R�z6�h�b=���o���o;�Md/��W�wK��
@]�X/W#��J��/ÑH�	��cfH7C�`�A����A�D���d�}�lF�F�#*�TD�Fu4�ۃ�5ڷ�	-?�xbxS����9[�nxEb���jY���f�|�4��͑�w��p��G��r���H�l��~�K�~9-r%V�]i�Oc�޽fΤDȚӞ5�멌�p��f}�Yqv#Ϫ)J�:��q��{��Lb�8�O�U!�F���M9��q(I'yR��ͦc�{�+��l傐�.Ff&�r�m+��@`?(2�Y�:���Q+Á�%���H%ّ)�M+&��0�vg����d�b��"����N���C���}Nf.o<��t�Sƛ�Ts:�Y���Ų�6%���s�I8��
?z)P
��h��)�Ώ�-�{��T��!`�sZ3�p���d���ӥ���ҫ2�(�m�!9��y=�2촏�U���/�۱=;���Y�Ca���X��6��%�Ty�Y=��o��AH"�w+��Ps\��u���y{����	C+�/Z���\�����$���c�O����s���O�OG]���������D+ΟE)��T����M�T��h�E��� #r~x���K�[�R&*���������r���8��Y�q���2�6���GQ>�7���2j˹~=����gEr��~��!��E�>�@�fv����nz߹&���h~��iI��<�����@���w` �Mu����X��EWk<��F��i\�Y�Tow2���@$dK���_��z���5N�^��^�Fh�1������▍7���_��b�����8~��xKӆBH�'ȴq����e�E����O�9c��L���j��?�P K�bN�����<Dִc�7f<#�ɐ%��T)�s���&�A?���zv{�"Kl�7r��4�t����|��ղMB��U��ݔ��Sw��c�{v0Vx��1���n8Z�Hl"�A �P�d�#mJ{��x|2�[�N<��4`NJ���1ҙ.�s��c{��h�5��x��z���LDD�y˲�T}�����ۨ�R� R;�X�<���SQ�R�����*�}�d���V��_�x�ޭ@����t1
��h,��Ƽ�a�?O]|��;ﳂ-k�|������G��+�xr�1�}->tϱ�Mg�v�:�囦����zj���A�Iv�!@ ���V�;Sӷ!(^@�8�	2���iKȰ鹨ɴ��~�blJ���F�!.��vn
"=Թ���3�Iu*9ag�S����2�ɨ7���x�����L�6<��z�h����L��"��F��*jLy���+�|�@Z{Y����[,������Q�L�TcO� ?=��$����C����=X:z�z����Gx皬��S[nBE�0JBg\M�՘��R��짌ѳ?d��BT������u�Y2B�wE.�Zw�0h���d&�Gʂd"ݰ_	@ٝ`��5}E�zT��4����i���J�z��/�B8�鷷#���)O`�ӛ���޲�0�����H6�`��.�}�H��4i@*�]��+B���=ɯ�Y~m��ͪ ST���XMf�_����7�κ8F�CpO�5�3�7�|�,2�<"�o�5h��⢖v�y���wH����D����L�BDK8ᠹp�KU��S<����n�4�����W�[��e7R�E�,=ly-��`�$G;����1?�7Ķ�_�!`�PQL+h��ΉO�!���Uv�P
�6��SP���k`X`L��2��n}��cS�~ڎjmWd#�t��YT: �*��.0�b:h^7֓���0���7�}
�z�;�f�OMе��v���Z��g��d��|K.Ows8�e�C�E�d?�w�S�?M2����#�>Lx���(e��>��!�cJ�o(@�,���:�sF�B�L��u-�]�~$�?���"wLiw�<���B�]��_�C�2�"��a, �ګ��5�_������p��锵F0����_j`�$G�2�{n�z��6m<LuW�/��_�`��������vBX'#	�	��vxl#��Z&ºC��o���Z� ���V���@�k�_	H���u@լj�ϸ�Z����T�
��z?�Ɯ@�D]��.UQ�3#���n�ls�
��B>()��R��� 8Vϔ��ڂ1��jt�wPؙ�@ȥ������~��-a�8k�t�r�k�����U:�����F�Y�hv�FHH�m��m��t��h�K�DƼ�D7���W<�S��T�����)U�`IE �����#�>X��TE$����b�Y�4mC���TD�V��?�t�"e\5���*�~j���Pw������NҜ��%�\���^���� \$a1Q�6 u=۹����s��,:Kf�[��j/��� ���eOMN?7o�f�)�~,#��w3��ٕ�{�k�k�{�,����7���c��Cbؐ�fNwɶ��ʉ%N����V��m�ze�7��$�%�F�Nֵߢ�K�c�Qx�콲�C��7X��6�)	�!�z3�u�g+�0/1
8T�y�w)]�l�����q�׆~ۑ�00?�ǁ��t2�K
dY�l ��f׵�� *ߓ�nmYκj#o/�%0��'5���k�[���q�_Ҽ*����Py�9��i`i����h����G~�K���|�� �:&9��*���#4=I(��-�g�O����u5���%����%%��[z�N9c�x� �Q/�`��Tg�d$&'ja.~][���'D~��O5�x���<�u�����'m������k�K����O�R\��K�]i=^���I��3)�G�<�_=��ߓ������F��/���\O�� *�*k�@aB��}3�(̭j�v(*���Ҳm���\+�?�U�ȳ�u;g���y�cE=�\D?$*{JG-�D{��NW�4��â�U!ۀ,8R$�xyNOj�C�+ƭ_�lj0i�Q�)O3�a�Z�c�)�;�7?�;��n��]}i���G����)�S����(9�881}���q����6�=��0�O��dT���ע��1�B�¨0]�?���%E�#q��p���1m�q�x���?i�f���C|
.�'�ئbܱ�QF�;��A�܍`wh.�S�;��$aN���<z>Ͽ�cX
XyN�M�z���J��X�'m���TԆA \���'&��vߕ��?n�!���d-㳱��	"!��T0%+�W���)I~m0��=�> &'H�a�p$��
�j0VeH���}�~rPX���>��^�-��7�����b�=��6j8��rp��Z�iI�06<̚ 0kiDz�Q%���D��uXW�W�`k!�5�
��w;ͯy���'9�>T5QjV�R�k����K��__g�����r���8����uo�#�3�˻��Ml/��װ��wd�k~M���	��,�.��h������e�`؃e 9�V�u�A���D���G4g� 7PΫ�����0琪ҵeїU]�/~)�Z�����,��*��Ut�$?��a�Zd��>0~]�.�{�N���]�����@֖�c���ۅ���b8Xc�[Tvh��}���H�?�y)�*D����Uƅ`֊(��CP'��WۻsBPp���2��$n�iڡ�b�*��L��#�+[�~�>9�w3�l�^	s⼲��|��n�V���6���ή�������w�i��t��խx����ME r��Pb�����zZ.ܠu�mY��˵�L��CH�7��^+~��˨��V����גּ'&��MN�	F��K �;$Q#��%���b������V�a�+��]L��=��Xʶd_�3#�F�8f%Rw���P��Z�0p�rsx�=�ퟯ�����:��N�[�i4�+W�>�Q\D~�Ä��Q$�l�[�>�=Qr�YޙJ�%��U��_ѯ�E�/�_D�A�e��� ��B��Y���=#���(���bo�8�3@	y�\��v^.5�����eB��aCB`�
�۬�q�j�7���_(d'��!4Z��ݱ3����<��p�J-��J����,g!�����ٰ9�ܥȸDG�5� ���W@��`�I�y���5wz�*M���}�Ko� 7��y�6���� g�<%�d-��	�h���	��e����E��*,	�J���78���Ke�o�6�.��ō࠼�����;����ܥ�%�%eBH��[��o2YWP�5���J�ل���FO1Ĩ��#&XU%3i �b�T�K+9�s}��� H���n�8�F�e���h�a����0������u�,��`�]*>g�w�Y�nh��6�#z��x-pe��_*L�2����m\���i�_�������)a�"�'��k���gI�lv�f�z�p@*I�%�h�+��5��FL:�}�bl���)�m���}��+:����O�P�͒�Iz:%��o7�9˦�a\��JN{~��8���g��v�'��W��U��Rh��Û��S�-�%h�����vF����(�fj��{'��7~�|4t����ÛE�j4�m0�&)�P���TK)�V����w���mC��RCܕ�va�q��\���+`�xTR�T�18Uy�X���9�`�˸�Θo"u<��E�N�ɣ�A٤�d�*[<\2�\~)�R	f�Vӹen��$*�z�ƘHaMa\�ꙹ|�f�L��5Ƭ���s,4#��T٘��Լ��"�z枹(�>72�&� ���bg�"�
;,zV^���ނu�bn��şU��*x<ɾFT�t�F��mD�@�2ߘ"�?�M�7\���ЮG�䞌�4&��
ѣ(g�b����D����X���i��lU���������\K�P`�&�������8�e��Z~�����4y��H�������q�H�m�M�쪐I7�c>P�y�Y�����&Ǖ��Χ�j-�N���*��GMB/�,���?j��l�&����9����&�� 3��/�:��.�C��{�_��-���u������Bg+U��<�K�q�)�=��D�^]�M����8�|P�G�g��^��+��,��+�RT��t�f�u`�8�:K�^t"��ÛW5�<O<ʎ��X�єo �i��6���2Ϟo;&/�tg��7��
��TҝV��y2Z�{�'"U���=�����>����j(GQ���g@�_�j�o��l}�$P#MFN��_�HgƜ�~K�kMQA*A�밼�w���h4Wӯ��XƠa�: 6��ռ�|p��S� � ������V��q���/
�G���3]��>�]�qj�(�U|��n���.���6-�U�k�*�H�)+w���"�\�;��:c��XJW5N4ؗc"�2�f+sL|�͓�$��߲��3��@w�!�;rF��zB��,�vX�3g�wOk��
 ��[Y���MBLݣ)����Z]7�G���aF>��������͚�;��ga�m�K#�$@noT�ZDLr��M���)�80�D0���{N�?H9��ufb/D��$ek��V"���Ʈ=��{ ]�H��;�1��B	�g>rxn��4�4X�>�F�9�a
�ŋ����ռ�!�� �bD|��4�NIh��'��V�<V!�#O�iD�Y�k��6l����%P:R�.���U=K�b��Ӝ����:4�1{/1?#$0���較@,�_�3Ù�t�z����l5�fp
]��s�F��30�nm�L�i/��\�$��5:pm���J&����f��J�Ф=@�ڥ��PK�<��t�}���`������wI���.����$Ec[q!��6��,�����m�K�K|R�������*������pB6�%ݶ9��	�A��+���Ou��>�����Òi�#d	;��#Bj�vq'U1�xAB�$�*�eiD�!��g�N���Wo%|�c/�"r���
�v��3UZ�2F���'�Q�9��N�䲜��w�!!#@�����-��h��
7��l�	!M_8���"�(��g$�Y��@k����MY�I�_����4�+D*n}�M�#�C�KKjӤ`���x�*w8��h���Y�[�� �E&�P����M�A}���#�|=��n�>J+����Rd��Q,��a/x�Q>]���)W�_r������cT_�@�f�z|�|c�XK�zLZ�\N�юŎ9�MՈp��'��#�"�>g��֋ A������E�����<�.��֤�5��@N2L��
�;^�R�⡫��ËdYUB�R�j�)���ϤڗN��6�2}����g�83KN���Y0��?f�8�ѳŸx�!��:��kk���j�����]]����~Ẉ��W��%.���+�� ;���"��}����tz�B-��~X��tyI�5�N&�7�I�BK�$��hR��ؠm����gr������Ë)6�<��;l�2��*F�56�od4L�&�W�Zʋj��_�j5D��rY#ܞh[��@ӛX�@6��w��Uq-uA?����u�.�\�q屠��H=١���������أ��Ka�p��oU��-'zS=�r�v��Ԟ��Z~xZ�iBn�r
`��K���X̠� 1�y��&���*��������Q-ܣxp6w�ͯ�j"��_�[�T�
b�]@E��Ʋt�Ώ��T5;�z�] =F1���bQ$�	��1A�؝[1���>��ༀ���<��>!�eg�X+�J��FJB͠ި�{il�OQvx��g���'�D���������6��R��|��C��9{�:��6S��YK�<���ϻ��t�8r�)��"\���^�&���s6:��j!>��[�r�9��H~b�+jd���2p8�(���Tn����Pbg`�����ek���	��D3��k�.��o=�8�mI�v'.C�t�K�8�YX_U�e�Hpr�ʏ���.{Y��� ��]p�)����~�͚	O�m|֔p�/��!)�ߎ�^:��SO�|Ȗ��z��ሕ�6�u��J�J��P;�pB��w�k��	NT���|H܇�1���u�튪��%������v�CJk��@�N�=d,���?�/���M��W��r/�|�� ZI�8�|e�t�4٧��-i�Y������:/:����9�,�]V�Gh�bW���50�
&8�Ț��ɾ���O�*J8��y23�#x�$��@�Q���[�gg����iT�G \8�Ch_s�!Yw�(�f��п�j��Dp4����\��lKr��V��ӧ��"	�B@�N�
���*��|�D��"��+�򙜌�����Zd�S��p8 $�w�5I&��=:�d�Xjk����(A���#u'o�=����Sk6^�p�&�x�ЕY��3_��p/�� Z�1r����Zp��\����b�������E��P�ez�#R~e�+nC���4LXhsy��d�	��XŪ����6�~���l�����w�Ͽ`�����ň�"�2����͚?�c�C(�#Ac�;h�����"�8^�1�q���ȩF2���2�Q��A!�n���vAŁ�D6~C�)��Z�k�S���.�oЫ�T�mU�񸝾;���>=(�O~si�T�=��9�������H���zze�t�vt�&B���w���E�#�T�	�K�A���!��&��X��4���X�w�&�C����AGD�tEܕjuX�����p6��>G�o��C�vȻk<Fz|��^���|���
���݃�
z�A�5>D,A8LgW��G�7���h9�?��|����[p�"G*qUdx
g�ހ�� .�{�|����ULdD���.��i����\�g<�7��Sߐo@���Ҧ�;�V�P'�!�1J�yD�5?�E�U~�#�zvN?Y��hw����Ca�,	N�?C�slԽx�_.6������)].*�k�yy0ɢ����L`���6�ߖ�����}�,����e�|7�������D�Z�ba�P��C�v$�a�i��7��^�7���U���s@�lr�٬�%�0�~9�	���Y�6�:�}���Qw�0���a='�:YM��gw�
ΰ�bT��s1�:���U������[n>�C5�7g��&�*tp�:���3��P���I���A�iv�z� E����<Pd�Z\e�y�+]o%3ޠ��W����5���^�]P�M�g�9��~� @�|�}XW)���B���ӗsQM�69lۅWΕF��<b�~�Į=��cm��ۇGu�(��f�^�͎�oR,n�����:b�|���%¯+�lt�:~��ţ��s(���X5^S�n����t2�'4���4G�2P���gҼK�d��@7I���싅�f�]�r��],3Z��	�{�	�߾���
�����:r"�$h�*�ko� P&&8�~o����ubc��1=�+�ROI����.c�/-�n٤�'�q�����K�t��J��<f9:�]�Xz�� ���f��7����í��	0��m�K���唬�z��EǛ�H���)6Mk�"�����ؖ�N�YD��C���YW�NX� +6M�G,k�":[�׻�F_�:��^�'6���}9�6l���k�����;�􌜯��:��C���t7a}�򥮤������D���e���bD��%Q�F3`�Fn���)gJ����ڀv�7���rj�؋
�����
�a���!ا�#݉��j=�:�z�*����w	�_���� %��ή�ۿ��M�[-��,�ڕ;��D5��Ben�Y֙"d� 3/oc��0b��k��d0�$�o#�����d`��no|����Kͬ��tG�F�[w���^���Ghtw4�^��E��^�^G��
å8�>��c�i�,.iX�V����L� dp!�]�m:#ҟ^~����� �s����O%���9r��4�m	��^���"/��Ӣ3: ���ǩWi�X:��l7V��(��n�[I..�#�`��c
2�Щ�398Xۨ�Ш�,�n�z��IR��w���0�ګ �>���C�sL\��:n� Mg�R��"P����7��������W���y-!���ʉĀ�y}��A�?ҴcS��*ݎ@�� C�.���B�C�a8�hD'��G�4a��r.������&�'	�O��a��L/G]�	|�;��N����S�����\ 5%6C㌹�#�:D�=�Y�?#�.��"1n�����4JVA����S�Gr5�av&YK!>yA���z�S�9Z�� ۄ[Аn����������G�}[qyLN�a�s���~J2iӗA-��0�C�-�l��R�h4%0<Sy���m!#Y �4P	4 ��-�~x��.�]�o��ʟGL�[瓡>}���J�'ޮ����764���0�T��ݒ�a�C���$^���M��b-��}�SUD�W
�E�c��P���BlX�=���ӻ3��z�3����1DD���)�Cէх=�/J�b�BK���K�w��'��>Α߬���l�������4K����6���|���S��YZ�n�єO.mތ/2>V2�O�# �9��)!'�V�@Hf
F�P��K/���iֱY��i��`�B`c��Z�l\?�pg�!nDݘEk���Εk�5L����,�^���ڭq��B�����&��v�Z��Y_I��Yc�����ԍޑ��"�w�Ö���rMV�S�Lw
T�~��,QD3=�L�)]��B�y��+A[�}$k=�לkq����`���l�wsn�9����sM\P����e��{�6`;�k��1�L
���k�iE�ux���c�3��eZ�>�{pAϮ�P'�'�X�"f�$Q%8I�.H�X$�А	GU��J��*���q��I��2i�>�O��;,H�����8����JL��ZX�ILc
���{��Z�M��-������Y �4���II���hȘ�w��K����I�y!4��RTkF4h,��w�W�!�!d��C`h��̌�x�;��e�v�:���;.\�������d��1���%�%p_:�N����R��� 
�Y�k�+-nܥ�&=+ˤ��`�MK��h����UQ5�o�Cw��ؚ�*;����`�tm|]���Ʈ%1�;��?��a�P'K����a��e?�H�W���~�li}ڈ�F���������u_�t���L@���p ]�up�#p��y�S�Q9�^��Y������F��B����5տ���p9`t;��yK��!��`�G���/lN!T������G�GQ�%�����RgH���?;k��ܾ�N+ߋD����c�)��_�>%��$4�Y]	��K,�#��q`�)��j/a&s5R2��� gX�d����@���5� =�0�x�w���Eg����!b6��-6���OJ�4��P��
D�G��,@5�g��2�{��G2��u�N���\ѲW}��UR�S��p��M{u���V;6@�:��/��[��N����/���s��ʁ"lq&��/xm�{Qq̄
��,�>j�莗:Z��/R�c,���0�K0L�֜s��c.r��W��jex@uP'�o(�*���:�}�����mb�'_��� k�!}:�sʭ�eD/�AIƆ�1��e5ג��4[��}�� ���p#��d���`�t���s��-�3`m�ˌ��ϊS>ee�b�<�����[���� ���	y���쒂��͋ŕ�>6����7��8�i�o�u5�����D-Q�o�Ζ��X�����S��T��i�z̴(�%��҃\�^����o]YJEEu�%����ky�Ժ�4[ו��:��Z���Q)Q�΋L��8��l�ȣ/�dOû(AH��+䴧�u�C��D8���'%(ԫ���(�������,�?�+��"��/�O��@��'�l�l�p�A�H�w�pW^t(572�LY߼��������\n�"FS�B��(� 2(�u���o��<|υ
�-3¯�����
� 1�x���MG
p��qqG�;ל\)��j"�B������;u%8��CS[�34���Տ��������[��$7�˺��-Fœ�Y� �⟞�D��DQ����:���y�1c"~�$MA]u�h-��GJT6:�Dq��X�f���%+ˤ�N� �y�lZض�8V��I�������/P@�,�}LW;y8\�Xw�@��q^�,F�����������V����H��5�P.]�S(gұ�ؕ��ד���Y���w�0!X���V���k� �<�C��f(�������
64�Tl�<�d�:^j?��8�)�	�ԁ��l��Y�2��;������-<cɊ��˗����4o�'���@�KF*���C��O��w`�_�*Z���S`{~K(<EX�r��7��� �Aݒv_��v�D�K�R����Q�ǎ���<FTh�jTa�� �2�V٦F���·1�ڵgơ$�f+ƒ# �Zn��f����	0�ٌto�:�"�n�����ӹ5*���9y&Hj�#%��(�:�w��~M���6���r-U4�.`�r�~ms���������\���ұ���v��-3�*o@�ǡ�&�R���o�vF��Y�s�>����y�,]m�/��N:��P<�r�:]�p�ZOa8���u5�c򌉑Į��0����S��*H�!Z.��)��yI�n�ɏ~j�n��2@�
��H���ڎA�7�i�ZR���~fz��ˮ�[����gsȹv}!7l�?�ˮ4�;=�$}Z���Oz��X�7��^
�aG�h�c�#S��F�_;�Z�����ݥG_H��R/�2�]��<�ߊ`�R�Ej�Hq��˾FY+���;��o�w
�$�
�k�R��م�����âk�P�+Yʝ�N�?�OK�F�oI��=�0�g�W��!�Ig���r�Ӄ"p��л���o�J���ʵд�?e����h4g��Lվ�� ��Q3�,N��z�u�i9�Ʊ%��Z�d�O�i&�v�5L�oVu���[X����-�)���;�\֣��yfq+o1��
�'��~���D�
<`J��.CØ͓]��y
c�
j�	q,�XmGM.GG�LW�,t�G~/~���ٌKߟ{��AO�w��=d�����jC�X]�?���	�(!N��=�����9�ܛ�),b � ��.}d������U�j����u�2W�i���8"1�G-�E!��ҟ�\shb�)��A��щ����ꡅ���&��6k�ɸI�H�{���ȍ^�K�ɔ4Kgx��g�h]{�!�^�Q"1/����S8��#L��n��A}�
��F���10��K����_���+���]�Gtq�})C1�H��1���R��0\��ޒ��w[���j�I�M���8��5�E�hX�*C�C��eDw\n��r,ikLU�E�<?�� ʺ�cm+��#J/�b��i�1٨�L� ����m*�O��8��ִRBi>9{I��#��j���m�H�GБ��Q��"e��T���X+����\#�Ui�x	ӆ''��v�x����4�u��l��ej�������^��v\D��$�hW����rE����\[���{�̧�~�S=B�������D���:7�'|?��jl'�p��r�`d�������/�����0��^G��G+՗��)��_L�ⅳ��:gd�����bt���E�nȚ�i5x2��bE��Ey��z#(��߿?�a;�����D�A����N���=�jf��{W�h5$�g�q��Qq�_�j޾Ԭ��������H"�/��lOe� ��ͅ���Z؀�p��fLϴ�8�x�r%Z�,��j{U��j
n�H��y�t~z��߯@�_�:�<�d�L�'Q/ѻ3�����CtV��\]edI�j��O�&�ZuZ�Ȫ�2�w4��H���+vC�{���5�NT�l��S!S7DZ����,+,tR}��=D.�jg�C���'uc�TEVq}��m^���F��|�k�c�Q���r{�jŒ��m��3cQ�ߝ=	7�M���O�3an ��[��<H�����oо�	uj�At�|��v� ,��ќ��xަ���]'���G�b>xfW/)��/��d��/Q�M�n��3�E3���M�I+��;[�KG����Xymu�
�{�VA����\]2�A���6̀=���D�G�x��h��2�y�Q/��M?���� k�������,j�`��L���;�6坕|	��Aݘw5[��U��僥�Me;#�ߗ�����nپOm��?���&�Z,�!��|^ ��	jX�za$Ohsy.K�JQ���{�Ӿޘh�s�9�X[�7����u�dLK;��w��a3�H���K ������{<�$V���'�$�R>^�e���Uҝ���R���Q�ʾ-x���q-̜�]�(���o3�<=u����	䙼}o�Iي	{�sW�w�2�s�k�U�h�C*d�۴��y��f�P����_�Pn�a{&�ra��
��~�2��\�����en�l��j��3b)ɳ2��̑૵�A�f�HFq0�'�rd���`�%e<2G@M��-ۣ6� �e*na�Ѡ.�~��a�X=�����<`'�������\1�������n��g>D�t\��ݖ.x��e�#�+"2�#ܟq
M��aK�L�Y��K&`:���f%��+0���>��5잺��E�s�`ҀSe�QtD�3lV<�k'��5�P�j��K��!&ZФ��%�6{�-�8��~���/����$G�(��oܽ0F���J&�})��B��,�� 7{${P��/b���4:���8^�R!s7��-�8�GL$�l\�=����׮s��t��:&��TD'J�Tp�e$e0��0�v�E�,����U��p���\RfV�q��y�9�p��rҡ��H��#��j�,P��F���y��O麝d�K}�^?@
ɩ�*s��PC�9~/�"�_�U<h���2�a��s��F�$ux�����B&�iç(�<���WƠM�;>��0����#��je�Y���Քf�?���2ޫ�Ҏ&��z��ƥH݉���+�\`)�9I��lrr�JXfp�+r! �� U&�X1a�Ni���E����cn���/����O�C,����Z~eK�eMv����1M�\����%����'ڷ��@ I����.�Y��!J��Dw �k���X��-�J��Pb��K4/��6:�a>����ѡ1�c��D./���uh7�l��R	��{{K����݉��+�-pWu�:!�w��x��2`�~��d|���GBN���e�b-?�C&3�Z�aiE�+�mt,6�
�l|���Q��6�3b�7 ж�� �MK� ���CJ��cމ5�ڇ]H�39�A��z_�*�o��Vo=i>O]���n�'�	&��	ȅ�A�@S�!�5��Im�TKJ�.�)b�i�X&�w�c}jO mZ��ᮍ��|�߀�0���f.�唫9�Q���p�{��,�D�1��� <���<��!�i�
#�>�&�9&��F4�A矋���P�W�V�Q���̻��G%��*X:��T&*��n��"��]��̚�۳�}i;��Y��� c�\ֺ�����jWfBl]� h#L2O ���N���t�f*�'�iE���m��!�*�AF�,!��/��`���n	�o�z�{�B���y{ ��p���\��r���1)�~g�rD,����m1�	D�ITL4�-B� �h���u�k�%O~�pI���w�)�4[b#���i!� �v�#rᨗ]U
�b-ʆ��FvN�[쎴4j�/��� ��)�3�ST��`�kZ;ۆP�g��3l�E��ׁ���Ǐ�rf>p��Q��������X嬹�|-�� ��	[���(���	#Z;�����\���:.@��V���ZD/��s��A�j-?7Kv���x��NĠ������q�S���\Oɗ���y�"w�B��*�[Z�=G��v-�6w�o���^K3�m�_�9����W�,�ݫm�7Y,�?S�1i�5W_XTp��wL��8�	Zw'�϶����hY��x��dEp-Y��G���tC�T����#n�v��q�t7 )Ү�p>��tB9�/l��CY~���W,c�^2T6�������ޫoG����D b@���옎�D��#�i솣�X+� �>`��V�0a͔��Sq
j��AD���&�\�8)%��w�k��b�hG~��<0�
JU֡YEF��ur=�~�,�nk.�pE(U�rX��V��]�����4�	;�r�l�p��*��+t�d�{<
��'[�����X�qg@��ʨܿ�w��6xz�BP���`��pi���R)��#l�5>0c��������f϶3�Qc����9��n��S���ń��<I�,����d�D��E/W�ę�K�,A��d|?Kta�˱(͌@^��]=$�����ȕeh3!��瘶�2��"n"E#�J���Q�6B�@L��-�|�G�Ѝ�)�0��|w2�/��HC���S���U���L��|��#�!>h~6*���D�	&��<9�˕���\���'D�O^����&լ��+�d�ꋶ�8��x��\���{�z��D�Ar�tA+�^r��;�mU��&�� �a�(tu;��m�Z�� �����t^?O��7��hS���u�mW9�G|I��V������f��ႚ��.����_Dv���r�&����尸�b�P@X�ӯ 3b��;�	(6��-��q_P~ �U[��?i&�Ԃ�g*-�!�_�z�~:�d~��������0w�>R1B�ݭ��X���c�uf��rj��h~7�69�!�H%�Hzu���^x{�B!��GX$��v{l&��X�&���0g���>�kUϐ��ĭ��")D 6j���'�����-X�2�S�L�x���٧y��x_��c�~>���~�[.��:����3ې�!���7$B�^��xDzы6J��s#�L*�G��P��N>ϲ,EH��˗!G���nU�pp��>֝��wI�.�\$fo	x���Ԭ!9m^�Of��h�~M�Z��7��'�E�@�7y,Y���������O�ȵ�L#S�yF5�*/BZ;L?g���Iu�w��brL@�v��^�2ڛ<���rb�O}w�^Rp�5{9p6E#_�D	�^�<|7nW0��nT&�������u`R�7���e#�I�p����4>���0+ݜ���v��oa:1�����Y4�W�	R��o0�;�c���o|����l&�A�l�lL�[]�r
\=��M��v��`�g�pV�{�.��yZ6z�B;K=l�趐�I�8���PEm�ز_H���U��W��A�;�:1�������, �5��`3�N�U\��Qe�F�#�@��o�J�2�B(.�� v�KG�s~k7�>:ON�c��+�ad�o�w��M���J:���_���όw�Կo��1zD}5Z�2*���WQZm��:0��9}�ˌ����Ę���-�ι���I���(����3h��1����������"�c�U�4:�)�-m�sjh)�!��J�_0<xaU��g�b�˷qo�:��V�"����CFW�4����AQ��'o��Ni6����(�,�8�N ��|�'���u.mwZ�l7�.A�3=
%�ܾɤ�F�\��^j���%����K:�'��P�� e6�܋1��(���}������@��M��+��O��x�>�%>M��� ��&��d��QOD�O��79��y ��ޫ�;��z�k~�紑�0G���G��kWR���T��v�(2�	UK��}�v��}�wOXb��C&]3�������҆f������W��@�R�	
�=�͍�η�	4O��г�6�yc{�h@,	eU!�[ ��`�S�2m�R�tيϗJ���4����_d�SJ�/��	�� �QmQw��O1e�Du!�Q2F�^�a'��z��&���TQ��1���)�	�z�W��蛐�B�"k'�.8F�1�]%N-xbs��A�R��u���79�ChrY��
��BA&��&�+LU��Q�}Y,rd
)/*g��~<��u�$��b>&M�Ũ�v,R���L1�B�Up���y�rP�avm�Z��9?%�>���gp�WT�ʋ�Fc�p������;5��Wzu\�M��0�N����H��}Ί�侹ŕ8��V��Q�40��%�Nh2�hJ���6��ዃ�*	�͐�v��\@|�L���t�f�Y���e�\o'��V9�/�d������bJf�JTԼ|�X�ˑ���k]�H2$�/F��2�j��O#+g���J�xz�Kⵖw�c��y:M�s9v
ix7R6�}IA'w?9��[H�ȄK.[�F�V}1 ������G�G���93Ѣ8e���B�RVe*mOV�!g�t'*�]5�Bx��DyK��z�D��R%?3S�w`ag)p�Ҏ\֓��ߥ��2K:K[Dis�XU�s���$��@F��`��	׵<܍HR��)�].�C������zi��8#��4���?��;E"#�'�Z{�K6�D��>���cM�eN�L�Rb����a��d9d�8e2��K�����L��͎z|�����(�r�(g���3{3m�`S��{ك,��������x���d��������J��G��e,G���On0G�� s�L�t3�Ö��'|�Ye��e���8�l����Ć�a��������ˍUY5����|\�D������V�VB)�DM�� ���E�?"O]�y��n��R�ȮL7?1��}����$Ϣ3N0�/rƴ;P}��s����>I��5�탃
)Rcn䜎{��]��ߑe}'O���mv�˜qe��5�Lܯ�.����6;� c���s(H��*��9��@J�D��(R4%��~���`�&-��όL�%b���$��z�u�����ŧSwЃL��=<d��k3�Cd�,[�M�_��	aܘ8�����6�;����9�:��;��/B��+�mf���9�5����9M��(ӂ�l�p��Z���Qu����e��ߋߟ*�'��(K��+>��˔���x����R�&e�������4�6�S�S��7�%�~�`y���j�$����͓#A;� Im�����=����<�QΜt�@��Yݍos�����6��q���8�L�Z\�m=tH�� �����Dr�_��=��
�i X�h���\��Fz҉�g�?LM�LjL� ������]!����q�Q�j�9�2���&����ܗ�b����Y��?���؀�'���$��h�S���]�.2�3���f��c+$��$��Z��w��xW�{Onb��Ϡ��~�0۴��l?7ϖ�)5�ߨ^\��#ne�jc���X����Y>+������g�R,�h)����%t����#2Q%����B���Q�u\���ݢ���ʹ��+Ew����{{�Ӱ��򓯋V2Ư�k�m�+BI��j�~�� (���V�������)�����@EE
���4&����0k�")K���m���UE�<��'y�ʈ	�?�G'�N*����*p�[��|� ,��p��k��7�S���Z �����;��y��N)�f�9����7	Dn��H%1��^zt�[j�i�\�@^��~�3���73�]%�+�W�ׂ4��Lޒ�G�錑�Dy]�)��`�t}��R�`��k�n<񄣨��K��[L)����)��b������^ϳ�8���oĆ���Q�PM50@gH����n�**�6�Qp���[!��c�S'ϲ���c���ԊJ���e�#� A��${9�7l���k�m�i}��Ͻ��כ"9
�g�fcZ����d�sꔁ�'z Џ݀hO�P<tq$}��L\�Ly_�`�g�c,�]�y�>���q���R�F�8�3vQ�Z�غ�k�I��j��M���7N}6C�K��-M iN�dN(<���y����X�n�*�t���C��Aj� �ި��/��{�L�ּA1�z�
_��_�˴����t�Зu�\=KR�d.�^sf6��ߚP��p��6\��0pv����HD��3����R�. �j�� �D�8CːPM�7Ή������}���o")�A6�eˌQ�RjI�U��1�0�v%�f�������#�<�/nV\x|-(�K�Z�:R��놹x��I5_.7	���7�\Hq�ճ�?|3j�]�(�����/��o�,��gWd�D!3c��0|�����<V���?�L���'�*��}+է���;������] ��C���}5��~GP-���"��|���5���PS�ǒ����)`Wr�mט��:Zk&u�f@��:ة��?�,��]���|�bt���H��B�������jh�벰�%��+X@9	&,��c�z�0$�b��Z�뙔#Xx�c�A�O�}�͎���ukd+^�E����D��U=?�L�{#�����	��|0�a�����߬�i���#�D�*���4�.e��.�O})?��b��Z����I1%�����%�h��M��ѱ�i�O�1U^K���W��{��4��E>����
5��w�h'O�[@��n�'���W-����#�c�Z���r5#�2N���d�N%Ǖt{e0Y�[��jr��y��D7rr��gp\砳�ףn%7%��t�*ɍ1i!�i%�����>�;��
iu1�~^�Sh�f)'p;H�3@�I*���!�q�Į�E;Nn�B]:��^	= ���}Uk�:��!%����l����$ZY
�y��[9�P:�P�x 'P��|��{��i�l�z�I۬mI���ז�G}�G�MGR��˴%�=ܾ��0Z�5Sy|��9�|�t���,v�U��d�y����=��>���i���Щ&/�n_ҬxC�ЩH%������e��4�s�y�����d�ؙ�a��FكNQUVL�����\[I�NXP��&�\ ��E~��|8��!�����.c��KD�NyѢe[)�}s����Z[`�wFDu>��o�U�8�Lh�w�t6��.f�aV����w��qq�������x_w_�u�X@���"1��X\[��Qػ(P� ��͢����;����;ʺ@��[	��m�A�$�_}O��f{后��S��L�@Lϔ��6( ��켝ŀ�j3�O��b�<,(�s�{���A8�AqT��!��%b4���&8��O�-����{��,�J�$Igd�wΠ;X���%��x�Lo_�?�$�a'Q�=ҟ�@�+竈�ڑ@���5�O�U�O�<�7�;:����d��'�1�&�SN��o��ES?8S���+��>k�4�ـ{'J(x��klϰ��{"�����(���
�T<�WPS��1ӈ�X�ö��ŵݎ��4��_P8]! �o��Ȧ׽Ux�/�?���?��9�@���V�� ���&�J��Z�~��ظ;tBL�G��4��-ɾ�*��8V�
<j�����ݐ<>~��+� ������^�=Zv6�ݺ���i4�V�1�s��VQN�m:0R�])mV3X�LΙ���`�뚅Q�x��V8�Ĕ1����m=f�&ջ\�a�Nv�t���9�(]z����0BC<o>r�
��( =�,���*/! ��u�*�uO��wϭf����ocs�w;K4�%ű�~_��/���;
M�b��	 9�c��-��]��+����c+c�
�C�]<	>��N�
h���8�-ʫF��W�z�q��P7�\�#2`ߍN�y�ˍ�׼'��6�N��7�ٻB��R1��������q	�ȣ��C�4p�����_&t���f/,�3�t��&��
_���&��ػV�9�h� 0v���l�ד8��D~��̹�+?�=�C�+C��ԯ�X-Co+ȦnY�p0y,�V!-4W(K` 9[���P���_҉=zN]��*q�-t������lpZ�Ñ-"�onw�	b4�A�����\w��#Q!4;T�
�&:�8�,��NWO���t6�F�P�W�v��+R��f�S砤~�m˞^d^�~��!HE���;�3����M����[R�!b*������ȓ���K��8�!��C�NX㳐���+c�o=��C�4�s$$�zsԕ��)fω�Am+�:F�z�����=�ka ��
��VB�Qa�(�D����}��"U�#�mV�	��V���^_�2U���i�H��Z��ܕi�P޶9�&��!���5Gg�ynD��u���t�{O&��^'a���0.dv�Z��X$�W�/ک��A�<����v�n�k3r���Q>wuuR�M��X7Pu�=�oT���+Jo��g�f0�Wݘʇp�#	�uͻ� ,7�ub�w{Q��}g4�2&2��z���u����G�L,#)��_��i%��T����w)�!F)��*?�ɨ��[�H �Sؙ�E�%&���e�h�� D�k���,��k��o��g�v!�dn���@�7pm��0�q��*��~J�]�@�#��v1�qҀ�hg�tqѰ����oP�g>����5��'"Y6������:l�=�y�?�"H���
lK���h�H9�v̓%켲��նDj2ĆRĳ5  ����%�Ie%\��l���T.��U>����\f��@�3����,�s[��B,0�<�<�Õ,J���^�_���Q�6}�
�?�~I�hI�����Zy���q��rV�r�a�+�o����k|� ��`L��W��J�������^�>�ch�������M����7#�ZO����|܌�1�?ls�x�`�N�,r!ڡ_�tD8��}�5�90��0�����	加g�d�959�,Y�"3���U�}J����KMU3\����� T "�0�!T��lt��W��_إ����<r U�n����]=��Z◑�a�^��d�].}���9w��*����9�a�Zm�����z�_Kϣ4���� �����Ia:T��mF�L��8n�"[�4ȑ222y�ŻVk��&�Ft��Ot���^���1xHۗ�f:�m��K�ZZ�n�Ã�۠y��Y"�P�1��ʎ��â��U�"5����(�J�w�g���
M?���P���[��R���=<�(qq��9��I��Y���/9�*jo��z�R�Ф�Bh�qZWE�< ǩ�ͣ<.�	+�p����$�_�R�8���K㚵bx��S�^+/xq3(���*g^��Xk[lWa�M}�a[������"x�V��5����*;�.j�`2ݦ�q.b�Ack�\Y�hyɜ�>Q$���������`	��9�ڨǖ��W}�2&�z6ٗ�Cp��Cd�� �����R,g��[Ǜ'1Y,?��9�3؈��sAr�.5�Y`m�֣�|��+�̷#Pʝ��)HD�M��̯ͼb�q"�I���)�	=�!�\��c�2����D�R~H�R�� M&�&�:Ba� ���#���]��u	*1��ڷ%�I8 ���<�ép�W���� �y�� ����6�n7:./�>��q�����au}��H#6q3�Q��E!22�	��P���^�Ԛ�D3�=��.e�A���#�J�.P���`��W�8]��wGஆO�h�=뷜;�+��q;���Ӧ��g{������:�d���@�.�S/���"U���}1��	���|���7ɠ�0�Ey@����r��֕��yh�yd����r�����K,"d�V�%e�qy�"c;@K=H��Y��Ӑ��&?(�½�`�E�󢠩��S��QĢ���Hev��Ʋ=����p�!�B5�JB�
�X�Uw�e3�W���^xv��Zҭ�-\ ��C�b�H�	��-�m����gdR�ul�@h%��S��@�K�k���e�	<��j/��ߓ�-M��GK:'�I67*ݍ�S��T7"Di�XR�H�UI��7�G4w� ���wK�2^�
Z:42,ׁ�4`?{��{?p5���Tˇq�b���&���X�d�CO {+^��
�7B,������$s7V0����85�#����}� <"��6���;ἇ�j��ȡ�_���$?����_:��3H���L~'<'��)�E��%�sE�`��O��E�CΒʙ�-4�'N��VF ���8�������]K͢�XU@/<:B����h4��m����kG��(�V��ʴ���G9!���E ���
���ˊo)�ߙ�p��	���$�C;�,�'�y]�c T�D,=3�Qq������<�Z�q�4�ϵTs�vGixb0��^�T�4��+ 8V����$N�h��<�N��pY��E�-�o@.������x�hG�FY�w^&/v��c�{*(?ҤP�h��c�z�˩Z�C���s�L���}�A�0�)������!GM��A
�=k�v#�.�51��>QaM{X����U�`�e��lx�oC9+��c�	� �}���e6�y��-W�T��� �>�i��U!�&�;V�k�sOt�D�3޾��Z8͓��a�ŷ: �(�)��/�T�vy�M�����r�[�}-���~o����v���{�������ѩ�]�ǖ W�̎��D�B��&����o�A�X��+���V�;�"�#>��k��c��H���d���J�,��UB~2O�#����z|u� �	z��i�3�ɅE2��y���]��9�[�N�u-���ε��gw�+�h�{ѠI�d;윸11���LO��H5m��͖��;]�*�6�۬p�	��]E���(wǪwq/x�	7�A�牪Y��~Ge,�Q�pu�k~��-�ƌr����SZ�I��-�'4!`�od���*��s��(�[�nA�wOf�|��6�x�'QAU��~eTg��4�}c:H�͂��������E���`���OX+����-W�&����~��a%1�� �b���J�x��9�GDCՎ��`;�o2�m�r��H��/��G����h�<���s���	��M����s4d�D�6 l��~��>O������6� rz�v�L9'���!���J�'�!�ɺ�r�^���l�I����t�F�|D���ַvH��V�@]��2&B��6U�h8"~-�z�U!k=���7������xo�(�qI�%����R݂�?�i2J;lti-^J�}AD���Y����w���xLo����`�w��'p�k{;n�X�!lH&'}^��]b��Vv⋚e/�ׁ���|4�ڻ�C������Gdp�*Q,���i��7��`ƪmz����ӱ��4�_�wZH���@�J
�hw����1t����TASNl�Hs�D=F3����-�1�˷�m�{$�v
�E;.M���Zb�!��6u\V�1ǘ^lޟYx�x~j����
���j��'��>U,���G(0��)`"��ۚ��h��Ad��[�����W�s�:�qT���#g�j5G�i��;`y�Ov��u��A&���W����~	����o	ovFqm��g���\��B�m8�A;&H��sp��<�`r5]$�R�Cd]�HmQ߅��^�}���m&��1�&n�#���CD}�/��vp�Î���3����O_������Mz@��70��[�ݥr��~��1���|��!��κ[}��ѓW�o�q���"�̢��ؑ�j��n��9��΍xƒS�������L�T�z�"��s�f}��ɞ�Z7k�X{�+s�/|��^���	��Ukź�6���m�!�Np��`�>@P��k����� ���\7-�.����N� �8t˦�pT��4�
MF�l���m-���p}�34ǂj�����(�}��	�� ���&�14j�_ca�0��n�e胓��/� 8�_F{~-������)���j>F���J�B1�Z�д��f��>rZ��?2�\g㝜�����$����u��#�i� 񄴇(x	@Q8,�Q<�u�(P��c�l�L�{ic�
^��[��f^�`�B,��հ�$��E('�����!C�M�	5p�H}�m�<�}4$�E(�y�W���Z���)TʥJOdr�X��{�-U�>{W���q��p�����K��$�K����20ܗ�qZ��QY/Q�Eh�6�u��-7l��yͮ���@d(�=�A�g�-k�x���%��c�4k�OJ��7C�C��鲺��(gq@�81@'(Wd�� ;,�߾D,��ݑ}�?\@���8��V�^�Uԏ�R�=�#[ܛI��*t���:�X	�qE�NIW�5�f� _Ǐ��"�X5?U�"yaX&��|�n���It�u}JO�v���Ɩ.��3C��n'20=�Ai����y���|G�#��K�! U�PN�R�����$q��c�ؼA���L���(�a�� S��(�$�����Fλ��O�F2��Ԓ��]i �Y�,�!JEK��ѡ�s�Lv5�f�E���p��|�Id�,t�f��:����A�� 9q@pH���hȊt%��>��׀)2�KtpΚ3���g��[�]x��u�n����v�����K-j��@���Y�&���^3(<�,�&���C�ڏ*T֐=dY��v�8#����|P|xʕKE���HdS)zF�Ԗw��1�BJ�K���qeޣ�5����*_GعX�B~�ڇ}�Uz��]���"5=joE�|��F3'�t>��A�G$�g��BW���4��<�<����r�b�_��ͦ��,X�h��X�g��ڦ!���`�u�`���ژC�.<o�"+���E��m������"���G�xc�#A��&0��lD�T}��*̫���v�$Sw�����s�'XE)����m��9�Q����	��8͎�&c��M*�tO�K|w�A���m%�U���NDP<"���*W� N�PVW�*N�Dk�G�4����'��õunGץ-��������Np�9�A�Jv���[�;�&0��c����w�����H�b{�ԣ�4p����l9y�����oc��S��6l�R�zSM��<���qtɭl��h�
s�+���Y��ǳ�R	߯ �
B8��:f��P��?O0A"��J�p�l�3���ʍv�������,7QR�-Ux�n��H��ґ�;��O~��Rd{D^��5ܶ�=�rݜ&	�Ɋ���]��!�q��VӐ�����fQ���L~��f�������M�:T�� c�\���;�ĩ�ML3rٔ+V�y?J_�q��2����{��[�@���b6�U3Y�y��\�p{5�aE/�bÂ��TD�v��5��U�@�p@aYV�)2�"�B��=�����+}��گ]������1��=X�'����
�B+C�å�ν�̉/~�F/1�͔�Q��	I�G[m�;5����p��<���}h	���]�}��ʗ�XbU��ja�ق���Z*�Ӡ�y��d��+0i�v��w�Ya0J@�)���3%<�@*%+��J gt��X��{����/al����[?���:zj�:AFb��@�/�:�W?rm����Ԁ�l�U�F4 +ۊl���<U5m�N�t@'��1�æ+�X�)�$:+ۥ�C����QD����~�3��}ј��	v�Z����+��������fw����Ԑm#@v�O�RѸ��hΈǡ�,����BC=�2^HW3�r<�sN��"���5%U���1{�ܠ��cˑ,2.9\k�#Pf�
-��x���=����{�F�<��Ü@���+�L����Khm	dU͋�{�?����i*J��~gC����~�]��aA�n-3$.Q�����e#�����7z�Rۓu�|5���,�$'���KrӖ�C��P�@���;� ���#e���֓ãZP��
����=6Q}Pn�V�-��Y.mJ�O�h�1�q��>�p@4��#T�Կ ��bϡ�z-�!f�#h�l����ҿ��M����l|��.y��ŬvQ�՟��E���GA�C���p��S����,���;#�c�~������K�����W�t��F��+��ي��%qAz��\�YC����:@�ޕ��Э�,{�����p4>g`�VEZI��h)���wv�4D��.�_��],�Sjpx3� 
ލV��>Y�cC䅄f����f���w{���� \�x�W%6��^��N%��␨ϝ5�"6.Ck� ��cN� �����_#P�9@+V�yC�2��:l~�ԫW��w�ߨ_e�Ol�}��A$�"��' aq��,�l>�
��]��^�$K�#A���H}1g�|DxD�}��@���B8�`�-*�0'���g�Mtz���ߍ�ݲF�	Υ�}$I��Ɓ���m�*�Jb�6���7�t�o�I� n�#���*5� �ⷪ��j�����s�Rt���]���x��D�;�Z�I���1PqA��b�|*�3���MԹ���փ-���ܑ�T���SJ�"4�H>7�͛ v��+p;�l�b��ݦ	��Pr$u-O��y�L�@�%�.�=#w�"��ņTA.��?���4%Yc��ɑc��I�����c� �Ko*�E��a}'��.$L$C?�|�}JZIw��"b�Y���I�S���Ԍ"4	\�w����u�+w���WLɏ�e.l�J��
��~���h7�ձK��*k ��ŕ^����D���)�vUW@	�I�$8��t��'�	�"�}����\H�S������@Hݽ?���K/�ȕ�c�g�v�ua`�A�V�z��W& !4^(%�����O��kH�;���2gCB�S�I�FߵJ�����b�r�<͕�`���Эư)9�5���ܖS��vhN�l&h����i�_+�EF��<	��a;�O��9�� wD�����{8�N��u�f�n'�M��WH�/�_#�ЮZ~ga�V\����z��,��P�/��-4���dZ����9~�kX�K�߭�\�;�3H�_7�(B7�r^��!2�^�A�q!�A��8��x�1w�2���YT5�.�>����?)���޳I�����Mݙ<	�eߠݘ�N ��as���.�!)q)�Ʊ�XB�4��7���C8o�*���'b�U��6��݌�|��k���W]ٗ�Jl��2�i��T�`�<��ЁY�3aP��`�O�+ 9-
A��+Q�b�&I-K'u4ɯ�Q�fx/<?�j�V=�-A�1�j�IZ�wj�ZE�̆�>�eq�YK��M{M�5_�xf�?�FV}w��fd.�5Z/���'7.�j�����a71�Ȼ�!Ux��4*�(]9�H��*�ɧH3��Ƴa������������6=
A�� ���'A�K^�������^��\� �	��e0������Thk��!fH;Mb&�jړ5��q?�y�~2��ì\ׅ+�1K�9�q&��/���z����G=ڊR}U&�ף�G�9�u���2d]�>������B��t/���k�[�m)l��NZ�����a�y6��\/�9�t��[��� xNL�d����'�5Iփ����?� ��mY;o6"R�i�I��qp��6�~�b�ë�&��z�ug*�Y"Mt2�x�~O$L����=��?Ă�3�䎧�A�@)���@�d�x���nթ~ƄvߜVN�0Wݮƚ�*\�}��h4;ɴ�ٗ4:��aս���~��#_�@<�,��e�&�a����"�ߎ:�I6b�p�l1�`�p7PT��;�d�z��N����!��c��A��:��U����׫:��w�0��8��`6�x.g�3T)�P�jLq�U��O:��h��p�^Q,�2����bNb�(�}�㒁Dt����س%[�y<O�$�0��*�H��j|C�96{ V|�Q�a��B��ߎE����>N:�7(��\2�(HM��6g�_:�NFsd��D�����YE�4����F(*~6T�(��'2�N+5�Gy�9��KT�][�E���$r�ܽ�y��J�[�E1��
� ���oX>E���O��e�dV��2�sK{A+���F�"O��M��i�\E���.C巆�%�/>_Ng��_d���j�Mr�����I�y��\+�D�@�����Q��?����:њ����
x	�nO2��[{�(W��+,�c�*)�Sa����'Ի�6�yo�~��,��"��>p�>9�Bh�{��{?ax���-�:1�5ʫ�C'TS��]ww�N�oɚ`;�/��x7����=�'�*�W6�
*wŭ�1\�<���0*��� �eQ�WV�˸E�j���#X�A�AG�$c+Y��]S��1pE�[]��<͘���;hs-�>(�ƶd�z�� �Xh��ܿ��	S��1��,`;%-�(�B�x�VI<�Fm*�ԑ�Xh*�`��:�/I�B��GX(٭V�)x5�!:zS�|���'{�-li �Au�����d>Pm�!a���Iq[�u��ﭟ��$���;-
�O�wA�9�}^�S���g�AKj�m~���:\����QZ�HL��ۓ8
Y���0i�q�`���&_�|:����(���*u�{<�E�������`F��<�B׻���N�6�)d��Xo�����n����v����_�Cq��e�g��W��Ԧ��E�Ʀ���|�?W�%2L����:;M2ݥ���i��ƅP*.� #�>�\,�\�� ��y�V�T��rC�g��Y|ma�cL��<�~��)l�	����oX,,
4PB�s	����j����sd�깭�/��
�}�3��tiO6ꐻ�� `}[�փBfr�D�q�=��c�Qwc3�j)�>s�*������������PB�D�6~�x�6�3n�؊c%���L�ݪ(��19<"s�;�rާ��Ưky=�����z��ʮQJ���:��Q\H%p�S{�Ы���~DM1����!�o.&H��w2��
�w�:g����ҼVq&>�ї��	��_v�Ϙ=������٩F�iCs�;�R3(H�(~I2w�5���� ��x~�uL��.!��_ܡԽu��a��"��e2��͑u��(�B��ÁQYɣ����pZ�F�7�dT������]��l�1?�q( �n����'^���Lң�Z��Wx�.�V8/����x�%ZU������b�d^�玑�o�3�2{�� 4j� X��7�]&�n/�y��T�KF[�Ղ�Zi�P cT��@ݍ�0D�!��0M4i���ɬ�W���a�����`5��Q��z����,}~�}ӌ���1b~���B��j�����E4-����B�݇��RA���.��"�+�k,Ԅ��zET�C}�:�{�W�T���M1�]<���iw�$^4CZG�QM{x��������=y�rbη�c �K0��$蚦p-cOgxܦ�@�تA������>E%���Foc��Y�<��`�D��Jt�C�U.��1[���-������ z�K?w��A,�L��`lg��}���Mι��eNG(+�����1� �M��]ge{�� |-�%����m��e��#9�o`�Gm�/�kBuFX�Y')-�=od�7i|�8:Bi ]&a"���P�^s�G�Ľt5Lz���o�y݃�Í�Y��i�x���Y9i��m�=���ե3�~�7d'�#��6��"F���|�i����p���RP%��3O�$U	@_���3�l��i����dS�Ӗsu()T5�U�94��)�y�}r�L)�K�'�	�B&̢�|�uJ/H2��t7�X��2�45���tg�����1+��c��r>��I%<���O�;��[rG���%%�\DΛN�NT(��p�R��]1!ΝB���sz�|A�'�s��I���_o@9KX�|�8n��@ly�}��]�>:Ną2x����S�������&���B��	�s��?��W_S�Ms��hs��?5��E@0E��U��a��:u˦��s����I���ڂP���+���q�̔g�aA
�9�6ٓ
{P�@�ص�.�]�lQ����n/���j���E��>3���S�K?L���� �4}P;e��j|��2\��|(���~"΀E_ #�Q"f� ����t4�l��&MNٷv�#s�kE�E���v � O���mM��S�����D��1"9W-e�g�zFr�\��	�h��#D��L�u#2��TJ��qdO�D-�#,��9o��^R��^{+�V��B���e�Ϣ��Ǳ�����襕��"����р�����lV&�IA�����袞��e�kˁ�\�E�/l�丢��Q'(��"-�30M �����g�<���<w��f�W�`������s��)a	Q5֝q�X�^�sȊ]{��(6wZ�*e�tf�!�)D'ye���4&���
/�'ګ�ڐ�%*Q���� �����=n��"�߽p��Of�v��!**�q�4||�\4��C�w�̃pA0���k{}���<�\�ұ(UWu-���f��:�Ns���(\�/s��y��7�Ԥ�]��.W�A�f���w�nĮ���s.�>����#��ZI�#n�22�&v!�6� ���*������6ceצ��M���6��ђ�X�{n�!&g9B
��j���Ƌe�V1���j�>��u�攸+�(LHu�2���2FJ<hN{10V3�z[�y��5r�Ӊ��̒�i��òu��S~\O��-����#�z[�Sȏ����r�IҮ
]�@��Dd��5V�u��Z�����Mi/�aub�V{�������2l�_��C���ܛ�Z�I���n�}&ZiwS?:��"#��]��/8�B
œ��ԕ���lV-��w�_OBҺ��A��l1A�M�����9���Ɉ^�Z�%M����c����?5�^
�z��E����`%.���ĸiD��O������" 8rj��)˲��,��G����gQ��8:�D�Ӕ^S�#���e�6��{j?d��y��ר�<���.On�7Vih�!�����ġ������68el����&�s��A�s�5�Hn���%Ճ�$�N鷉����^Z
��9%�I��A4��p3G�ЛGޟ�S?����i~�W�\�<'vA�Q僞`�m�!_%�( $u�\Oڞ��#/Ln����:lJs|DR*�zb�Hm����|�M����\~2����oΦ|+�E�V����h0P��M����y��).�J#Ҋyj#�Ѻ�	D]��Ϙ�n�RTt9��P&���d᳖�cѸ�46B$ʏc�}1�	���;�CM:�Ѫ棈�Ae�6���� ˺@��=`������3���݊e�2\Ϊ��L�>}D�Q���ıx�7��kԵVq:��!��d�ښ��z~P�����5B,�Ʈ��k���j��<�%�#fR��bĂY%��n�8���w�U�t�8u%�#q�V���O�)w�����B,�Y�^��:���/Ek�c�(YQ�lY�̖����?�28[y�lǧlf�e���$µS�ǟ����!+���{�,�
��8��b���X�!��k��M��� g���z���[�~4�X�<����A�MRL	�������.z�F��6����u:�i�m��-�_&��U�*kP�_��4ٿLpު�'�V����h��J�^�Yj~��of�2�L�7vL����fj�f%ۻ��S��ε����c���g�}@z�����:��U�S&<>UFP~Y��$
�T_}��(s�h'���c�1T���0�W_}���X̀zO��?���	��*G�jH���ֿt92��r	����'�S�����Aw�T�.V �{��V�we�'<��"+Ҽ�����@8�6�����I��cm{\���� [j�W��y���Q�C��krz�Aw��oWЀ���(�`Q��S_4��S����s|m�ѱh�ȴ�m7�KS̈���9�~U�^2o�7Df�"hA��O?:��7�����uv�Y@�Q��@f5W��Q]�����i��`��g��[bV�X�����,�@�"�n�����*kw��k��O#��>P��ɪnp�&x�y�sb�VV�I�є���O����51D����o�?*f�/CL�g�ٌ˴o�Y���Zԅ�rP�4k�Trz0�o9��~b!�a��2?���듁�.^g��K#���*n��K(�[�d���I�
���ɢ���O�_Y���JX�+�	\ښ���I^Y
1n`�YЭ��TAgs�f�_ B�b^��G�����t#��'�:ro<	{�\�z$1 g������^倂c_����f�dZ��aH%+�k��~:=Ǽ����z۪M�e`�]Zg5׌7���aRo;�y������C�
��N����A@�ub~�'8]Z=݈ǩ?Ś]:�i�k(N��~�h��>�A	\n+V6)uV�y�81fGsXчlb[;�*�0]:-'}扵����c��ܰ��7�����A���W���F9V�PcdH��!e�
]-�4)2\�:��ӷc"rш�*��9";�0�Y�B��+26�}��B�ϋ���2�n
�ü��K��,�ն��	Z�n?F�LD��E���������#X��0�ޑ�i]p�Q��|Z�O��(z�<��d��&𠡀r�c��M5������ȥ��3g��g�`Q���=�٤@�� 2㱶Q ��m6\W%��~k|	����{����&���/�������:[�D����6��8x�f)e�ïg
��P*EI� =���
�l���Nt��^Cm�D��kf�
��B��վ���h*�w�6�kuIuKZ�Y�������bT�v��X��%
�
���� Xy��93�LI\"$5�ңI�?�vH����qΈ�����=fDaF}"du+�K����fU�2ﶲ��Z�
���g|��pd �حc�/���Y�d��4���7�[�W�幽�IDB"f9���3���p�nDB��[n��rG�)�d��9&jZ�����f��r�T�|�ĉ}"��(��K�ebU��mU�;Ʋ��y��r��JP��k��:��~X�&�+R���fS�n�n�_8(��/���Mf���rY���_��_f�<۵ Q4�Z��"��bf[����b��Sw��9E���^F�	��y䫯�Sţ�a1���>�+)v�7�c+�x�_�DLfv]�^�G����hJ��^��n��Z���B��~��F:�>��y*�&��K��Rv�-a��c�H�:�ģK|����"��Vz�[��V�24x��[�`O�����-8܏�v���Zr��-�?LUގ�����!�ξ}�UװL�[���+��i
u?��B�a����hǚ���X�*��J��L���G"mB�Ρ|H����+�~@��@���q��?���TrǛ�l�o蒛GM�1��H0�s��
~��s���y0lW�.?b.�B}�V�K	;����v�e�7LfM+Ǳ}�'JbZM�&����t�����[*Ҩ:a�ɮ� �Y�V���Ó�y?>"���p/�ONDjw=m��tZ�ƨ�KFJ�D]>��Ba��?K=�mc׽o[�O��A)F��;�H���JZ~_n��/�ڑz�^�S�Ty�A���]���c	���c����q4�	�彇����y�3���J#���*�� �h�dY�᳦��j*�T?�p��n�Z|�~)q�w�P(��k�����#���f.`����#{�l�]#�I�����Q�XZob���!����!<Ƣ�.T�J�w��_�.�I���l��*ؖ��["�AѴ0wЎ���Q|[�OSX� ��[D��i.4F��o`>,Wn���4he���V��G�A[�3ؘ�J�ta6�,� ]������.ģX��}Y9�x��V깙tf!��Q,e�I���$"J�c��\Pք���D!fb����w�NZp]Ys}�	[��iܴޗN&6��)�EJ��v\�M��.�I��ly�.n�L, D��ߖ�8����F&.Ÿ��G8�I�������<yo7��ɘH1L����.7�K���YdMjWb�V5�S�2&¡�������K�U��\����W�n��\:jd�`/&���g�[-�i�tDL5g��3�9=6^}qW=	�7�����{wr>R�eT�4��W�묋P�"�1�ԉ�4='����͖T�0��m.�ж^�z]Н�QW��l�p6�U���a�a�a���� A�K�MG��bY����t����)��<7�B�4�z��qF�.Qm���UYY;�]��M�2����_T	me������K�2I�^,�'}N��
���/�2`(�ޞ�|�" �Z���MG��0�e��E-$����^#($t�Q�W�R�8���z�g
���E������M��hB�XeZk.Z���5I�|�� �����϶qHHUq&�v��7��`�����<�
r��x���X�G/y���1(�=U�lz)��+`>츎������Ŀ���	���G)#��PrC��o��׹F�8״�w�⸜��ʐ�|��|XB�B�o��r}?W~��v�eX��K�s��V�KA(� �X7=ā]�L<O�A����grpI�0����Q=	���d3�`	���Ͱ�P}����`g	  EAt3�Nf�����M���]|W1x��	�_��H��2f��*tT����>��A�`TIؖ�c��@�aG�m�d߰	���bA���3�K�eg�BՖ��s��W���ܮ�$�oa�J~441�asO|-�]�>����!�����D��	^)A�C�ş��`ܵ�h3N���(esʰo}��_�\���;vv6�>!����ͤ|�i�Q(�8k�3Ǩ)�����z�4��B��!'��Rz��@L,�}�Va��7��$��cv�iHcB���Sdc�i�[�/�Wٷ���[{\"��q&�ʻ���Dba�f���( ���$��#1�-U�C-�c�����>�uYF�{ `��k0E�$+2��Q��fH��'�yhu�ףn}@�:�`iuNn�ev83��">x�0�D�UŰ����Rodn7B����j��y�;��\�E��_���pމ��-�NǪчʧ�z<T��s���T{��]�̵��J6$���6�����u�OV� J� �C���R]���t~��0���Cm4�	&|�H#�G"ս!�C.�bT눕g���c�:^;�y�1��6�%\v2.0��Wv���
��2��	�qN���^aO�6ZT��Y�nƆh�B�:�����EUX۾b�U�	] �lF靏6�iCU�>�oi:��J��q���$zB/`��z���.|��+LI]��s�'ymM�U��+��	�%�5Nj�"���vی�q=��x�F�V�#��e�z����I�ϵ��gή���R..��[�>=+_���#�ONA�:990 G8N�h�NS���y 	Xy+�&Y���wfo7�����6A�ڗl �.���P
��&���ٲ�S���y$|�7��VP6��H�f\��7�MV��F|���^_�#�����o��Zcq������KE��{�R�I>tu$����d��cߴ:�6�g���e�T�fi��^=�Y'�|L�hPT�'��;���"�.��뢩8��$���20GE�
�䌧� �x�Xc4�hC������sߤKN��*���mX//1���Nf��2TȢ�2�Hᒴ���$g��<�CF����� ���R�!~a=寎�NYy���!��d������=E �P�M%Z�}�����h����ʺ��i�+n!O��!%�Jj�P������^\�*�.ㆿ��"d��}\�Ow�~lA�Y�-n�N|YX�~Z1��}EY��W���+�)A�ម��_<��,���mG�����v���?H�c��W�,�<��o��6OT�!�Z4)�=-Ѹy�nuZ�� �=߿�����/�zpy��~�x���]�fJ��;�G*���	�^���^�aȹ��^K�y %�ʾ�/�E�7Ix뵩H��Ik������vYz����=�jP��_��ѣ���H�寳�5&\�X�,���D�7<H��z8f���؇k�FA�m��#L�zI"�R�iGi�2}�g�����R��j���d�`������XV7�à!/Mpa|A2��,�m�Z�;�Cc�����~�y��\���Q��ķ�@���}ɽ�P�~�}�s��e~��Fn���U�z�9�`�ck�?q�AYs�3��Y���N諱�$Ȏ�|��	����Xw��ϱ.�k�>i�W%&.R�� �H�*��&O~�2"
!+�
4-������CD��{ V[S�(×�%��Ț]|כVίb8�L��j��I����� �q������~ÿ�r��c*�>�h���W�ƢaʮOƜ^�?|ϐ�ćGy;K[�,\��z{�%�94F�r#x^s�����=tl%e	�⇤G��b�z�1v�ˤ��MZ;H���&���b���5�I�']�Q��H7��m��$
K�]DN��pX��n^�uC�UH�����0U�@���� lX�'���vb	�Ls����AV���ȒV���w��_)/m��j�Di�'�{�r�|�X�[����|�^G_�pJ��R�ږZך\��Gdo��#)P��S�㔩�<�K(�U�,��w����3���	�������'�=�CF!P*�����t]ĳ;����A�*EDԁ�����Q��Z�2'�QN򷾧�>����pe-����9��^+n�,a���F5M��s�+�h�ʥ�8�@����	���δ�5R!FW�.���qZ�[x��r�Hk<�z�~�`��Ԅ�o�H$+C��B'|$�]�N٭�� �g�D�%t����Hތ��^��b�U� S�s��;��^����W��¿��'dy�xjJD������\�ZF��.�=��)����v׷�Գ���������{q2'1�?�"���G\��qǙ�e���5�R�r>_|h�f�[�eLQ��^��WB+ū���Gﵢ��J�C��R��U�[Q�X8���c]�0�x�u�i��W�I��?ȕ3M���0T���^<�{�n������EQ�`?I�|4pm^��R�OK��~�F:ԩP}���9�q��Y����i��,2/4�,q�M�U�Kd���q,�g%_^N���J9��tB�4=�2����CR�f���H��ś�N�a-� {���3�OZ8#�t_z!��r������!����l�0X{�HS$����@ʯ�{F�c�r��䜲+�����Z$Z�?l#��h��>���K���8�Ӵ;�e��Ԋ[
8�
LaP���F�^�ԮšQ9*)}�7�P�V�E��k$b���@c���rY ��x.���F�"�@2���Y�L��{�$��<�"��:9�D
�lv]�+�0�H"�*�1Su)�QT��d���Cm��㋐?�Ńi�� �F��&��#��o���*5ɻ.ǖNS>h�+:�f�'��3�HqC+,0�UZq�/�gN�Ⲹ��|��4#ِ�G2^���d��c�*c����b臻,�3�N�1�ϥ��@V}���ۍE�E@�}Ƈ��eW�̹^\v9��
	�^6\��'P�`��6�"j~VFBp�G�x۫+ʗ�=��952�ol�ܱo7,�ߘ�U|icn.JA'@�V������c�on�{�Q�R0O����O �̈��p���j[�	������	��W���k�|o7�&��v�*�3l�l��\�_-��un�p\��qV_xd��B��&�Tʡ�ܟ����IS����}������վ#��D	6>�V
�^>�ރ2���X�h"%��AZC�d�@P�N�	��3���8�A��=�K���5��R�6��Su��K�4�GP�j=h����ݒ����̪�P�@�k+�6�ut�i=�����,T�}�]��W�wqiQ��'07�W����=��ʑ�ч4����G~�i�d��?VW�m�W�8<������*S׎����F�q��H:�c�[k*7f�=c�}�ngu*Kb3�$eͩ��M)�m�Ɓn��x]��9E�T�m���������>�P����T6>�B�M�����]��(o��`s�	�j�]ƀUcE��w��mE&�Y�m��!�K1t�DR����%��!�u��PW������D��w'��c�4h=�C-���9>�{�m��b�u?�K�ve�OlH=a�;B�imGÞ�g�:��.MJ
s:!s0v7�+��\G��ج��g���7U2�2KAcm�E!t���5*��hH�f�\H%�)-1�2�%��p�xcQ,��+6X��j��$��M��;il��IQ�:��w������sZ��f�b��>�P5:?�s�p�]ʄ�)f�$b�2�1��٪�2�*��p�h����{�"�:0�@+���?L��1[2�ꀓ
jF��v�FU�ؒ1M��2�L��a3!9 �㚛�h�t��x�L�\Xa\Ub�k-�P�x.k���lFb�V7t�ӱ`���ᫌ-g�RnC]5��˷��r�9�l�g@��<�^t�V�m��ϛ��Rt���R�T_��
MƁ�K/d��E���T<�T�PQTS�♉�y_�+�`�y#�G��jY��?R`�9x�� ��L�����=X<���6�f���}y��ԥ�O���r3����fa�K�I�v+���q�^���敲���o�5�A�Y��p�]�ړ� �o\���uT;_�Uu�KCN����S���5[��
����r��huH�  ��P���Pm��w�%'�d�][+M�隙�)�g6j9�+��KX�Q^)���a2z��9wϤ ��m��ڽ&i�L����)�wF	�	l2MN��^ t)����yץzN���_m̍C��ٚ2��tX��}s���1��M/��w���W�I��*G��l�7G��[�P�A��nN�1�7�%�*a/�����@���м��1��!��':���	s��։+U��*鏬�yD87����BѰ��t+<�2#���+u�?}U~����e�3���pՎ4&J~�}��6�c�Nn�]�0��ɷ��ӊ��"
 _�����ܸ��>���`2�Q���PiC:�'����-��|��:��+�D�#~��4Y8�S ��ʷJ0��Ey,k�0��K�z�x'�N����_��s]�@�]����M�L�1{�	���(ӆ�e}���k2}�*�K������*N�ސ�+m��!yM�3��E��<m����GN�x��ȴErӮ<��.��_�����8'd���+�D�R��S;��Vf�b{��<������{5;ݝ�U�!��n��=��������s�l]��ME.|;.��'�e:�@#�u^T1N�f�|��0�s��ǻf��"_��G�fH,�}lM.�3��7ʵY���0r�qJW�ߚx[+�*�|E���u7}��!m5���r�
��^��=�u}+�#Vw�C@3�j�#���^Zdt	&I=̭KK�9l�T�U7���0*:�;�|v�}c���5U%���u/~{�a�pQ�3�=�i��Q�+ ��y�L(y��-Uu���sS���Î������J:Ճ������'���vWo�&P���A�]���C�攣���@_���wn�\5?��@b��!G
��*�δ���s�&n'�z�.@��k����Ⱦ��k�G�w���G�m�T�U��y�ov��3k1��P�ϲM�r򀆮�:�9�CV9�<��A�I�(�@z�Q��I��a築c�&mף�EZ���0����Z>!��W��UaO>��p���k �S?O��^�s���{R��D!�QE���ݛ��rb3�z�'�TX<�_�W��і���%f��}]f/��P�=�V1�~䄺��ijm@���J������|V3�m�M�9"���9�����ׁB=h4e�\�G1*_Z���Psv@�3�J*�m���<Wl}od����qR�&��"��(�|�\v�V-�* ��q�gߨ�P�"�{^i�(�ʾ�&��!yj{\9���{-��y�JX;���8�~-��'9<*dj]TN�%q�Ђ6 �/N��x��z�����b���b=g2�/-����
��ϫ�|!�`��G:\>�y�	��&)����yć�j)��rӆ7 ��Jn��96oM��h|���1eD�`c�*�d���6DSo�cV�1Sl�A��/��p��W�<�gq�"c�0�@�c0��z����1`-ZQ����y{�K̘�݂bZhs�u���S�I��s~�`��������x���z����=�۱�j���������fw�s�ȅ*���}2P�4��03��tb�/�o[� �Ɇ$����ǳ'e��Q,�5���LJ�}h�f����q�����=F��ţ�2ڲ��O��q�bun��ZZ�)sS�g��6��ׯ��>a�?����w8��5Kwc���}��;��3&��I�i��G�婒]��zrȗ����\�n`�*�T1�����f�n�	��io����^���嵔�~�?.�t��f�).ݎ�Aje�~�lk!^��2��b�[����Hos��xd,��@"�Ue�w<�]�9�)���	�n���I��	�E`,0e���P�u�2���a\�e/Y_ҒxQ�+��A�D"dU�qQЭz'�jg�M9 �64�H�o:W
�"e�'�u�n+G������i�b�y:���qqXY���~�����6�5��'T�Gm ��d�̶�h�$�T�u�W����-�[Y�C�h�p[oޣ� 3��II#1壓7��u_��U
q�C��Н/p��D��55�(#��� ������ҙ*��H��̓S42���в�!�%�.LH5�B!�3ǭ1�y4K􂨴mDrk2sR@ڞQc6�#a���=��V�vT[;�ȁ/����3 ��t��e���ĦP�PJ0�lµ��WS�9��B>~v��૙zq7,���*�{��K��IC�%���Ü�{��
 q�V�o�S�X���4S3�O."c,iO���K���7�"�g���GȰ$��Jb.�}Eh��[���<�>�z��}6MTۨ��s_A����R0	|0�Ly��8)�C̪nFa�[a��=3�x�Te�5�5S Z����4�_@��J��#� �Q�1KX}�,���n�F<*p{�l�_�q���k`v-e�����IY&�I̬m���p��?�A7Ģ��4ec��o��3�|y;��|��v����UmŪ!�5�҃�ejZ���%e���E?�,Jl�hC4!�DEE�7e?1��D�I���V��,��.��p�l�A��y�e%NSo9�Tv�&�+W<#��^�
i� Y$cϕ�nQ�ț��Q*�s*1�E��;����fx|����-2��+�їH���@�(��N!y��Q!{O�0���y�{u�E��G�,Z_���9�qa�1V�t��JN'ϩ��ݓl�
�y�rV�EI�:KT�$uq-@�#����p� +J�1�E��� �3�'� ����p9L&;�'��_��|0���$g��à�n9g�	&V�Ť�g&��u��H�XO>h"����ǦX!��o9�'���EDg�{�I�E�^ɧ� �n�IyJo ��W�xG�a��/�(F�Us�&n�ƞ����ە�Us�& ��V�\�����"�Jn\�K���VuN��Y��a�`�Uz<J�i�{�I��_7�*�8�f9�
���2��s1K5�Iٷ�1!u�?8�H6���U�i%���ca�U�O쇸*ܱ��:I|\���h6�-��w�m;�m�6��k�P��$s����i��n�VŶ��*EC�N��>�
��P%Ĵ�B�*I}%�̣�P��7�>�kr����k��&�f�&�ED_��	���\x����䱄��s꯿�]>�t����إozh���5i
�m�v��&����;q�&mx �b����C�<&ԡ�@���ީ��KAl�_�J�9�Ţ��� M�Z�s��50�9� v4�Gfk�W];ݦ�ܸ<$,��8�-�����~c�^:��''�K��sj*�r�/@_�2�2�4����߲��;_H�;�V?�L�C�RI"���|#%�4� �lP. �#� 	��a�r���|�1b`=Z8/>+'C�ܠ��='����7�F�G��F�U>k雍9�O=�X�m�B�y[�ɮ��mB���
�^�gn�!��XR0��/���2�P<.�^�S���Fz�_�R��hF�T���X����!
���|
Z��pM6�L_Ì���� &w⃎�
Y4"}r�����7�fc������w���x\2B�
%0��kiH��h����ϑ 61N������i�Z??X�ɯa���q�=f���u��I��r?���vm	zP&a���4��*k���;o�����k�4�h�����(%>�����F�7��}����,.�(��N��=��I�ɣG�ku�I��߻t�� `����[H� ���VZ{�R��� 	�6�O(��5�$rvh�0>`��K�������p!�z�M +x�D����E����ةRI #��M�H\��G͕1"t�&���G9��'��QnG�#�I�T�d
����Q����2V��T���G��7udU�v1䑵,�C������.����+i�[9�7S�ת�i}P(��s�?NU-?XI �M8�,Mk��#��� M/����=�1Z�8��7D���g#�>��ڣ�;�����N�)��e��nF��CUi����U	i�		8�) g�&s����V~��5��ޚ+��3S�8̢L�,X�6���F�V�^�|G?���"�|,wB�|��1v��[�� > ,���>�d���bE4����	�r4>w-�Gk��D�م�t��p�gok5���k7,�Y �����EX��z�d'�3*E]��ͭ��C�����_������U׹�kN:�"�3�	D|�o�*]�Ǽjb���/8���M5ra��#GSjq�2+����<�ỿ\T=J���>-��e�B��e( ���=}M��*��_2w��������K��.��G6���	1��[l`N9_X2�����A8��\<(��P�^T�_�R�X�G)�����mU$���ȁ�o�ϼyn�X��s&" k �葭b��p/�4Q��"���H�@�n���vס1�)ۡO ��0*��`�v�:�,<�`��E���TC���PM�g��[�u�}c��3~G��� |,r���v��y")n̴B�y.�U=�<�?u��#NG�K�N`��-=�]j�x�ړ��wZ��nH1��ˋ��C"_ƕ ���E�l��l5���"��L��<n�v0"���Rm}�E��/�23�9�2U?�Ak��

b��4�K&�m���\��e;�2�%q���w{w�w
��G&.�lŻJۇ�&��ڳ�?�S����)qKiJ-�8b���Li�vO	[���ŏ~L��=) L��Ҙ\4l:��t�@{�q����0�l��dOUb��WĂ0ɉEI�h��ܽ�S�bld�Ypb�*b廾���C���Ṕ��&�Nn��*f2"ﲔ$:�Hgc�W�����mū��)<���a����z����y�s�dI�O9S�����1���kNZ��͕�ma� �PrJ¯Q�M
����]%r�!���u�YC?���6�x_1KD9��|���=
b��5������쁱5$у�f��$�~��iU.�		��c�k��it�w�9����� �$��Y����X-\U��"):~`�9�7�S�d匼$�h���/_;x��/E�/��J�P�	�s�F~cR��8�V��3��	�Ȟ(4�hԻC�67�7o&O��*�a�E"��ϼ2J��w���_4��-�׶Q��V�;4�!��2��6��Ál2�_��M��P��]�T/��:�
.�>��J"�Gb��;3 ��)>tL�!N˥!�z�UjQ�ݬ��T<�ZZ�~�A�@gF�̖{js@�Ng�1�ux���a�{N���]�e\"V�P
�<܍%�������҇6YgҔ���Rbq�R]z����	AjT$'6:bUk]lw�8�F�B oPs��>�Z&0M|'x�	 ��&�D�A�w8����Lk[	4S� ��zD�!~aA��ǲ։��m9�U�L4�cʔ׬�W��1}�ߦ'R�^Ht)������~b��d�F�F/�����.b��G
d��	���
$���T?�pC5�����(52"t�9GI-W*���� Zz�T�t��sl�A�V�މ�t���h�&�A�:��Z����ZO:i����u�����"����t�~r��*b5����f�V�\�j�VX�*?��ZnJ���ݵ����ѧ�J��������q?��)q��JZ���$���`E��w�1��ة ��zҩ��z&�p?�G��M$��Z�ϡ�v��bh�����@f�Ե��h�_��b����uZ������ZԍHX�!�r�1���%tR��3%��#Q�mT5x�6���]S�<�~�F�I��-㗤=s,��N��>�lT��r-�~jJ^9�`D�ҫ>�{Z?�ǋ1��lٺ��
p\t^�unE�'�7*Ab+hq�N�6�o;�7c ��#̋[+��[
��ա���Y��s�_�g�k�(}e5��1;���T�π �YW�x�*�z������$�Y��r�M����!(
�xd.����x��R��,�U���t"��Î�J�Q�>1Cp^N����S�N �qk;���6��dW�<�����:�x
�]_n�nO�n�RCE���Eex����p���9���Jc�����6��2oH�Y���ߚ�G���cC���b9�`-�1��JΔ�|�`��9Rr]�NJkܢ>;hFMh���p�v3g��1A��Y��eg*����+'��ԡ����7McqM�d�Ӏ�Y��VE*;��g�J�9 �7�u%����c����+��H��w��H�~KhWh*\�Xy-^�Nƚ��a���Ak�S\��p2,�fU���[>�g(@��PZTv0�r���/�Q61�5P�͚����\>� v�?�Ck���X$#�h�N�r'���<��A_#yD�JfQ�F�����5�*��1�8쨷�4��lA�q�&���<������0�:��n���G��
$�I���S�'ƙ�6��5b�-I��	���m�'�e�����59�\NY͹IӒ�s=*�y�G�:27�J0dҚ��-��|7��]eW��W�q�����L�c��"|�)}s���8��ZB�7���&
�X=��  [u|{�Gt�����$P�!/2T�"��S����>.C���@~9�� �ˉ��7	Z�Y�	C��	n��݋��ݽRp~}v������Vo|m��f6)��,,�*x"5��K��Kz�l���op[���P'������ț,���>v��E1����%����D���ѫ�W�U�/0�퇿\�a�����z�q�wFo�˯x2�p��#.�sV�5:�>��h�k��%�s���-�&cw�Wml��$�gi�K +��!-�r(iGo}� ��I.C�:HQaֳfvV##�$�@�Z �.��b��,Y��غw�:��}����[a_�k%Ewn�$t�u����:Tq�W�,]bHe�z��C��(�T�Ֆ���c;_zR^�$mH�k��-���3k�-%��G���n#���C�q��c`Ur�X���}K�`������|�)3_r��U�O�H���e=Rzv�1:,% P��`Ǔ o�y����W���efبṳw�:oX����Ei%� �&^ꔁO��I��x�8D��3ivk�=J�J�Beo�I(�霕Ȣ<-R��fYVVu<���=�&��n�J��$O�����t�r����7�X�g�Q�ۘ2<S�#����PL�n�_��A��Xʍ��y����[�;+��x	���Ԯ�S	�Q�8��ʶv�٧��E��6FA��Ja}��hz��@��H{h����ۺ�<0̙�N���T���8Ǭ<N��)�1�dk��_>E�ј}j� �I���O�.�m"������(Jo��Y�@���ˊ����	���AJ�0������|a�͍�YJ�qz��z�
QO��h�0���R��J?i5�}E_7*�_3#�sjP�c�r�U��E4��P	��U�=֥�k�������X��N2�����2�
�Z)~e����J�R?�T$��LÏtI������`�͍�
���uzKz�|T�»���y��x��F��[�'B���(W	�FD�C7|d|��ۦ�6�8"U���A�f�ި�UZ�(Ig��xh��yM�{��)��i�O[ϋ����L��z>9�ѿP�.qd��O�p�âO�NA9ܣ:[2�����ْ�x=TQ[ٟ��Zo]��(&�/�U���ϣ&���b��k�ЈcDM�� �O��Y������>>6	
��C"41d�Zmv�Nh�c�k�ٺ�P�(O�X��v'�i�
��l>D?�۾p�()W=�;-|c���%ExJu�E̠���	͂����ny�J�F������k���LX0�*���S���p���(�U�t�L�+U����vf>&T���Gz�K-���X�.ۋ�6ǅKe�iCJ;\E'�tL/A�r���ʞ�M��M���� �q~�j�k�n�����n������[!��eU4��&!;~S�Í�:�\��������	J�l���轀�jF|�����9�2�6}GGY�� ��uZ8D�w�U@�%hNW������(�3fi��J��L�=/��Q�w�6�qp��|p�o=�2R �T����6��x��un���tW����G�r��:��DO{g� �D#󠫜��8�)� �L\�C�a?ue��
4ѹ����RX��,�����:��-��M��a�I�Аl�u&w{�����X�w��"��!��Jg��5�H�	x|���.�^Rp�3�[#����Fj'd�ר۷�m������8��2�z6.	N^�+�[���9���)�Aiamx�T��0p�w�!O{�m)Jm���Z�y�n�r���+�~���/j��c�^�=[�8��b|?I�����]��1�S��ͨ�����ɝ�72�
�D�P,��&���`P}� W��)�+-Ev����A��ePX���hW�5�N�Zȯ��b�9�	��{���K��P���>�d�<��{]]y����HxG"�m�	����s@b�BT�k.M���ܮ��s�ɴp�=g�/�����
�8��(�5ݶA����V�k�ug�h2ɉ���}[�x�U����Ӥ�-��~6+i���i�Y�
�^�n��~�t��E�OAG��F���G��nn~�} :�5��Gٻ�r��a~2�q_f�����ЛLB�Z�f�Cޜ��7��ޢ�OrvXm������~\dM�Ħ9]Dc5�-�Ef�}��
�R�vn��~�������l�W)8@��j~�u�3�ȹT%�@D��m톀�}��A&<�2�)�\R���W��U_ej�E�>��U�o3��X�k�j�bG��Kօ:W�Z:ￍ�n�2�)}�J+W!�X*�����ɂ"E��k��S�Oί��tc��j�ʻm�]���E�{hTr�l�2Qa/t��G�r5&��NeЧ�lI�F��7�*v��x�eg���ĖP����E�G�{�B�W둒��I,.ng+?Ҳ"�dڒ6��5�Y5q�C��
ZĂ/D�!������~�M��ĴÐ�b=X eOimh����7k����7�{}>�߼�Jaz?��^c"R��}��{����۠T�/5��rg G��������?�UZc����ŵ䗴$�����>����hR�3&�0�-W�5'/�?.�!���z���S��L�@%:}�2g(�U�����)0�;��Cn�g�HNL����P��4m�0�{��r�J�C�(+�����$�Y�15~_na�D	i�D}z��I�9X
�wj��޲��F�,�G����}�u0��SX���f� ���[�E���Ts���ҋD���uտ��O��j>�7�d�b[�4��@���V*��"�zkg�f����|�
�`AE����ڂ�
���؉d�/+ki���x��	��iO�,Pm����O���m�{����2�b��or�Q��e���)4�[�A:)'^�NY����<i�#�n�*?GR�ֲ��W4�c��J�J%�М�hu��q[ܳЍ=9J<I�&� �!Ĵ�B��gr?��������h�,SzO�O��	�NZ��d"TqA-���p�a�x����Q?U9�/�#o�6�ؚ��),v��J�\�����`+�/��~@�4�&���Z3.����P!	���W�Z�EGV���B�r�~H����CS����Z��w
�7��~��c�*e��ZX9ɺWY��ӽ?NuJt�v��ه�R�y��Kp�6���ܚ
&�d��5��!��H�n�pr�e��ٓ�L	b�7wP�+TM�P�Ѵ�4)�e�$��M��^��/l~�⁡�d1���R �J3�����O��?��Vo��b�n�%�n�ˉxŎ�\N3�� �~��U�d����d�s�-U:j���� <.�t��������څ�����wV�F>�̽:/��+i'8@Y`̋_L����r1�x�CG�rK(�dѩ���g�}�8�-�Va_i�>JСSn�D�AS?��}����HwU�jМ��=�K�����91`˓�6���Yr�;�N��^w��-\�e��d^�oE�YA��&�Ϫ����=�j�����s˄��2�`�TmqC���W�N�P�Y�51��N�kt��)�g��t�!kj8A�N�XP�.�n�З�W' ����&��� ��P��.4�yн~�����fbm���K(y��Y��2��-#����� ��<����s�s��/�ʵ����2s�T�>��
��E?$���KL�\R^z��a��m\�F1K���̬h�A=��K�M��O�#�R��{�bV��l�&�� ����Q�s���H�U�ˤƢ�~��;��G�{p�|��;����Kֽ4��W�OѶ��m�����=ֶ��S�{EP�	*Jh���۾�9�X �����>��]7��;V��AzkB���8�i�
����Yԥ��zd������;m t�����f���
D�\4��I2̣�����~�P��mS��� �����{��y��ک�$7�Qs2l�Y/B��<�hb���{Ns:%vݚS��%p��Q�@ ��'8��|�����4�H}��R�Z�?��}=6��6�_:s�y}'��<I�w���L�����15-`�KƐ'�ޤ]{0�@?��KM���VFԁ�vG`���8�kN�t��s��p%���/=Q�'&)�2�W�֟r�?�lTa1E�
�b�k�G���s;���ؾ����0+������u":f~AV{2��FGg��\)~�w�7���@� ���~��J����'�\
�8�Ԁ?���p�,C��h�`�w��32��m���d1zw&���P���F��:���jflSxЇ/�lGC��T�q����zjV�l�D��3x��$4����eMc��:S5�ɅT�4���p�Kā3L�RgY�1���4r	q�h�I`1tc��$�ۺ���m���MA*��-�����R�Œ���L�`�Z�e�$�)7j�t�o�-���c��5H���d|۬���Fw��a���̻7������K���a�|~IB���	z`u,HN����mlx����}�<��'�j%fb�"�0���<}��s���L�n� r�|�əO���e���%�G�����8w��3���t��{ƕ�d�(�e�fM6��U!'�
����"���,��p�@M��"2��4�(}=k!	 L9��Εϩ|����-w��b��Ћ�*κ"!q����$�P����s�Yі�G����8�8/Y�/��_7����F^$xP����6loQ��X���sZ�e��M%K��!A�Yݪq�����X�����R��C2�/��8i��+!2�>� ��n�����|=�l���2W6r��6��/�̒*��U��nLd�:>$�ٕ�K����>D��(oK�A�x��<�Zռ	���}�4��oMN*��˺��&v$�҃�8��INyn�^Z�ص���R�b�KTC<1�$�՝�gȭ� �K�%F+(�t�Z�6�C6%�쉂���?Fa�_���GS|8�5ٴJV���va�흣n+wX�ӵ�>p����g�ؗ�$�Jk3�o�<ˑ|�Xa|�'�#r����ڲ�Y�KJ�C֏�M�1h�ŕ��	W��J��θ.��^�����`�
��0&E��Ga]����<�쌾4|���Es
�$6ˑ�Z�-zǽ�TKCzu�~~�|����n����oհ�GS��IF�;���+H��E�.�K��Y�+�G���8��-��xД�ލ�U�1�Ǧ"u)���U�٪44 �99/ V�Ӱ/}�ܳ8G�������ceZr�aGl�P�w{�x/z�"���a^㬃	���"'�_�dx͟���ab�$�pcʁJ3�&����5w�,��r�RyI��N�oWՙ�� ę����&ۮ��Og�.G����D����|=��Q̦������,�>k�;���k���Sh ��2��Ǜ����r��u�;r���M4�r��!y?D�l��l������I%,��n�r_����tT�ч'EB��v�@|��+�H�I���Eb�5%��0�c�U&.�"�}�zֆ�FL��N�,�g��V�V�{.9���)
W8ħ�9O���w	�G	�2u���s~�+5����Y1x9쎨��^�c%{�(Ǳ�h�~�<�D|4~a~�g�^7�r�70e�����BG�Ç;,;�6CI�͆��xP��׏v�d�]��e�,�F�o��_��&H�R�m�C9�ir��o6���؎Q�M���f�+v��aY�0
�/[;Z^ao?��b໦�E��>C�d���v�ɇ�Cl62��׍3
/�?^\Y�7�ո||Åsm=���J�q���$XC-��$7������������g`���p��Ì/25��`9 �Z�eb��pfM/ ŔdjD�y^%�����U}��w���:S�;��(��\�+���h�+A�Ѭ�f�|.�ʇ����Y���;.H3�{Ʌ�'�^<���j�쩿����'�p�y��c����2Ղ�i��|���T�#$68z�Q!u��0��A�6A�%AW�N=���>��,����J؄M�tkl��C�5���ק&�o��W��qC�P>�TC��K��^���ی<��8d�a�!���/��q֩z�Z��g��k���F���5Ɗ3e<�\'��p s;�ex�#�d�ч�?���P�#�x���A�IN�2�M��׈��E�ׯ���,�U�Η�ж���*��_Yg��F�?6e�s�����e�5lS�5��BPƍ��N`y:O�#~�7H�I��m�F�n���N�M��v�b��^��i��xR��zC��y��+�U!��mH�_r�����,k� Vb���>�\�u�M��Ձ8�~�4�}pd2$xA��QŴn>_ʼ
e�G,�3�h��s���qQ�� qu�`d���%�[�eBd��r��
]����F!]�Q��^���F�[U���$4]��	�и9e��ÿNFZx�m��U]((�]�`�l��v��z�u<�#�5HJ����ᇙ�B�MmJ2�%@�q��g&qpr�]�E��̥���6���[�Z��_�
�m���������6��XT M䁉SH��j���z+b<�3>�4!�-�m�l�b�~�b%V;�Z�L�w�KF�۳K�U�M/�pB,ER�BRp(��a3�����$釃2Bg����ա���S�#zz;a���r�L1�se^Ur����w�Rw���ҮJ�>>Ŋ���I\DP+��O'��I1��D-���yaF�@D �{T��m~� ��F��lD<dh������ݶ��,�~]����8Ό��������1(�dmY�Z*Щ�c��p��MO�}�U�L��Kqlg�S��df�M=�m��������d}�9R�+H#��*�Z�8aw�D������a<�k�8�<���@����zc:�p��R�ǡQ�����D�:��dw����á�)2��w�l����N�?"�R;��uL��!
H�X������^Ń��	\|e�f��y�\O6�L i~iI���w�f]�5Y}P�y��C���v�:w��[�2����#�=�eO
.��:�]ǒ�H�� *���	%]ۿ�V�-�����`��2CiB�b!nX�ue�a%����� u�+��b=��]s�
��}��`��C��h;�!p��� � ���������A��G��wK1�Q z�����rH��ط�'�r���?Ŵ�?t�
�[��=>E��7�Fu�a<�	zj��
�=�����u0��KܑD��;������앷L$;��a�� ƿ�%�r�@ݛo$�0�T��HZҐ�g���ʙK�)���~:�,J�א������L@���zt.$\H�N�M&��������T�Y�!s9=�H��.y?O�p��W��b2�B^2��?��_4�/f�U	mG��1����EiB ��:�������F�1�j��?��"��V.rP$.j�W��,�� ����݄����o1��U��*tT�l���\�X4T�O�b�����kKܯe�{6�Y$PS�ф�N�=$�~�V��D4#���m.;�@�7B[Lˇ��`�6���NȎ�O�" ѯ��@�L��;�yZ�k���N�>�11��$n<@p������!6V��qD@��=K�m%j㰭��k�:Sa��
�=	��-q-O1��Ú��?X���/fƬ�8{E"���3)��Z��N����a�ԗ���~qAIˋ�L+X>(�\'�ح��^�͞��x���	^1C�Ϗ� �Ij+�3��;����Q�	�]��<KD�혠2e�e�P3�5�4Cf���Ѳ�N��3�:s�
ͦX-#�ʷ�R��s��-E�{ė��>�����+������ޯXɦ�.)C 	�0Y�~I�,�U�7��u�t���pc���=�1���^���Dy��)l���T��|L�Z
�	�e^? �=k=��i^�ƪE6�C�@kc���]�w��Ei�]ێ�#��{�ϡ�����E��l}�����q�8H�������2~��E��Y�	��|hLe�z�a�:]>||v�P��&I!�ƫ~H�<���ħc����KlCKI��h%02�|��!S��W���9��X#,�杹�AJ��}п�t�E��|"C�]kw�g�y�0]��h�h�/#t>v�AEb�"��r�|���
V��n*PpF	����$?FG|^,�����K.�%,l��e�A�«4�Z't��_�o��ô�A��1�Y�� '��l�V*)�d}��������u,�4&f��D�����kn֩��x���<���U:�tw�!�4�b �e7��}�G��o�X�v�z�>"�)�m��X/��R�����L�;�Z��WE��)�90���v�G��?k�~1�/��
�4�R�g_�p��
�ٽ)	�����r`�K�	��5O)i:�Ț�4W�Fs�>���i������|˴�e�W~�;l;!Yڭ�l4Jl!%�}��+��$�*�)P�9�߽��Q�i�Ao�I��V�O��p4 9�%f�����ѫ� ;0������Q"��]�[n����m�:;'Z(�3��q����Q�k��j�}�٨9�����EG|�6"7���&:��1²!����p�&�p�Jxn�gK��?6�8�=�"D!������B(q'X"GVo[�o�A�z�J�Z�ʲشP�oCR�"L(^�I�r%6YDSa��e�=���+T��R\��7��Z�D+���nMj�f4��2�q<}����؃Z����O=�]�f<�/x���I^�.%T@B��<����D�!�RW���0?[��ʗJ
�tG�X��^9��bƪ�o�l����-�����ߞ˒�j���N9����NHP���"@��~��K�,Wu���V'=�@$ڨ(�d(��p�<�C[g'��ʷ�#	p|��a&6X2�J����V)�5�s�l���~���0���?�C���q�3? ��$+���&t��x���h�&|����&�`ۈٰ��8=3G+��k[�a>��خF��X����U)��h��T�B���YX�U��V ��5�p��.=.,U�y��>��]Мj��
��RF
�
o����M|�\�o�YO��7�%x�(�07f6�=�[WQF�_�F��O�}���A+�&D^��?������������v"C�]乆�n�*{����^0q�m�&�-�h�D�o��=��k�A@�\0'؁�eԺ4B���L����s���˪��2�j���q�}/<�Ո�A�3�*�ORy�J���u���s����?��Xျ��6%�3�5���r�4`%rH�% ���������Z
N�ӻ�$�����2�U��d�{o��y�e�^��=�!m��TCfF�� �0�N���L`i���1���P{?2(�<zu�M7z9;Z�iG5�k.�݀;�D�jƑԐ���R�W���������M��c�!�3�����^�uS~��܄���f�p��T�]��)�*�g�ˇ뺞�lɪjN�o2O
K;�8Mʠ;�|!��ʙ��II������7OZ�[|7Iq`�a�y�Oyny�s`��0?�l;b���֬R�q����9_1x�f��'
������U^5Drw!m�k�V����*hExse��TD��g�h8��5�h#�B7N̍.�O�@ V�b�HE\2.͒%�Ƭ������Z���]��#a��*��nJ(j�ͫX}���.�YC=�#�*Mj3�w������<+<�Mx�~�ϕ�eq�p4J1�O�8�YV{�~>/8�<r��C�)UW l9Ǎ��ꦽ�S��<N�6�_��0�PL|6�Ul�wT?}��� 媏$�����7�O��Z�Mz�bd�dK��8~�k�#���?<8�J/�||�U�]}�z��?v�yɖ����L�w�b�`��d�:��@I\��@xO�� jE�}e�^�	艄�ؙ��S�sOp?��@���h�m������!���m�LL��s�D��4L�^G����w����t��[�0K�D��pG]n4��&tyI8n�M؜69\�4
/��T��׀+@�Ñ�x��v�<�u�o�ZXh��	��%��~���rʆ=M^�_��ɿ��$��7)hkYbu�K���H[�/�@Ҝ��k�f���wȗ��{Z�uf�`�3�ve�@���!�=+
���hv�j��c�S���
�J���HDy�]��f�Nl�9�D�S�T,OMY���w
G��_�?�z��7'���-��LF�'�}@���E�����Ve��v���Vc�ZW�bòi s���,H���"D5Ti��p������6�\穜��k��,�pyx�_�pC,��KZ_.�����rg��<!��ޜJ�D>M�V�
�"�����0x�����3R�Fx���ዏkC;/� kӇf�֞p�?�RG,U��\sv8��f�}T�i�lQ�N��
|�#CvG�$��K%�l��$�M��8�ף�z�4]!�܏8���p�n)���5��{N9�PN��<m|C���[i}�n��e�S���m~M����tXUiU���R���F�P�c���	W��-�=O�/�Gp��[��SY+W�(���]y��c�|���D��ޙ��'�F���դ���u�۔>jn]D�W��]��z�1����7<e�¦u�UZ���u��R-&���-w�V	-z�%'�m<�z��02)q�Z���l�����)�� ���-�Ѽ����A˷�s���Gȇ7/��o��E���RM`A:�dz��q�RO`ƞr����w�8��4�Owe��W1!�d�p������_��~y��1*5��d�%���mұ�x��䗞��a�@��OZ!�*��7ʩ��H��8�h��t�m��%�\�G,QC	t\/�5N1?)e�e��c6o�VWߍ�!���B%y9"`c�	�e���%����SG*>ig7����I�"2�
��5�bv��]	���9�C�	N�<����I��
8�>�:�mx�{zRL���1�:I�qnٙ!�U\�J�'ѩ\�� �ծ�5��-WB��f�2L��
��_��&q^�22�_$LM�R��2:vy胼�i�W��
*7�y�r*��q�N�|e��"��F��|�7Y1�}S2U�1y�����:G��z ��fcq�\�,��u�"�&�A{����4
Ln�~�~$���(^a��R���B&0p-0����`���+��3/f�I9k��h��Π����p�
Ы>��"coh$��H��!^QA�_�����jM%�߀��j�7�o�gD`��&���gp�q����9M�;�M�1�*RN6�#��A;4)�*&kP��H�p�魻�n��X�kZ�`���OĒ��bдd��@t��U��^��I��3�-s��R�L���o�V_c䦬K "�k�+dR�}�x���6fR�� Ǧ���Q�ޫxt;�g�����/Ehڔ�T��9 g}
Q�,�JzڝR���4��x����o5 �V�p��@K�ߠ�ѳ݄�Roy'��*I�H�?�ٻ5�����a�&e�T;qe���s<9s}�::���=�B:W�b�PĄ�\�Q"oD�P�*��w��L@��24�8~����L{�F���o�P��c�@���Y�k��$n��7�`��	`M�xUV��>aYO��"��9wp�#prV�Z��~��&����I�͗��Ԑ�=�FX(Q��o��]v�����lSDʨ�<ք ��-F>�����Gc����`��>�IM�r�
��'�]--�B���b�4��[� �g�;V͵��<�����3�5���n�i}���N�W�O�����(t�x��{>f���!X B.	��{yۈ A���F�4��է���
�Y�c1�3��i�*>�P�o(��l|�ο�돹���#`OͿ�Y�?n����%vqr'@�����k�u��t	�P�����=������ڊ���h͜���0i���Z�����@du��Z�=�o����.
�R��p*��oH�^m�JnhQp����j�`�)X��W���{�^���t��T����e�sK�(U��O���x!���S"��� i��,B#��_}����R���!��(}G:�Ϸ��C�L	Q�!�����(��]V�v�?���ɑ����c`ޏ
�;�I�xY<5�!f��ȱъ� �ّ`kGd\�V���O*9��IV*�֔.�@������ͻ��9�uNl1���2�o��N�L�[��ɐ��|j�;�t�J�4[a�9 b���ό7�c�=�	���m���-ʻZ�m]�l��$��0EE����ܳ`E�r���d�:tS�~��P�CJiX=𑗜R�7*�J���[o��Hl��\�=�C�����Le,Ts�k/���\3�0ʬik�J"��*)%�}}h"˴:�Ǉ��0/�h��m`��K_I[����a�8Ab�i�����Nteh���'��ۗ�%d1��`Bp^������In5�q~�QsVh�4q�F�nc��p/����:�I�$I���=��`���Ǉ�w[r�/okx��2�2;^����-��o�b4�{�|��T�sMm��+�<3q�5�W,���o����LHnj
rw{�|�����g$��|Cݘ��2��x�g���q4wK�P��՚4g#@F�&�����W�v��*�:��D��#FÜV,�cN"�x��X-NgH�G�2�o����rC�تV�[Z�W�em�xv�G�	H�At�7	�UlMM񘝐cu��B��9f>���]�ۢ�{��y��]ضL�P��W<s3�@�"d ��N���RD��Ę����Ȑ�_�̧�WW|ce�Y�ML]�2J�#����%Re���{DO��{��٤�0���U����yt����%�q��g�����c�;��$cr�1T}dC��6<�1�@�S[��G���S�\�iU��D3.�}H�	W]V���fw}���� ��g�n`a���\��7�X�Y�sǡ���xa�{��+���ɴ�4�LC��x��r	��y�Bjg:׊@�©`�� ��>��q���̰���b���Y�9}�XA�Vn)D�~���&�FC�l a�1K����ʠC �~*��(��� ��;Yp/Q��8!BV5�1�~J�L]_/��E�M��o7�s�-�U��m�2��L�����PTy1^�PUr������O�:1��0u���:��<�h�e��%���5�S֎9qc!t������y�E�Bξdrb>-*�،^�ox�-����'qNos0Yj��ĉ���/�nT��X�!&.�5Bv?s���Jc�6�f�0�F0���א¶8�'�֙�gM`�搈��~m��?F�������j�H�^L���0��������<� �tő���K��	s��Dd�6c7��˵Wv�lɨ*�4YԆ��	��Yl��-��%�Z���SnFц��M%�j��0%,e�PTC����PO�^�d���ec���H�]c�^������ m�/����y(�A��Yxq�X4U>���Iw.�/Lʾq��P(~1i�3��Y��X�Z�M�?���
Ԛ��`�+�  �ٮ�ŮN,g���G��M9����9 �1��>-�Y�@��"�ȱ[��Ԧ���F��Ȣ��܈�m�w�q�����/�	���Y���7&��`�bv����2�ֈV($�"�i+G�d8I�ߞ\թ���Ls��It�3X0a�n6o�{[��<�#,�e��?�]�Ese=1Q�@���Wϣ7����h49G�bN~�s���~���$�QH�o�ݥ2����B>��
5W7N����x�P�̤׶�96��]�z�;�R��̰�*����;-[F�J�n��d���gO�g�)�a��Y��0��(���p�JHN�`;=�V�;fI�S������W\dl���xs�|W@JS;�����	d<��}Cq$[X�A��$IV=#^a���:|��!ⷐ�%�Rz�^iK���:�9�� .�@���랴�	�f�3�Ư��xF�	Ű��A�Fn*��K!� Vz�(��2�O�$=��kEC������2j�&?{��s�K��4XZl'�Е´3�B\�E���m���}��/V�I_`��!����x.CS!���U��k�:�Q�Sa���9�PO�H�&:������[��H4����|�)�������f)��N�Vs��/})�"s��َ�x�E!J�]�>��5��ݨ�T�8t�bUl��fF❦�U ��A@l/��Qr'+�^E؆O޲�M���P�� O�o�����.0=R��j��*5��
�.�O���ki�Ň��x�18��A*ºNQ/�3��%˨����4��V?瑷��n�|�,D���D��PS8ASD?�g!�.Kq�`�|s��T�TI�CH5�N�0̀>��� ?ֲ"���cu�q���g��n����)g�ޠ�q �$o�-Q���:e@�V#����de(w���lm���tJ�2��X+�ں|L\���եa.���g<M�(�s����� �U2J�Q��3��o4V���R5G�Y�FE��:�	�g� ��H]�\\�����!@����9˵v���EEj��z�gt���[����`�-B�qO�Mo�-�@�nOX"$ڕ�k�o!����О{c丙5s�	p>$�bC���$ͨ�ھ���zX"g5:�z�3Ҳ\�� ԣ��6Sڏb�늬�NCzZ�9���l�p����RB�B���+�P	iI?D>;���C � 	.[���u�l]zt��w��x1��I^zj����;��<��=�����sHE�K�\��_����5Fg*��$�B�{��a��,�U�ji���#0$��2��e�������9��	�έ����5��\�D�0�zm���{�gƹF�`�S�J�ݷ�Re{���?�oH��";�YL�I,�s�V�EB�+D�rr!��,��;����v	>�uv1-v�6B5)x�"��}���4j��8^����ӆ�K��W�;��u�F��0�Rc	�r�b�=uUG����9���������2�L<