��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��&���i} Ĳ?����D	m\;���k��o���W�c�$'�sĒ&�� ��Kt)��A9z=!� ͵r�hQ|�{�9G0�&��o����ų5�غ��6H�T��~��QOI����b�� ���k1�|^�fD yέ�L+�U
�����>�DKUf33i�^%�;G@-��y�A�XG�в�|�՝`��;�Zߟ�(��
���?2?�� f5��6T".�M�2�BG��D3Z��O ��ߑ=�x�`���O��
��-gv߾?����+;e�(׌�-�2�r� 6�@~;���	�h�^c׽�;�N�˵����Jh�y���<\*�^�՛�:��@wȰ���i��G���#���A���1
�6v��?��]4����s�&��xX/Vn�}���Jxm��H.�ЍMZ�6#���{[@W����K��x�8�zi���A�h�� ��6��-��P\���򉙫�xa3�=Ό*��D~��穡J�l/�|jlach|_x{�]�0)rR��^�)N����!�-���ϩ��	�X���
��C0-�7a�� �^М�:�l�8�,�oق�Vԧ���Z��!��-~�]:W9"K����e�g��O��˸{�5��{f;�a2��ڄ��:�_�'�=�W"��ZW �`v����gY9&�lH?n��ݍ	�7����#�'��F�x��bjp���6:K�7�D,ረ��2�˨.�����q���"���CVIԿ�F��WGT!p��#�\4L�w��+���s��Z�m[E�U��z�P:��l�wً������=Wc��y���y��O�-y�!"Q�~���_�G�T\�J"��2�޷�lBZ�RATr�lJ�[����Ѵ�Dp���4?sd�?L�Z���eXNE"����K�V��Ȫ�j8�?�O�4%̟Z��`L�7kr �F�|���&���2�ksŇ~�vRu��=5#����������-�L	��;����V�J3EY��)��R�#�9Ɏ�&1����zZr�p��s�vgВ�ҍa���睺q��[�A|�x������!�����NL��Qj����)I�޾E4e�r�d����XD�y�8?	� �6J��|��b�2��^�~��¶`�>Wa8�f으�{�zn�d�3y�g�@�=?�v�e�,���[�1J֛x�#���D:x?T���/̉5�#�U{����`n�2�ّ�ƤS��C����WQ�uUg;�!5*κ���$�ٽ�,�P"��h�A��U�1��|�c?���]otB����0����2r��F�ȊV;ތ+dzn�p~%~L��z�ҒK]�X���lַ�$&�a����Z�2HY�Y�i��Q���WV��yh�0�����D?�7���1�������4�|�ゖ��ZE���UPZ~�hS@�L�l�r"�Ѵ�(���=���Bz�r%ا���.��V\D/O�$mg�α�RF�'`HuV�ui�d��͹Ÿ�ő�ֿ\d5��@U~ e6u� <E�%b�)O���dc]3DM�.05�E�"���0}G����J��F��X�Vύ���C�R�2-��L뛶���$Ȫ��F�*[��2����Kb����*�	�T�[�A�넷��n���iKFl�ܴ�Cp��F�i��I���B�.�f�T����f��j�Vն��������t�����U�Sa.X`2z-V�ǯMwl!�d���7i�7��X�
����I?��O�:�q>�P�����쉪��K�{�Si-l��֎�i���a�Jj�L�:��OI�f:n���׈�����?P����1��$@����K��`Pc����P��'�����h��N��P�����%�4�-��|Rx��{��E��T�ߠ��w�i��l<��)��(��l6m�i͛e�R֗"V��=J"�Z��91���OA5d ��H/6�3�<�k�������&�����W������7te,	a�.^c*Kwn���
�bK5�q�u�(/�M�Rb�
"PL�j�G�=V���l��l��rCv<>����σV@d�5�@Ԑ%>�[�/+���O��넚�	/ꖥ�t�gK=��|������ƿ�~��6TT�^����-^���c�'�j�3��J�۳\�:jG�S1�;f���wL+��iD����_ڼv���*�F&�y�/�9�M���<�CƉ�L I���6��HD�f�}v�8��s�U�,���l��A�9@�6�.��n\��ͽ��b�r)�6��\�e�п�T�2�[(�c����"�}�!.�ܳ	��V2|Ů��,g]���n<P�N߶����}0�v �t�x��>��AUtjTn��%"��;�/'��5����D��� �/8�r	%#+�.rd �dD��e M���O��b�O�oU��?�t/�\^�;g�&����
����[3����a�O�\�'+�.�ё>�^�`�d�.���Lyو�2!g#�+�]����1W���|�)s�r:��������g����UI�=��*�5�i�ƥ[��'W)�d����9X��_MEҲt�0����s��!��.0~2^�Cnq<�R>r��w>���-�JBDM�l�Ud�h;���$f��*'{:��b���H�� �;|΍��O2s7���"�N��ž�c�����&�:)����	�m�A������NcF���s	0�����nlgR��v���"Y��U���"�\\+!�E@�
j�u���zW���'�f�V?��\��R������hFO�y�\`'[��.%G8�.-lC�I݆���$�O=\G�	�Hti)�
9����i��.�	�n�.Ƒ킶����xѤ2��q(� q%����(���ėi�q����h�)J��ޢ�]�w�{�5�g<�ls��tm�,|��	O#�j�ǩƤ�嶲V�����ϥL���@��L,�TG�lL����`�������~��E\����[�[���{]�Sg�Q ��z]��Oް�W͐��z#�O�N���AtA�@2�Vc�Z�c	�PWL���~�Թ5g۔d��
�����0ԥ�7ц�MdP~�;��Ӱx'�!��.Aۆ&�+��#n�?��<!J���S�t�r=�4
V[�7�[*8���BTף~)x0]:$��̞�$��R4�1���mom��{��8���/�J9[2Y��k�'G��#yw^����ӂ�i�r������&������b����I����{�J�0L��z�z��$$��P������`�5C4�����H�uX̯XW�4F�aѸJ*:�҂�K]A��I�
dr��U{��w�`��ϱ	��m�2�|}�����S��)SS�tܔŦ��W��n(�Bg.�=mȕf�%l�^���ˁ.ȑO�+�qgm|jU)oz|�n�ɦ�ߢ�dE�ƾ�#4��G��$���:EG¡���8fz�J�91âD��Co��-nmo�f��E�}�:9��3� �<�����*��OjH���>��5�EY4:�FX"�Α\ï���2�wh9���$���~�DF����>j�-���<��W~a���4!l!��́b��<�8����%[b�	:������0)l_�D�B�����gf�vk��f�����5		s����������Ӧp,ۚb��ȃ9����=�؁F
c .냹_�j	��R�K�O�U���P�5n_����y9�'dK�2�M��� �8��'��:EDO�\��"���9�o��)]��R�u�r%�԰,�"��x�C�\Eo��u�,���~�Y;Ҭ8�Z��^��X#�b#���m�OϠ����Ԫ�M�w`��%��M<�~a���եg�h<�=��g r���90��PՋq���A��s%l6g�ReJ�*�+�kf������7�?�����ֲ�#A-V.�8�H�Sv����5�|�{mߕ&��i,�)^�/�^���������)%��b����eo[,&�'^.~���a�ʟ������t�t!-��ߖ~�I�Q�E,4�c��?��I�H��������%fˎ)�{(�YH70��T��m`�[Q_�d�!$�g��T~_o�5���l[���4K�EuKa�R���m+AX���A�����l��=�G���FǮu��,�����Y;P�!�|�Dp6#c�k�,�#]���Jh���-�8Ag�"rmDv�d�EEt�m��|��}A��x�10x�B��HqVT��ʨ̐�T����[W�be������iR�n��A�q�B�u�R��:醳���K���E �C�>�B�M���k�5x�9`�\,�����G@z>Xf:K�)���cJפ�����k�?;���&����}�k����t}U���R��\�&%}u���trrӉ����C����U]��N�fU��D�ҽ�/�Q�����xV�0��)��Vtk&�I�:�_+� ��@&ht(�T�/��,5�1<{��ym�ˡ\U!��Y��[rO���k��E��7FV�V��چ���	j�'�(w ���b��Z��y��rA�;,e׬y������ֺ���_�DL ���*4�,��Y�C[��tnd����l��qOّ���	琓�7���F`�3�72���2���j%��!I��O,�r���K���Y�4�>�q�ė��9�Z{/���BYm��^(m�CuƂ���'�ρ�S�Z�L��W0_9��8"b&�w�ҕ���Uq%S{��s͡h��1c�+��L�p,�t��w������l������*º�
a���c�����X��l��Q�࠼�#%�?�A]Z���-�S{g#8�=J���to�T���ٿ�m�h_q-Vs�r����K���ͬ-��&,zRq��j����4tbc�u��:�Xr�I8V�I��z �b?�Sx�?ͮ���s��L��hr��?#F��[\L�M��RWk{O ���q���$�Y*H�;���T�[H���s C��AfyA�E`{<��B��$��dN�=��с�?�b�t��_���}o�c(�֍���''���,$��tѭBS���(�r��%3c�uOz�a�wP����*�9�dtu��c��gF�AgHM��x�seE�'��A�k���~�?��S-�a�>g��y���*y��c�ziڙ�R�%`Rq�8k�it���@�[/�0%�JF���歞/ȑ�τ汣����F���K��j"GQu�S@6N�7�����:؆6��@�U����4i��7X�][�3bFw�u6$0�VU�yfo�,x�΃\)ؔ��w+����㥓���Ï��  �����3�q�h���`l�'���&��	��g�#ܴ�vf��D��+��U��[:�Wz��@ �Iy�ÐZƆ��مPSl�p�OZ�&�g�zA7P�v�6�LO�K!�ڒ�ʚ���_ӛ�b�ef+�'�/�]TM}�˂-�y!פc~�;�����kL��Zj�����;X�b��&*�'�E�c��S�@�)@T\�՜F�x�k�<7s�iAS_��Մ�Z"J�T��$���h�d��SvQS;s�:؏t?�F�������6�Z3+\I�!�V��)_��q�< �+j7�)��#``�V8��XS�a	S����5H^��ew�����v�C���u�+�̰8:��,u���_�#��19'����-�L�������C0��J-�J������Ɏ8�0�#�sh�3!o�����eA�{D��ȳ7��-H�G��ʖ�\��Vw[7�op�Vx��J�:7*�y�6EuA��daF��C�b��,	�B���k�q�|4�U�B8]���8���\PȤ�f
���nP��6%���I��Y�-�L����	}%���j ����G堾/ߚ�{����1q%G(m� �'�~�%�s�czy8-��`�|�K�3�r-
�n=�]�H�� z�9��t=�ϥ�n�Ć,�mW�l��y����@�f�#f7���V�)<U�^.�g�Q�Z�$���_�M�>ZZ�e8o5�	?���j��'��m�{y�'�ׇ����5�(NbU��B�e����%�;Sl7*�]\���֪]u�1�\	��D�4jw����b.f����U
�����?���w�2�(�v遜�X��W ��궫�)"r��)ߤz��AM��5�2���\t�*<��]#��nd:��V�ws��@x�V[���!�m)9�b�YВ}��alNQ���������o��ۅB����Bj��&3�y8�T�bTCo�T�g�GY~#s�����G�M������ͯ�N����:�"{��+<iA�M������������5�~W��ə���cB7O���ą=�g3�L���$�E{��+V"��8��"�#�kI��E�cY�T�4���[}X2u`��)����"e�O�����`��H�Y�X�ç�f��j�L(��c�� y�?vu��tu�\��E5F�4Y[��Θ�o�/|�f��.�!B&����ch��"�kR�-�名$jp����)�5A���@'�a%r-�qw�\�1C�u���[~k�-�D1�H���w���X�K�J�ʐ]�Zl>
��{�Q>g�#�}ȶw���L~"K��u�,a�)�2I�R.�$�/�T�}���dN�b�ȌR�P���a�n��E��(���p#��W��PV�
��gg�d�Є6m���$W��:�o�x %��z�E��&N�b�=��kI�xQ�:A�U�&T9�&�Ŵ���kg��kEH8���_�J�Mf��:��K����+�oM���ǂ"�X4�1ɛG�'H1�	���$	d�n�y�AJ�.�J�J����"7�6�s���H�g�~�2fu�X&��8�L���H��`���G<��!�&y�T��B���W�k��}d �V��֓m/���[kew�W��탠4���·u[}�\rL�ةF��o�0�Ґ'QP��4�N��s�G�{�Z���o�)�e�8�2�=я���6�T��]wh���la.ܖ����>���w6�!��X(��^��5���|��LkO�ZȂgS��Z����q�u��~�p����h?�o|���i%\p7vB<��$P��k��d�	@��9J����
����c�=mDRA�����?�E��!+7�n�ڨ�;����pn��sZť��o�� y�6bkt;���زa� ��.�1n,��I��wu�D��	�����O��W��I猆\�",
�;��A�du����x��.���\\� 	��|F"�y�C��&��?Xm�B����r�2gt(���?o"9]QTq���O�y]0���[�����>\�%v�2 �?f��rm��|Ķ�Ě�H�3CZr̮�	��D!������2P�#Ҩ�[��A@��{��*#�5CM��B3�|�U����􏐞ė�%���:r�v��4+����uoH�\��'��=�����Eei���c�u3��Fi�|�f}-=Br~?K�\ː��:�x銝H~S���7?lS>��(�^}������1L�k�P�O�
���!��E[�	����p���E�jږ7] �Rd,h7��tg�1qUŗL/����;T�0��N��&��先e0���S����UȢ�I��e���.ҭ�W?*]���M5$����FL�z����zJ����hHgPɴ��P��g 2s�@V�����i!ZZ���WS݌V%Nß���Mom���9T> ��g�yռ	H�T��5��*�g*�s���ߢe�����s��~��Z
(S7�M��=`��n7s#qHn��C�|���O˕}��E��QF�Sq�:jo�>'"��k�H,cO��B�e���I�s<���?�O���c�"��(�/L@�T�S6�:	ع�1e�F�+N�=��_[�>\H��Id��f��S�ܼ��yhx�%� �R��Sg�7����.]��^�.�&<����T*�+��yj�2e0���*@*�/�R����ٮ�Q�b,r�Ӓ
�?��ըt{�ir�l�x��XiaY��ug�&E'Ǹ�\bS��0����ecӡ���Nh$���FK� yqp<u]h];n�U�B��c�Ѣ<z�$����j!4Uz�������?��E����jP�x�Q���;5qwٍ��7V���D��X�o��k��*�+;8���X�W�+Tu�Hs�S�����O����J���<���Auf,fA���h�"�޵��r�����^N>B5=�=��5p;��F1��,&rnd#����C�Y��%a3T9�h�o\���n���N��6��p>�����4�&��Q*�f1��v:�����}�]R-��|VO����� �5��!��]}�g���S����Wir0Y�ytA]���nAw�)��lx�Q�R(��_��UpG1�cr��kv媛�w�)�(���{�kV��E�ig	>갪?�)�*�s/Bٯ)��|M<��Z)�6:w�9]���og�dͥ6W?��M��v5���K$�pd^��t�Z���ą�+O�#;�ij��!C�2f�<w�u�XČ�#ys�\�-@�@B�*0�ر����d��9�t�۹D�gkT��!�|���Q�Ҡ �B�L��&CлB���<N'8Oi���ܞ �P�&+�e𯟏@_�:��8��Z�f�f�Źɨ_�r���$��Е��NCֿ"0`t|_�\�Y�/&_�᯦KZX�,:e7�CJ�Z�Թ����h� -/�m��)����g�q��q.Aq��cN�o������mkE����_�[#Cp;d"I
wL����zuHt�����=^WUeT�]}���u5�PҼ����h.�r��u�����xRjX{(k��ٟZ�6����u�hn��|�qr4���6��Ư	s8����dZ?�~��X����L)�L�L�HZ㠖�{���5���@���ݐ�8/wpf.���������W�%�ؗh`vV3�O!����n�I�h�����ϳ�����Qc�����(��f����ﴽL{�������q_��bKe�m�d�B�N:[A���ם=��甡�D'l��Gn���@<�΁���Ð��"0�Y�i<G�F����{h�����s�fآZV{�����`B5��Zq����-�G��ȶ�p�MR	���2�uU����`��+�@"�A$�}��}������ִ���W��H�L;[��#�R��ı� ��KZ���Y_�?r��C4��1��U�h�����y��{iİ1;p5��L�3_��-A{����YXF�O� ������0&��d��U��S��j+�\�ӣ�UN4N	�Л#�Ia7UIJT�����ll�!I�"8�ņ���R��K���m�0�����苗?�اj�K
-yY�~U[)�.<C�؊���i���
�h�wE0jO�M�O��FV����N���������ERh,�_�ƕ�@|�XBwM���ǫ2%"�R�x.,�h��Բ��Z�B�Μ݈-Z @��q��6B6g���f�qm�_v_C��(�8����.:^�=s��Kƌcy �Ȧh��.K����`�U�a��2���w� �3>����<G5,��� Na���N�T4$�5�xKiP[��Ik��!
WX��&���V���z=\Tj��%�eq��f��0,R����S;|�w'_�����Τ����?.�d��s���j���.���s���**N�� �4��!rK��E���~�wU��NPb�F�����J�ѕ�{
S�_H �:�k��-駊X�%}O�P3���[��3�W29:�$�݅^�r#Psc�D��>0���3Ѓ���'�M���
��5����)zG�bS��w��J1�M�^u����()oJk!F�-��_�(�����;Z���_ǎr��Pǒ4���1�; ĉ�9�qw��N����ʛ��a��CM6�8�}\��]T�Lw�La���y�l���iG�Y����c����Б�d��۝����5�!B�{�c11t$�a��7����R|ܖ8=�A�zht]�`��w(�8�(`�t]OQYa�a���kؖ+��~i���c\��hhD�6zRV̝!m8j�|� �i��K� �(�.�㡩�� _@VɎe�M���#��<>q�����:�>`K�0<.#1�U|t=�<T�#L7���\�C�����1_v�ۧ��*�J2�%��r�N��zw�Pr;��"&��ȶ:��͝|,�>��D�dvʾ@���}_���]���>X8%�#=�cm�Q���Q���
ח~���oBI�wq�p J0^��aE���H�{��4*g8��*��+NYd�h�ҁ?�/�Zt���j�1v��O�;�O���ksL�~�gj��Ib�rB�S��.�ó��a^����ʭ�]��ă.�'�S������>�/h�$Y��(Q��:�|܎���8�e����\�V���@\Q�[,	�>f	x�b�ϰ�Q�����Q�$�7f��L[lh�wv�/����M�ua�F����h�.+3A{���!�VA�ѹ���A��7��kI���Q�)j��ǥ&��9��r.sJ�0w��m	|%Й�����&��h���	�M�"?�x��q�ƙt����2������ �yc`���Q R�b�6��4��c����խJR��W�݀\/j����<Mr�&���r1�C`7���L͖�z���N�oS�͇�F�-�5���`)[��]���tS[K�B5�5}1Co8 ��TN�n�d_����L=Ё}��������Xj&S|GSB6�.
	�O���?2+�.*��C�G� �2r$/2Y<���QbKH�����������(�` ~B�������8f��?��p�����	1��y2  ���\ƯEX�m�.eɴ��˶s��"�P/A��C���u#��h����~��ލ�3�A�����  L�����d؏�пH�����>=@!؅�Q����/KK��Z�u��!��gXĝ<��3�$:�F��I��_0�`���_M+��d_fd��=po�k���	'��}Ѳ�Ц�F��`��/�� rr�\�~@�%��n�ïht�3U�i��'�,�|��?ޠ�Yʓ~�rX��~O���x����پ	��0Py+v��fҭ)��u0�0n�>�vvt�X�mn4>�_l�Fd��a%fGC�L��8���q$'�S�"��}2��(����Z�R�٠Ե�gOpP�h�l?�,Ѷ�c�,ȾYt#O��\�ԇ/��"����^ouT"�X �מ�������KV^.Z�
�`���
E�(���QuDm��]>_y�$�Vn\��w�&�%GJ��:�-	�����SV�WA��a�qFE�~����A.���g�u��I�ȸ��4����q�M ��s���ͺ�2G��BN���+��.��8Y3ι�i��l�*̲��8�jв����*6�I�F�tTT
Ȣ5�l�c}��Xҙ�Ѓ�a�	��^��g�Q��[�KV0����;����d�Qp;Y��"�?�؈KD9;ĳ�uۊ_�ʊ鍷��z�Ã� ����^������^��샦����O,��3k�Ex8��r�[���U��Ә��ȿ{Ae��܇J�������d����8�>�U�
瑫9nK���m7�C��h�(��H$�����i2D�^5`-p��]ݰ��6q"
<��{�w}�d4Ӌ	�b�O��䗇�K5v� �	#Q����n������([�c#�p��O��� �s��Q��T�Z?��M��O�R�e3Bp�~���;�}�W��	��M�[��H�'��_��C�E������CXe����FϞ��G�R����� y�Mz�ӔX/7��&?:��v�=˿+�?I�z�(a�y�w�5�q�Ѐ����:7�y'�t
���z��Xx_XN����[�4 �d�!��bT5*��9	�.�6�L��"���*�!����b�|�\Z��6!���%_��
c���P�6!������3�m��v���{T�3�3��r 7bx����d+@f�k�$"L�s��׏_�v �����1����oWk������s������̧��K^'Ih!�Q������[les����kv{+�q`? ������1о�%�t�'V(��\��̦.��B�>����շ	�&��/��2-گ�7a �Øw��m���m�q&����%�n)����-��#�.ᅯO��8�Z뺂H(p��ƹA���ͬ��LEؕioaUqC��;.xd��Ф@�km�Z%�L��v���+�Cր,��dch�tP���0�]k2��]�k����w0y><:s~��w
D*^���u����J�fW�p~_6ξq���(j����������O���l1p!MEA=�ψ�,�N�"�N��ڃd�\�7�y
S`�%�zOx�����j�E���»���1*o<_^������ayX�7L?m�\����3/���p�_�T9_�+P�HT�q���y��MB�S-[�'1b�w���0��� ���������v���M� <������+�@�]���p'f���1���E���}�2�)A��Q��U��+1����d��Z!E�K|,ƅȗ�L���*io���9�a79\!��9�hr�6ܞ�{�A�p���^$����>�%T�g�����|��3�RR?�y4=�Ɂ�h�~�m��yd\�g��g�"w��X�8܀��9��R,=�2�Q��4w�I��7U�:��	8h�M�-"��6C�WbM��N��m邏ڒ8��b�P#{P��WK!l���z`=�Yg�ұ}����U�۰�����Z����I6=�n_��8����!lSՑ��:���"�~y���_w2?Ǒ{:`���l��"m��a�r6�v>��o��3�1�dI��*��}4��!�-������(�$E)�y��(q-
25�j������u��b�\:����+�����Cks̟��N���� g�te`"�R.�ǒ2%���d4A:I����P����3��NcXi�>�ڣ���,<Ct����+c����]qۺTO�������Qj�7O�d�w�X2Lq�����y��!�;}^	H}���-��	K��5����1F�����D�ՇS�ED��&̕�g�&~p|���h�a�= g����W��֣�K�[#	{��$n�e����(1W���|Սk���P�@(KFY:i��'yN�Gl��+�j�y���1e����1)��۽�m�K�'�W�������IXA��*-?�D�kF�
�y5�-�`w��t�&�qS���Sy�PI�t/(�����hB���a!~��T�P��bP�w!�ٻJ[���J�������ۀɏ+���!=I�F�2�Ux]�\��[�xJqnoj��)��5�좋L:��8�5�DWg�I���l��a�;�W�i�Ǵq�(��&0�`?q��\n+��^Zt<�Zl�&��Gd�[3�'[cM#+�½댻w�Ł����$�	��#�AZ���Y^}�2=;mR4�)נ�M�Di�#-����2Ɣ��=��g��N7�8�֗�b������a*�u�)�@iOE�)�����������ōn�� ͻ�uje���k"��R�E2�8z�˄�Σ;M��}@�B�3�XI�������q����7;e:@���&N��[2�b�=۞+��o������M�N�=��������:>>���c�����]��[�*q3r��{*���"O����PO'�W��z<�iUD֭}�`�bZ���,�\h�K#�!|�?PΝ�D��Us��F�Ĭ�X�Ƈ꽘���C�΍�����/��nvhz6�x�PqӘ`SUA]�a���a��,��߾4]4����{-t.�~�(�UkM!7��qi�6���r��}��حdGu�7/3�DF�βb2�o�:'�W�\��g3�;>��u��I������<x�0�!�;�}5`9��r����΋�~R�eP�!SLH���׀+QX���k��O��u�g�EB���R�m�k;Ȳ/{������bփ!��Ԟ�d�#o����`�1�h�nE��."B떋z�Y�e(Gp�)�P�ܡ�j�x&�,��!C�&H��Vm�C3�E����`��$�GT&"Y/%DgM+Db��[U|�#�x�H|���a�T�=~)ʁt%���(l��O��e�0i�����*��E�V�$|���m�3��oQ�`��#�?�Hex��\�S�kj|9 �gˇ�8�?�8YRY}�Þ���f�Z~�_�;��q��I�⃹;�Ъ>�
�1D㓄qj<l�
�/��ay �5�����K}�l��~�Aڞ�ȇ�!����g���w�ώs�R�K:���
A��)��^�&hI<��ͣUOO|����D"x��������Z'd"Z�%Q�A^{��#�$��H���r�$?��=2�6)ihU5�]K�;��vy$�G{ՔN t��hf���D(LP�4}�����Q��M�f����5BqKA���O��8�fԑ��]�g�iߧ��r���F���&�0d � �2�ª��%�B�y���!>�"7�O>��AĶPw��;�
�|�{yEA�$x�[�&���h�_oj�_5��S�]����,�!1��ZÌ(�>��V�/L��-��M�/4��-^��O�Xu-�e��.ˍ���Vq���k�� \��T���& �Lt,H�Sy�ϖ�P�p��q{P��=��v���At! �?У
������J���J~l&k6��ȭ]	���S�m)��0+lY��3t}M�H��`�
�f)"��p���`α��<��9X���4�u"�!�@�~�����:�EwMu�V��X|�*��'d���^���D�{R�R�=����3�S(vE�D���NF��`S���6.�p��ߟ�������-�a�Q��=�qr�^h�>0�~����s�"��b���W�8�ͧ��t�(J*��9g��!��C6��R�&���7�[u�@���ø�ha�0�f�8���\u�2���5).|k�&��T4O�6d?�S?�E<Jإ�W8Y8Gy����'���_˜\i�f=�Ģ߹{�����Jt� g�����!���p�ց�]Ŭ*
3c�������B���w�j"�h_������2
5���j��_
�F�#��l�1�T�aKH�sh�z���.�7~��T��ݮi	l�@������d��fQ>}Gǧ{�N���K{���D������K�Ú�f�o��#U��dh�/��`�����x��;@��z�'���h?6�s�I�Y����7(_��(|F����ȷN�W?bWZtD��c¬K����u0�%���LS�!��6i䣳<�!��05���U������.Z)/�ѵ}��yR�XVP[q�����fR'8����(�~���U4U/~5��e�Aك�:[	��	��
�%U������J�Y��>�J^f;���_�M�K*��3� �K�.~j���0:�'`!�M0�z�R�o��I�h�:S0W"WE�l�g��z�A� ��z��_Q"���M���g�"^Ԁ3���`�2�������N�<�[�H.�&�P~G�.Qi���$l�X6|���k�ZqKT]p9�+�+v� C!�m�D���a�8�J�K�c# I{+�T����	���2e�Z�$-�.�1/D�%~�
�p#t�ԏ�T���ɳi-<c�6�HX�`|����x�������(L�ƅ��9�,wr��:��:��fE|��B����,����Qz�i����N��c��sY��VL���ff����K�*��xϰ�\Z�>�99�/@�rjǡ�WWY�8Ռ�7LՐE�x��؄�5xS�~�Z�7���A$�f:I�Z�3y���x��'�-�sFo���X !;�3�n��dq�s��͉pnOX�~�㨌v�`x2I�o����I�*wX�e�6���v��e���g����Q'��ZO�kn��݃���aa��Q	tG�7J3ss�ԡ�ݗ��Iй�䒂�˶������l���h�+�#� �}��b�E�GGH��Cƹ�Ћ 5M�R ����MB���(qJ���\v;�QUBM6�$��|�4Ϸ��	��|A2����R�*G��M���/G����/�<JE�z���A�cũ�r<�M�Rx$ ����@#�طA�t%��:������͇�PGXP��Y��q���B4?���Ȳ[��!�F�%�[�������@1c(t�>�^��Y�(��o����v7h�\��msQO�6��
>LH~w���T�	i�~�jF^�V?y��:F�4c#�\�hPӼI�F����8oj��8Qu9�P�����$\g��gu�� �0�Ѣ�4�pHv�-?#���`�v���/�h�=���t�"�[>��i���,iIY�ٷ5'��ίi�r-��A���o:����`W��1�=���7���bp=���N&�G��d(� �!X�H�B#�����<���4Z�m�R��ݮ[!��}�H����#e2%٥�t��O7`��6xP8�t� �2�U��!Ǵ��h�-�2SH�� ����͎dz��aN�俄� )G ��:�#$Q�ƽeH��3�Wue����^���w�i�]h'���� l�*�4�9%rWj���#��‡�ރ:�n��
� ?����@��ygZ��9���=0�%���|gX�fOhk���[٢rO�Tj�W���y]>#�O���X-�<�8%�嗇2W�_�k;�\���@Be��*t�o��;���+�gܽ��v[1Z�7� ��r3.���k��i\"�u,·�n��`�δm$`�:�!Y��5�h7�4�^c�&����/�)�m�|���E{AB���64Rw�sr<V��6��L��W��4���,�s�e_0��;8�fi}� �it�z����-���m�T�U2T�nb�����r.�b�L�(7p(t*�6�*x� ��d���c�Ϙ�o"߹ЇҊ��΄�Rݰ�[g5ì3e�	s
l�I[1�W����H�ԅ�{�O|�'��N&�Vu��v-�;�X�v���p����O��9��$'���̪���,Yþދ��������m�*�Z�N#v2� �Ъ�w)ל�v6��M%~0��bu� (�L��`�Zⷆ=���UE�K�21n����(���:�C����G�d�[d�z;�TMi�qsz�0���wO����Z��L)G*!�2�Q]+��|s]�t/�pcW� \�"+���G_���P���-��X����Z��r������ҥ͏^7��2�d����>)u����ߙSo��xk�˯t1�W�牗yW�~9���4�k����T�t�Ŭ*��O�۾)c��,K� ��&����t~U�Q��	6�{�GX�љ��a�S��LT�G��d��W�������Z�������>I�SX�A�� �t����ư����E���	��8�;��v��FA�O��G8d-�;��m�o��W�� ��U��1s��WP��Ѹ�͍V�6��6\��Gd�S�#9��JcT��:�ȉ3�X�H�@S/1��� �7\F���u^�[2j+3������~"W��B�'� �:�h��kJ/��f���Qr�^��o>�&,R�α��sV�,�/CzK��ޒ�t�pX"���TX��#sn�}���,^��]R,�q�{�	��'��8E:;|��co�m�(2��pç_�?��2�~��wTv�v�zA�?Ȫo�M�!���H~ֳ�޿����&��F�{a2�eZ��*�����p�q$�x�{D�{�����g�w��a���2FO��R��e53_�J%�������O��N[=��,�T9S�`/������-�@��Yy@���w%֠�D���KϜ{I�f��ϝ蔇
q�<B��Ep.c�6�Q���Y(�B��9�~v�Q��2,�����yuʘ'o-�Y�g�f]��w��a�o)��&�4*H���k&�v[��:JR�����J���$?X�B�&kQ̿��rA��o�u��Ie�i��`����uRd�^֘T#ċI��h��i�xg�˘���b�D¢кN���L��w�_�j��%����>�@b|�yG�=379�����wo��Xg�ԧ�q[��1=;3Fj�9�85��
e����`S���6,P�(�B�J���"������=�ŽlBc�&tu_�LZEu��Ô�!R�@�9-�
����4O�&F*o�A��Op�ކɖ�!�J�F�9ϒk��M������z���o|;�q�-0�3La���;)*��v�D6?:���s|�nmcO5�N�7��!�Q�n�D�i=�-*��Z8�I���X5�썞�&ǐ��c-��+nQ�X��E��#2�faM;\n(}���R�%G)�)���<�@88�L�Cʶ�;�� NK,���h� �V��+y5?�[�?Ǣ��$��Ujf��� �5�~��~
q��_I�{̘h4ֆV�e�~�~6xL�~iՃ ���t�ꏙ�gx��J3³��/�Y�Ի�)ȒhH;y��P��cI�ek��-t���!F�#�s�*b����/�y�Qqq�ݳ�] 5�PqnN-g�����w-��w�N�~/ji<ҁ׳�BU߭J�u�G��"1�K��x�&p�"H�Kn�P*5o?�R0ٯ`�qv(\~ǁ+�#CW��,:�Ǒ�]񱁖���F^���d�z<>�	��F\D�WJ��#i	��j�3
��U�ߏk���p�:&������x�Hޅkg\��旑;��7?9��+M��7l���4�B���Ñ����!�S�p\�G��CiL���y2��y�r����y������D¾���0�q_żM��,�ªo���k��֘����N�|����������G��^�4��LR��>D����s��b�]Q�i�fgߖ���S �z�g��Xm?�	9C�����GNP=���,"��ڎ�=P �)�ל6$�lmWdn\���I���H&x�/��ȃ�O�V��$�˶\��Y��q������_q�>us9�H뿱�V^��z�16� Së��<M�)���Wސ���D��%�X9�w}��c��.b����\����yImO�����BO�����ց�)�.�<k�	�_��1u ����=�@Zȫج+i����ⷖ�U����<5�k�|��vs�*jϙ9��
��ź����ZZ��l֌C�-wl����P��-D;�gv�ǚ�Ax�:���i�<0lW���+ht���3�6;ț4=�ؽL~��Q�gu+�ZT��C��+@O��%��ׄ�J���'�6m�59��Kq��}I�i��*����L`UI�+93|���ſ�#oO�G۳X}uo}�(>%]i��&V�jl�:-(�d�T�m�F+�u���:��Հ�F�4��S�ۻ��2u�*��E��8U��J�[~$	?�\ኜ$]Z�a"L~�䨵,"���������Ҁ]�(O�b[Q�˿�c��������F����ȇP���3���?�͚����nsl�KU��Q�'r�⥋1�]�V�_\!|��!ź���JK��/��T�,�6\�|TGE,��)2�#��M����,�r)�#7r�
�۽#���MB��n�-wx����A�u��B�Gd.1��'�x,�Ks��4(e����x����Ycnkʠ"g)�b�R�Ҭ���V���J⍹t�Jq􉐖XG�dIe�Y��v���F�?`���E����}o��c��v`�Aw���k4O#[��Z�}u�0��Ňl�E���8�V�Jbb���^�`��$��_K��-L̎p��^�>��^{^��Y��⒧"9�ױHE�(nY,3؆��\��I���*"�����,ȑ`)�L�o��)�9�*d�2M���-^(Y���x;�&;�����lŧ���������so]�Cl�x��4I9+�aO�R+;p�a��"y�xl��0��� �\y�߫u�q}E��y(�Xt� �T�xr%�+e5��U;�YYâ�'<�� `v�s�l�Y����^�h�#)J��YW����8��^��S�WO1=b�g�`�Lm�Os�j�cz��֕1���t��,����4�n�eٞU��ݧ����8��:�LlUR�1W�4�
����HQ��8���"����F�ɸ�7�$�{�X��9H�2`�8b��oty�E���_J燸BQ6���d�:k���_�v���@�Յ��م.W�����a$K#s���@�W
{x*��Ҁ�^29��zc�%�͊^ѥ�O��+�
��{�v@�)��Tx�b������!��Py���)��&s�o�s�ў�J�~Y7-4]����g��Z�����xÿo�� );lκv'��-0L��X�ޘ���,�$%�N"g��p���b|'.ɼV	�������Wٰ�����{mb2��ulp�k��ݸ�KK�-�P�&3��%�Hb�f���H,�,{�_��@t؈A��'��yvRC��ۻy�T���5~��5��qx��n�B�R̾c#�/K����N�3�Y�*�JF��`����5���Ҭ��������*�ک�t�P��PA(ƽ��_���<߉�.1f)���ۍj�T ��<�V@�x�d�H����c%!�߄p@���=Rd��㎪����V��.�ﱻPke��!��Q��S���4�,4�r�ٯ����1�L�L�|�hW�1�Z<��l�RT�\�?�~��}��7Q�<�^�E��2S>�zJܲ�n�^p���F���2���L6�_M6��?aWv4I��S�wr0���=�F>���4�[�Δa�g��N�Δ�u�?:�/�bQG��!h�`�M�	d�T�D��'�[2j�q
���w��󲉊F{�H0?�������84k��qi���9�{/���:�������X=�>��4|Zxp8��p=�LG��[���ojŠ0[}0��4�i�K�7+ِ�U�چ�C5`,z~���3Y���h�8�Ss��ܒ�����H��qⶉT���J
@:<���ދ@b4��,ݙ�����:�|+n�Ȏ��Y�1Im�	�
0�ƴ����ʁm�{����߽�`s�1�f�1��g��ϒ�P����cu�4~��f���F�d�B�P��1�j,h�%xв����.��/�wj͹�л���3��)��;S�R��� P���,#s-_� mg��nޘ�T�9��{N�V:)��0ךli{2�-3�q�K���>�7��S\obW�k0W2:����_ڛ��hEBmg��$FJi�y��2��c� H�=E���DB�w�*����?Go�(9��\�o����߼������nY�`{rz�t#��ܬZ<R��k��n��~������Di���%{��p|���{���`U��6q�F͓������OVe6syP���Q�b8�u7H��|!�������Jp������B]���wta6d��bi7P�1��=ah�_�،g��t^mѷ��g�?�[{x��a�����d ��4�1'4*�r1gT��ٝ��c����o�P�:�미Sy>
-̀�;���"2{�cD=��}L���X��JgG|:��
��,��RS���`����G��Ì���RD� J��}v��ۋ�
i�l5e��yj�E�Z�����e=;k+c�M����_�3����wTP�\Ob�����2ND�L�������|������401֩/�E؊�h����ߩ#UT���M ��b�I�F�Z�ƿ��2~��_%�����qW���Ӄj����:mT����)*�&��as������J�X��D6�Β�� o���`aP�@}�TҠ���)R2�9�~K�'��Rq1�u���3�g���e����`y�$;Z��7�I�uz�+Sg#0P�*����U��)��Ȁxb����Nf�z����$*��g��P	���N8zM�^A�y�p�9��F5�ݳ ��3�@l5���:�cR'���eT��Dl�yc�?$F���Ip���&�>Sg/�eo=��oa\��J:uV>Ć�O����]ڌ��F<��\�1KpII�w C�/<Λ�\� {AāZ��՗<j���s֒�oN'i����������8����.L�h�Xl}���M ~!�i���9��y�nMg�ʙ�<_���^j��u�3�|%Z���^��u�H����ɡo��Nl�}I�9G̾��_0��^g�B��%���Yx�'��Nշ2&֑�t�&�����;�N���ֽ���s9�D6�t�ӞE�ȥOCU|�/�Z6-%��,�aSFm�y߈6��m<�a��U0��RAA|cMd>4	���/�[rgfp\f\�3=&�ն7�Z��������b���]��pN���v�+cf"Yr�K6&Ҷ��������}�Rꀓ(�s!�'�Q��'��+;A��]�p2�v]}�3_��ǈ��$U!���xM	�|�Q���tR0�I"
��^��o��ޖ+�k&Bb�'�����^H��i;7 PG�W0s��NO��ys��$7 >�ő��D��k�-n(�]X谹��9�Q�3�A��!�tV�*g��ߛ�}1(v��jb�|�m��`1xse�o��Z#��G�謐�K�R���]�����M��Z���RF�+�m1�F{2�f@(P��-�j
��*X�L�3	ȱo^ԉƝ�������I�.��ڌ/����6W��V{@�VP�/it�J�:�ߔt��f�k}x"N-[�����nYTH �-
�wQ	R��$����,��ON�( �/q����E��Ѻ�vY���-��?��a�J䬱\g�<T^���+�3�ѮY<��:��<a�%�I�?(���.���kB&���8��P���Ss_7'k�i�m�ӶRB6D ���t�j�yf�!��`�>Y����Ȭ����z��Gm�Le/����[�<����n��:���#ڛ9=W�O_��0�)�<�TY~�{�{܋����ߜEW�6Y��{<��&´j<F
Lvx����n������p��Η��:LN�o�W"�*?��ߞ�1��d֎����Oܶ�J;�X���x�9�C�o��D,
Mp�T{�QT�o�̓Lt�Lt���
[n*��W��L�,a��.h�a�i�̋���^���d�!=(U�Ӈ�)���[�:Q�G�>��29�<S+c=CY�3�fg�����c�T
��',@� 05�s4`q.�b{%�ω��E|�̤�ل��޶��r	.�_i���^w�`֭dVMh��S'�s�cc�8Ne�b{r����VW�Gj�y!�*�ڸ�ʕ$���H	��R��q���/`M��ߒ�����UB