��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htd�����CB��Y�a	��t�g�0e���������u�7���1��7L0}�d��>�n<ǐu�
�sC38#�1jŏ��z�(��sGvL-�~�� l�W��+��8A4�R�['`�p,/��l`�#� ��9p���>wD����n�Q�Y��Z��¹X���M�]@t=3�i�qO����,N�u��cadGY��+}ϷúP�G���"
U�u.3~�2xi�C-������(��;tԞ�2~$Kyq���@r��.|���['5����Չ4��UD��|�'~+��fc�U�Є�O�LV����&y����k`#���h������� ������<�XG������X�W& �f�_ѻ��Ԁ�is���5y�-�����)����U�Y}a�ԍ�Z��kk���s�g�F��ވ�}�NF�V堎R��Bb��S��h���K�S�/�p���)����GЄ������:g�E\2RRY}��u�/~���/�K�+�7$[(�58�����*�����7����t@�8��.�[и삨xW��ʾ�s���g�[Q����3o�LL�ϠI�����vL2D/�KU��֨��Y�^2��*0n�~�4j#�]nr?=/�+į�"���8N~g-eG�u�9� �V���GϜ8On��g�dHN����P+�-��Z��y�q��C���ͬ]'�E���d�[?��ݒ��r��H��A[�y3�6�Y���w9�x�C���F�]�hCR=TM�/���Di�yځ,�����E�T(���@w��`Pj�7LC��LS��n��;!��W�@�5h��َ@��B����=J��V)�	���U= �j��̝�O�П��ҘJA�d;ڊ�<J;����+d��x8�c���0|ilp�u��XZ";F���)��+���4����,Z��Eٜ�e�"%���1�0��.(�ڢ2M��3�{��x�m�1%�6�؛^1��lz��UP������4�$36VYW�����i"8@dk~����F�9����i�j����#�n5q� ������#�Fr��Q�.�AN߯�6H��R�3>4h��Ѥ���Y�%f0�����q�yǐ(�Z�Gt؁I������B�\���a�ɟ�Ѵ���j)h�t���ŝ��Uϑ�����9�������߿�d�����ߵ�b�f\��>�lŗ- ��WP���7�5�K�)�� *����A�Ǿ㜼R�b� !>�/(TDi��y�eFm3R���?c� ���<�F±*=�U"�(��v�����YP^�m�T��?g�p��%��+��=�01����$)jz����j�e��!u�#�b�)�}u�������o��	���H�ْ�i�B�Ak�w�3p��&n�/n��4��=�'or��NP��{������P~�r��CA���	o"i��{e	�1���wr���/>�dz�z�u��֯�����sе��e~L�1�N�띝C��h^呫�$����Z�|�{j�C���h������^�����Fvf2���'b�����苦{���2`E�*C�*�\=o���qX7�=dFF�j�8��{ �H?�I�u7b�Qw5�{Ҽ$`W������wX\c�cI��+Q�1�>���3e���[L_�&��x� ��[$�Ѩ~�aŭ��y>\)s��tI�ZE.�/iGӬ�5���m�Hx8-ڄ�e>��w)ϐ"��A��5�����c����>\��p���:	��:U­h����rkꅌ��/|��$�nmb�,�F������c��[4�v���]� ��������Mub���e
[�o���=�+�{
?6�L�Zb��n������^��E�4�> ���S���Wq��p<����:��a�o�	̯����]S���0�C�o��{d:�EC�}�#i���9�5is�/"'�;^�؝`���b˽�mB���ɚ��X�ݱ�^^�uh�Ϳt��[ j[Z�k�Ǳ�����������ij�����~�r2�}/`TW�i_�*�n�
������P���+L�����#@{W�)j��D���*'�&k+��!��+E�s���%R��2�ES�y@�zB�1O�3IK4�9#dܖ�(+A�[�L?��0����X�aHr�)��%k\�V��*�(� 0S!�Ġㅫ#^o�!��絆3~]��8X���7|���}~Zڦ���͸���0`�1b,�%�����Ȉ��sa��_d��a�,�i&�F��ʯ��e�k�'�GN6��B��Ce�*�}�Ghw	�s��{�9��'b�h�6�o�Q�kq���}AK��ѩ�?G�d� ��9qcViGy�~���sa����b�vyX.�@�\����2u�n�P�r��)klFT�����L��.�Z�H
Z�Y���6[n/���Z��p��kn� ���X��*:�Ֆ�F4k���V�c �A�#a� W�'�X�M��P9����K��9����P�R-��݀?⢺�Ui"ޤ�;S�+�.,|�֗��_XT(9��v¡&;������Ɛ�[y�X�pFR�s)�nY����>;q�O]���]	FX���XC4s[;�Gg�,!��g�ڻ�!�x�6Q����]����J>=Uj{��u����N��HM�@ �%�rݹ_8k�bە��{�X�'lp�b
�*�`����Iw�z��eA%q���ҚT\�l�3�_����}�V�JPn��C7��.�̊�5������m��?���KPy��K����+c�K��;����R�&�@M�4�*Z-	G���?9��h���)�v��e),���R�\Ƌ��9� �q�q��Fj�xQٮ.�N�|��V,��ݪuK�7�U��,}�� �Oa?�)�ѬR�]�!�ư5 ���#Td��2��7r ��u�����-Z��:�ጬ��9�����Pʓq�L�_�hj4���y�t���{�����
b=:Wb��s��,\	��b�*�i��7�f[.aU^(���N�R�B0 q�F
��s�ru4y�c2����ۼ�	���KQ��ξ������б�?4��oh/�lN�0�����,*\A8V4�������x�B��C�1�'�A�&�����<\1��l���=��������s�F3¢VRU[�e�`[�W��-t�� ��R��`�,Rplߜz�����=��P*�L�|��6�_qR%�[��ka1|�OL]*�A�ి�џ�77*گV�pgfO9�m�'��+I���LY'���Cġ��l �݅_��h���8;�}��A