��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�۫k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������"0F��}�h'��8��<���9���-�j����,W�_/�H: 2���x���CH�^�g��$�Z�d�5��K�S:�Y���~��n	��]H�C1��C�#V�S��7Q����u��p�Yp�ľJ8�so��s��v���l�OK�i�ż��Q�LLa��&GȹH��i��B��K،Mʸ�qzZ�a��W�[�17�#>i,�,s�l�>�����4�Z��1�d�^��{֐�S��6Ux��҈��դi�{� zXh����\�%(�ܭ@�0�qyi��S�UvY��V�5��_\C>c�1��/�`�	�n���L�0u�c� ���Tx/]�ʇa$�Km��8#�S1�ܴ��Z��j2q����/�����C��b�*�#FDLr��"�7?������FF���a}Ŝ���_�B����7����d'��A�@#^������ݐ�S�p��Du�ұ�~�5{�N���K�m�m�
(�����������t��rqA��G�.�n�^������&y���e)%���<j��F�1�o���¸E��q�*`���d9���%�i/Ͱ>����1�I�S:�BI�A�+����_���X%*5.&q�$��-L��u ��
+��.b�Q�C[���o���������>�T����`��i����2Ș�q��5��JS���Y��-s���M����R�l����|��/��l>V�Α��Y�����ς��Z��6��P���;$ߨ��x*��~�X� ����E�zPi�*=]:sH��m���Hi����V�N��z�������v��Y:ē��ZN�3 �X�G˿����&��j�`�1�7! ���@U����-m}~G�����+*��B�HT�ԯAsk o	��/�*wۻZ�W���� ������<TnF)��8g��>�{��M���R�<��,+#���5i���Ad|x��'/�;�����e�YJ���L���/8��H����ݽz���3!.���!(�V<���0c� S�&wVm˿D ��L6&#4%����d��M��O��p���#��a�
��B�QȠ�
9��TK4����#�$����̕X��p��t���
���\sC����q�U�$ڗֽg����������@oǕ���C&(x�U�gP�h��}�fy$�+�{渿��4I�P��'jA����N�TX���=}U�4Dz{���3�������e���US 'C��ӵ!��&��A��mT5Q�]�<§��){l~ )��,m�CX���vȅrVP���<+��N�1Ǚ1&МԨV�5���nҲ�~�:(�x5y+�?�F@�L$�kX m�%�4�������q�^�'
�o���M� ��Ǆ�ْ}JR�����2���z�W��X۴��� iSQM����s#�]��9&�њ��1Յ����$���T?7����#�Hu�hS�K��ӊ�̂p�4�d�o�EeE"C���G�n8�6on�U�&`Z����7�ds�B2S/_��&%��f]��a�̃S5�a�jb����Y_�̀e�A8X[+�h4V���l�Y�Uj랹q��d�O�C�ؙ�����`J^��,%͊��xV��UoNzs	zk;���T�"8��6G�HAA�hL�e�t�g6,Qn����rR+�χ�Pv3���[:�J�z�K�A�C� ^"fũ�\�t���נ���mߨ���1��ϑ\!��$<�R)��i?Ȍo�#c�p��XN#e�簱e����
��m�A��wx��O��G��~%,]h{�d �-������f[fb���F�&��3�3�P�\4��ŉ�Q����f�wg��ɘ)}h�%<K�Db�P~����ǖ�	ЩT�a�Y�xh��4	X�.xŔzӳ��?�ML
�Y�/���FMQ/&!��L�4�{�L�����Z�9.��F�L^;�2
 e�s�@U�%��H�葡;*��OAC腂<�7R��G\���1VǨbL��I|�>r���	���i/W�{���;`/���+�޾��d����&�M�H�_��Sz�j������/Qm���E��f��l��<z���w;*�I��!��@c�W������=к�Ph\EMV54�LG��'�h�z�9�P�D�CGp�|��X�P	�^L��U��+�&TA�j�4�*9j$�-�3�r�B��\q9�G-�W��(�[�����W떬�'����ɳ�����f�>�I�Z�q�Aq�0ړ`R4~8?zJ1�b)�^��0ݚ����B�~�s!đ�ZC��ΝS�+�2��
�̛��,����2U���גA���p��%��M��M�xL��ޔ�߈��Ϥ_���g;;
����Y� � %�� Ym���������I���JI��^<��=J�[�Oqw>�g��Ld��S���w�`vކ�w2#�#�{�3CJs0��aZN�p�+�/hql�u�'�i�S�\5���\;�~f��џ;�� �b�VPT�m�?r�T�v�]-�F;�Y ��qKN�T�9��h3Z%P�C��	�(�O�7���qq�E�snBC�]�0p�{P��G?��Z��_>�o�6�?�ދK��lN��x4R�aQ���Z{Ow<)�.W����K�(s���aF�����ms�Sr��-�����daf_��t�)���-�e��}1<��^�>�T�k�2x7�d٦��I�lR���iE��l�T��%.�e1�F���?�s��uu�>���4�넊�G��'
��9{!��t6b���u���̚�2|� W���Ĝ�	8� Ls7�E��������#�T5]�P�;�7l�{����7������m!�"��D���r@�����Ƞ��[/��U��}0���-�/"ƫ(ym�����w�]'���u��
2ޮ�(��P�p[�ӄ�"��<}�?���$�"�n^�
�ڧx���|~���2W����M�ϯ.�e��hKOQ�78���� �mǶ@�I�plaW.�\ ��c(AK���U�}�%��I�9�"qPZ�,\��$����2�7�� җMV>�x7���l�sv�}2hHԉ�W���%���\��B���G�JT͚f]��S!D]�6W�����gRX���� kf���d�CPr�ɏ��7���&-.E�z�h��^�����߫�[X�Ǻ�`�71.@��n�+��z|b�6KS��v8��N���)*7�J��R����Y�{r��T�[T�7!Ht+B�%chꦈt�<f��A�͓��s�Mu�<��蛣f��zޛ$0<&sQ��d\��{���*��ɇ����|5��"��\ct�+rr����Z�($�t2�N��8m��.�(AJ9�J����Drq�I���@Hx�| �٫�B�N�7/՛;�[td�Rd4O@�Æ[cŅ}��^��nO� �'�B��A_��NkI 	F3�]�XZ�U H_q�]3?	�K|~�G��.�7����,��@g!�=��Tu۾}o�e�J�h	a�XyŐ�KP}d���p�U�c+�e��������޻@=)��T�
;4f�y]��gs��;���{�<)��_�E��(��}Uk?��~15�<�N�O� �����>���nw;�����
BŞ䯉@�R���pN�p�a�)DM�������6� El�ު�(�Gl���~����~�b�q3�-u�wfN�RO�v!�5����L_N�h�����c\��_�]�b�ް�l�.�w0��y�rf%&[%�z�#8'�AG�,�aj�ջ���)�D-$C� ��v-��U�aC}������e�}����/,�a����(��q��?�c����)}E�pl
�l��S�'�`��8�x<Le��㐔�a8��ޤlGsGU�0c�9ڎ�����P�ᢆ�7Th��������������O%�x��J�)�{����+�+��ӂ��L�~�.E��#�p�ڞ8��^�эàJ��i�0�h���4O|b�zxr݋N��0J�Xñɏ�!�J�:�0o�0������9>a!��p���������m�C�݋6Z(-wV$���	LK'�)a։��Q�[���!�Y�"0P��ނ��'����P�|���?�����61�����s6��T�4�	_�wF�s��&�����AE�9����*ϊ��t$]��6���H����"e���V]�q]�7;��z�Y2p3�t��<]����)<6p����^�<P0&'�Kzj�77~*t��H��<����N2�E�x[�?����AQ$7�`���͋u~���9'�Ξ��	�ptK/(;8eI���{�~M�����YJ9�����@��B|E�Llƻ��1�W�-��Qa����"��|�5*��i5�G�ͻ
Fp��LXĐ���HQ���؊ף�̶e����ґ�A��t��� �_-}E�_�d���#ou�~)2�Ec�Gߙwga��-��+951=N�-U�b��@V��D7���A�$������������!��a=Z$�A�=7��[ϻ,Hf޸9L�ϒh��I9=C؜�;��WƄn��H$#�qv{D�F�m�EbK�ka�jn��!�N�KZ8W`�(�7�n�h�=��Nԇ �sz�u|_e��.�F�˝}�#���n�8�-C�K���z�
���UW��<a�R�:h��{t~2ٻ�3DoRg��w�.��2]6r�u�d�Bzj�B��jR�N��\�<�O�l��?�V�G���hՙ8j�#�@�m��$am|e����w+���V-:1��H;�9zUD��Sܶ��2?��^��z���8["*��Z���/_�_D]��Ld����m��z���-LLHFV�b���.݀����|]j�� X�q\�OB�+^~�)�*NMb:�WWDeL��[5���a'�|[�4r� ҷAq�zn����^�V�x�
�2���f,�&DB5��̱)���٘��vv���]��ӳ��#Ȉg:�O;�bȩ�|,U��y�V0@�H�<�;þ%�r�E�W�l$��^ˡ/7�J��>8u���+WUe3�dB�����{�UQ��rB`F��>��e&./��������͖L���F�qY?���8 =��á?sG��> ��W�f�l"����%q�8�����D�_+X��ԑ���/ʵ|��.�c��"2.��K���#�Ok�t�B6�W�3������i�s��zcR���A9�[7�O��_�6������AusI����?лT cB�B�;~�W#��l��[)pf΃�,n,힬�_ۑ�7�e9������d�efrYQ�_�xyF[�<�qÏ�ab�c�f*Q�݋i
i�4D �0G�Lcj$l�zٹ�O��m�f�p��eb�\h}�hM�~�V�d�$����uN.Q����܅���VGQF�������6�Ai���o���*�t!/�+B�:E��`���~Ms��w�E� �9Y����/��&�?�Y��-��+4L�����G�=g�j`C`��a��2lT8�����pw(C�l�y1�{���q�c�O�hW���^����$���P�$l���ճ1Z���ʖ�$A8vk!8���/ ��_�*
!})p������zaX�Y�;I��\7c��ʍ	-��������b=�͒	c�!�1y��1G��r�S!ܸh���c�b�BV�CW�ڞ�P�t/C�>R<x#7T����[𢡊�Ǣm��H��c����oDP�Q�눓۹�a����/�t�))�U>g�e9�����_�."x�3��A���>O@r�� V[���V`Z�
mq�xEey�h�r�\����1�!Q�K�&��$$��F����xM��a�L�.xK�ߵ��;���ƣO	>��rT��Y{�ϫ��F��J���׭o���P��������(�9��杝$K�؜ӛr1Hf(+���8�DR��Q<0D�& p��G�o��s��X4߰���uc�N�q�y�~�^���[��+:� �¸�m�u��oc�1uN
�yT�S�n%�0�<"����r���y���[�+%"�ya]w�7��.j"�w���U	�p�7K�K~ϼ����Y�~ʫ	1������Y��n�X����Tdy�eI�j��cYQݎ�u�����!b���|�?�Q��Q�OS
r� ��Ȑ���q�T@�WZ��v��|\�	�w;a���_����7��"p����)��@l+9�=�g���W̓����錴�4@}:�gf��@���GM���z4h�x�>.�=� ����<��z�������ߔm5[�*j���s�{�'�V��+8P�F;6r��1f6����e�o�W.���Ta-e��
�Y�@�A�h����ԢRF�*�ْ��ii����RK-�bZ�aʘ#�J����#u�Ƕ������KD�3�V�������ǁ������ٸ��#�ˋb�[���Fp6g8+���el�����h��W@!Z�TH�_e�_����a�a�%�^G'_��T�J�:��,�,�M�o���aY^�i-��	/X7���d���0�F��L�K&�mb�{���n�k�L[3�.�������6k�\fl�kF�-�c0/'��s6�#1hڸ�
�[���j|�Dc����`Pn�1���0��F0���Ha�����h�ӓu;)?�S����rEi��4����f����������v�}6av�t�>R�\�2��r��4��o��0���p��4?|2�)"o%`����~��[[�fI�&�3�wLHl�>�%�������P��|W�i}��C�	��^������B*�!7���q���w����.��|"��||
��?k�!�I��>}.���y�H�!���=; f��@ϔ�3�e���=R�2�&u���9��]/�L�w��k��>��'踪υ�G��׏R�K�[:N)�'̐��7�#B�)U�h>>?�l���3�N�����?=�����ͦ�".����ɣjYۆ7�	�0F� o,�I�wq�;F�4V�)�p�C�Zͣ��5({z�n�P"X/��ֻ��u�JH�"�ϼ��Q��d�h;f�ō6K�Mڨ|�����e���!_��d϶vDJh�q��)7]|�(�<����B���v��߭�
�]#��09]ڼ_��0��2�u%�nF��4_@��-]�҅Z�^V!H������wrVI&��6Y:���M��:�_$+��a��m��f��YV�r��<�����#�V��lvU2�t9np}?�qֳ�p&'�ōd'��U�i��2b� �]�aw�[����c�[������ԯiq{1�Ua��0YH�A*�����z��3��k�5�g��G�:Z�}K�Ҏ�ڛ���G�v��!�Y#Z��8��q+����|Ԅ�ԂvT����>��{�</�u/3/c��D J��)F$��ү�̌�4���qV�ɷ��$ͻ#!]1+'bWJk�2��˜��x2w �����/c��s�`��Z �h����'���~����.t(:Nm,�[��Of��OXN�W�RU����
Ҵg
{ߧ�Z ��1+�}#Q}D���ߘ3&.Nu��1��Y^��� ưiȼ�*�W��< T$ŻAwysgj���|�,F�&��x����7�#hyP� �����rܻA&�clG�p;����H����C5�t�7���3?N�uSG/^ѽ�ҧ ǌL%rGl�T�j��ڇ��,�R���Jv>`Ѐ�X��@�Z($R=�(��٣nw�𲋜�s�d��}K�zA��V"k�9W�v}|1���FM��$"�$����a��7,5��-����ƀ�i� �Ւ'�%��ަ �Y�,�p��B'd~0��ӽ���K�4�¸���y���[aHR���Ey{�:�y�������8wƦAA�w𰻡�rJ���GN� �&y8����@vl�@��Hڕ�F۫�|��t��K�]�$�v�x ;=�0"��\Ҝ�H�7d�6V1��O�1~	�ܘ����L����^ @Yh��Jo��!�!q�(���`Z���]���H���*�葚-�]�QU�B���o� X��y����6jI$?��nޢ��T�������(~,�C*��w(k�<u�c�^�������Tў���R�p�����dd�('7z�9W���q.2��v3���	C?6Q��%��7Ń�?,\��cԴ�#G�T�i]?w�n��`��w �˶���o���D#�3c��{<8}��ņ���(M$3oſ�<�/��������ݕG��5�_����*>s��afH1)�}�t�Tr��~�lHf0r����
e��dJ�i�����f���z����8�.:kLv���ĆC��l��!�"��n�tJU,���|���Pʗ��HsE˖7���\,n�O�;�2SX=�[�PAs��#Un�SO������BA����f{D���j}�p$���!���N��^���\���6���Q����ɦ��E?w�Kg|�[� ,d�m˻YΟZ� �2 �_�^-���X�ɏK�M\c�M_���:=��SJ���!L����)+��,�3�~�C�!nDtD^�w
�ɺ���Ҿ��0	}@|���-�,Ƀ�O��T��H_������>���C-�}��a�� ���'	�|�i��IL�ש���={l�Q�(�]<��BV���4�/O
O��L'��UVS�#>��7����&���/�jҼu�l�7I�.��P-�fa$<�=ʖ W������Q�#�����&�����O�cƼ��R=h�-�/�N9�
^9V4�)����$d"zg�����i��N���z�{�8��#/�5N3H-PA�uЌe8��:��T���H[@*�ϱ1˷�x��#���l�����Zw�U5�[b���Gw,
qڇ���[�c��j�g� "|�g�td�����5J��2�ӝ���`�U��
�*Rt^�`�<4��M8I+�T�
VU<�:@Uicw8���6���Xt�%e�Az] 3��6,Ɖ����ăR,��Sm��ikpV�����u7J���(+������e�s$C���5�*zʖ��q�%�%�n�3O���w��R(-b�eG�$<l�fd]FV-�q��v�0�Tc�(���>�z �0�A�B��JO�89h�א5:�}TYO[��>Op9�K9j�hty4�=t�� ��u���'����^ʕ�L�a�V/�w�ƻ��Q�0���/�Ȱ�i=݆�řqt���8��t �����8�he��A2L�{��D��t�)�[j���m�qi(B�ԯ4���\��{���"������5��&Y�ݖyCq�`q6?_� Ftdr����5�v�`mi���a��<#*���]Od�Bؾ�x�PVE���h͍;�;��E��b�1pp�ܭ�^b�6��Ti�Ι�?�:��Î�%�4��j�j[�cD�t77Nz�\�T��g� uj>Nܦ�#T=K�մV	����`�h�W�
~$�\a]F�/�KZ2�Զ���"�(.�h��s��
�F�dΙ[�Z3�B7�4��|����>�v�Fy�Q"�	��tX�] �9����U�X��J#�`��5	ad���d�!�1�
�af\��#Y����YnT�<���ח�[Js�dc�K) ?��>+�W}����5�*ȁP�v�-���1+�_JG>�<��y�30���Y�B���,!)Z� �M�=U�#o�Ky��>&F��J��s�b������]9�ʔ�h��hf5y.�|V<E�?��;�A2���z ��g���/�uB�I2^�t�+B�5�q`Cض��� �LG�C�YD��w���\xT��~�7��4�����wa�ոU,ȇ�����S����X��&'�5(���T�����5�4F��)n}�2�8	t#��G�7������Ϫ�g��c���|���V�
�q���&�Rw#�net*�D���\$�'H��c;���W>�И�8��"g���b
��W�3����R\���J\��M^��v8��%�w4��W�C�,BO�'G�G,�MC��̋���d"W��=lߟ�rf�s�C��J��=[�^��m��f杮Nq;����� KY،O%�=D���k���(�Gr9�=��0����3�m�V{����,,w2;�b�h�����ፏ�V��`���Iè�"�'���1P�-������pd��)/K��#r��'/�T�2�Rq-��`.o��W��e��D�$�w�H�!����k��Q�:�B��`�l�v�����i��=������x�a@��"]���B��̀k`Wg�?��^�˸���\6�� *�F唔@7D�⢍���F���3c�4|��/��]������D���j�g�N>��������l�0i��V�.��.v3R����2(.~�^�`YAdU6s�4V�v�<���Q�ɔ
�)Q;�'�*dX�5���1����"�$ie��>G�*�6�KB	c�����	Ѣَ5�_�rO��3U%lf��Ԯ,nf6%-/�u&%� ⶦ]�|W/��4�$�q�0
����f�u��K MD��"[����c�(+K;���*��S	>���|�� �����<.��	j�������<It��qS{��kv�����nS$u��r�};5�����sz�
���@6�?	���β��>x��}jq�Y>gv�Vф�.Z�[�fbO�[u{�4��*9�y���t�^7��Pk:
�G��`} ��c�F�c� z	���_�ok
w��v��![�I>�l7�`�Nb�cp�1[�*�Ee��۸!D���G�,��E��g4��K.i�t�ֿ�b>��]��v��dxCW�m�>#�f��s�j�:��Jr��V-���/x���\�
_��֣��l%"_��ur���,~P�X0V7��[�U$�d�[��<�|mَ��	Y�g<]nj��d2nR�A�sP�E.#����@���CIC!��AD$�<�_?JW-���	K�����{�^��wd!y������6��Y�