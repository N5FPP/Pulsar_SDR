��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0��`q�M�'���2&��Ȯ�W�4��д��|�6�K!b�'mY�`��L����Tr�AW��:�O�po�-��0"RW��q��3�+�f<�d%x\M;	�0�ND�P:|��[z*��ܳD0��o�Ɯ�?�t$�k�l��0�l�o������&��N6��@�vR��?�mKE\�5R2N��U$\��G&�v�,��*(�WztwXlU �|u@H��wڅ���~�D����M����Ce���ut��B��y�&:j�T�N޴�Gs���<���?�VRZ�t��D��A����90Z�lN�hHL�Q��$�J{4�NG�.�p�;*���"��D�J�炔Y��'��ΎPq��~�M��w�S��/�ADaQk�8"���r��|��a�Oh7��t�y ��,�z�1Qp/��ȏ1�Q��9p���Pe]�m\f��F|����q+�qϛ4��Qh\�ڲ�֋�NW�򂠼���fI�=�OA��k�D��ֿ(�Y̭zo;���߀�b�8.T��o�?��@�CX:�;���y���sLt�?��������{l�fi�/L8���wa��Td�������f�A%ߪ�B����ˣ��{UƢ�I%�@��������#�FiN����O���5hҥ�\(��T�)ƀ�ą�9������%�
�IԺ�;�
���O�
ϊ�D��7�?a��'##[d�j����rY=��r�3<M*K�R5�~�qaE~/R��[F�ג9S�p)��6:dY�O�w).[�S��FyH7��ɦ�"y5������`C×Mғ�p�{�y�ər��
o�b����L�K&z�t��{�ffSry(��VP�	;7��kd����7�5S?�D]�ʃ��>����xr}��+`�e3[��D���&������*Q ��x.�O�-`"M�a��jd��++9���J/)���L7?��5��X�81�3i��?��[J
ucW��	�����6��>���">B`���S����!y�:⁑Y��v+��ڴj��/������%��[�
7s�G��#�����q��E�Ǖ�l)6|Us5����M��A����~ۑ����+�b�{��'^7h�y�E�)�ؽ��-�֌���K��e�8/�qn14\���\v�&���G������j\����:zD�`˯\L�Z�G��$���	�z��6!,l-92頊ƦZ��}[�(=Kņ�B2�@�`�5;��*�
<F��ݵ&�\� �����Iaa��Eu�w�!��Sz��]&��2��5�{�������5�s���Z?b�)��E��d�y�b�3��-��VT�P���NJ�������iq�U��f�Е�[�ق8O��_��^���֖��!��7�j�q��ޏX_��58䄽���%TT;����"s�GCj���X�fW<��W<�#�ի-=�nú�%<����hK�4;���9��D���2`V?��z9���Ì:7@��Ƚ1��=�"����	�-A���nZ���^��cTKS�'~��󶓋����u�I8
a,KS9$��%���-э�^�tX�j��\c�t���"[[�g���sXD[����PJ�{��L��٩M30X��C�p�:L�KFn}�!���l*c�#S����Vի1>����Pw�چ��+X����xe�C8H�\���Nr}{*�؀B���x+�I�"��&�F�n|�ᢐ5�R��q�_�˦�mu�m�;.?*�=���*yY��؍��٨\9`}rɁI��U��=1��Ӂ ��#�e(ۿSDI��]-3c�}?~��%��ڨ2���{��ѐ6��L�X3�I��/�$ ��x)�RI�u�H�S1Ԝ���k� ��K�x��O:%P�����Cɼ�+���j4:2����]u3�3U5
�s?#����_Z��nm�����2a�H9��|g@R݀��i���M��q�b�a���j<FTZ>}b�CqA$?���]o��*L��e���l�|sS�_2N#m6��2�e���\��K~5|��{I��xWI�:S�Rg���c�t�8���MہQ����&�V " ^6�D7������x�;f�˴�g���4� (�}J��k;��E��_$����|���#)9��;
�?�����j���-�Hg��6=�Lz���Y)�+�] ��i�jX��h�_'�������GR�����s�uL������Ѐ1;Bt��߅�A��T��N(�O��)�?��B8�,�#彽,m�kӇw�Ht:椋yx��3jS}��AK���1/g��A_�Nx��R��&WQ'\�A���#�!�5#l�fuaK�*x�ٓ34h�u��0�-��D���fD
(��Y=���k�#�P��	
Қ��{�
���.�g�0٨��y���b:�h��ɚ\�/k]��,v�~x�ԣ�Ʀ���|�QYs�����7,��㋵�0x���@�&I��'>يF,�+��>�.��ǐ�$��>�v����!�'�m=�ܸ�-��N�)�=hװÛ��AW�B>y >#S�|��n��@����=��/�|�'K���4�	���
���a�_T�r@���
�;�_@m}c`W�Tzn�C��0�$�c5�W�T�q���������sGPR��d}�U.C�+�.�.��n^�l�����z�6�o"�I#�j��-q0���U�f����]o�7;��v2Sџ����R4��a7�g���cD�l�j��}���?�U}��r��������v��f�[��<j�;�0x��{��m�>;���W ��l�h�ˢ`=�]7�A�՗���V{��E8�;�_ni��-�f���y٨�vIT��O{�o����+�
>XE7��D��+����Au[�SO�)�I�٦�1��O�4��3=����˲��:u"�9k�����i���h������Ը�!+T�{+Tגp�^�)�0�颔�S|tug*���|! ��څ?~R- ������_c7�72�.xj:#��"���B[Y�n���_�9B��Б�b��k9_) %v^Wݰg���d+�Ņ.^��n��uӔ�O|
4��=�����T�b��Π�E0F"�˧s��#h>y�.Լ�U��b�$`0�7�N��Ϫ��$H���FN+�>�r��/e�ZÊ>�C����0�'�,K��m�鱞_~�Vל�6ݺ��cuJ�a��&��P�M����?��RI��<���1�b�������O�Y>�d;�G%2� "<z�'7+�dG`��F���<����I�$�Bt����t�F����=Y@�<K6kWejB��f�JL��T�І�X/g��R>����I+^c�z��8�נ�����\!��yy�(����e�)t�y���t���k^Tww��#3m�K��ﷸ�F�Y����)~�?
��������+z:�Gc���!|�Cp���BI+\�Y5��`�P�	+h��V���jCU�n�	���	���ޡS/|�n�M��I���.���dr�-�d@u�+3�	H��l��t|B/�%EL�`���b9�tk]����:LA���{Z�PE�\�悁O�Gg���\N��FO=���.�ރ��E��W$x�Al�����_�2����:#�~HJ��Eѻ�n�}�ؠ��(��Y�:�0�hӀ}�����?�8f_��c�����d����!�f�nk�n���y�Y!8�<����-�����KQvJ��X�atv�y<E�<���%hH�Gը�+�Z�����@2�m`�漦 ������!��r�M��c��_};��W��YI��Ph����r�t�>��y�!�t�l-d J��ď0�5�7�7���:�U�Q����b5��5�Jm��q��4��o`m�O"�>l����Bx�@�N��_LX�.c�ґ�A��gg�AA�U�W*����#�}$���Q�\��� e���@�m��G:�`����3�~���ٲ%��9+Rf��g���2-=��J��L6~�Yo��O��@f$�h��ԓ������P�"��	�X���|(�N�wM��v:8
��1�rO	�����FxȒ�L�����p⍗#���(��L-.���=�H5�%����	���S`����&�#w�<��x��%�SȽ���#d���k�Ɣq�ޠ�%���`m����P�L�"�P£8$�o���>��3A��5Q��Tu}]�6����#�:h$tilB f8��H�2ލm<�����&�0X�Fl�m�ꬭE���(��)�ؐ�����.�r����2,�5]vu��vV��9H��9����^�B�"�<WS���(Ck�/#4��%�No��P2(���>kTd���,07��Xh�)w��_ ba���>>�|[@�uT�@E��*��O��H��/��{kä?!� m)��&؉�qHe;Ęv�Y���_{.�(���s�W˳�V���u����"��Y��B{�){{:8�|�����������M�^��(�5���������1�Y�6�s���0%`6f�2%"	��4��b�L;,���$�p~>�f��թo��2�g,YS�O޸�;�88�@���M|���
�U.d��U�f���pB���h�Ck$�Z�@5l�ˡ��=��4
F��ρ26�~g�D��/�p����R#���M>�:�4k����j��s<�1F�Z�D�fa%�`���Wz0Bs�M�M7�#��u���1�.�U�<��kl.����:���`�9��xW'�uЊ�h�̥RMM� ~ǧ��#s�`糞Rm�y -?\�I��Gf�vcTS^�!L\�:���TӴ?�}�4(qi�<FَĽD���iw�����Ό��-�iQ^�dRB[��UQ��,�C�i`�Z��&�5hm=>�f�Z���j�_z���"�lg?=��%3g�\{)i���N(�����蕑VP�\SV�A��stny�h�r��������ş�6?�2��PHH����pX,Xi�~!�9��s�$,F�o�k1Ա,�eِ���.�Z����$|����j���b��(�m�&�\ƍ����:v�0@��}ʯU�49�J$��rɒ;׷�n�b,�]� 5K�����	Bj�9V�zB��qC6O2]�(�;�^ǁ��~5g	ENP��9l1/[�C��K�^�-����U�׮=3iG���1��>q�8�[��V=�^I��iHƲt��6C���_H�N-�5U{y��#+m� e�!����Xy}�
"Ӥ��+E*RM�|Q>;��ktf%1�ٳ��W��S�?��Yih���
�����&T���/�m��TlAx:��M ��H>�{D{j�=MC*�?�XZ����#4kz6l:�슆�� �(x$���G�ԛ�)iƆ��)���anJ�߆Z���7�9��g6��l�bt[����]���@�)�'�1M��I���F��E�Y�5�çBp�#qB��Dxc��N��,x��J�����y<hϢ{�8��
�-��?�� �D����8�9�A�a)|��]����T�H��B̀R?Dw���
~0�Q�H�|2��|�C��>���J�l�����6�~�J���炑U���ւ'�����Iwx��E�U�p��l���IO��U�iC�@Q%w��zB��;)=ޜ�>����q[��$5���^Aϧr�6yr��� q1r���\N�rV�0-"tL0�� t��o���#��
U�e	��`���O�մ��VxNt�̇Ύ��YX���Ҫ4A��Hz&m���a�Հ�E��CA5���$͈�\f��6��1���E6,��&�L�s2U�Q[C��tf\d �9%%���9�T��WKC�Il%xM
z��w���Xkt1��cB��pG�*�ֽ�yv����^ۃ':I�85f�$�k�X%�Ӄ+ͣ���<�(�(V��6Ѳ`���ѳM)f*���G�~@�V�����v���#U�3.�(5I� �D �Q�������M��NK��D7��`8k����aR�`��Z��v��������UڤL6����X�|T�B�*1�����SP;^c��z�P3��n'��}������"0���ĩ��Gt` I?��9ƄU`x�P_�����{��bz�y"B��V�t��Qxt�М\��^�-�o�B�%��d��p9���~��oeX'���fד�:�0���9{�+�M{T�ig���o���[nn'��s��f�%[d0�6%��C3� 16�����Q5 6|�t��`@�xz��T��pݽM��@��9��E�E�K�z���_}�z �g)nW�T-,��%���n�);�g'����% ���? 	9(����o�g�����jRa��/:�ȥz������$����Fm�~'��h�R]�C���'�F�d>)i>���~���(j���@t��L(�+�+ySv�{%���nyu��7K#��ڛ>�߃Lr.t�/�b�6��y�U*IN�>�[W��!��d�ŉ-=�`*N�<z�� �TѤq���T�;nj�?8�Zћ���U���q��+e��k���piB�4� Yгgce�4Jr�ٚg���{�di��[{*�r���R���:^��ް�KN�D�Od80�k\r{z�uD-��2�t�p����\�d0ʍ�_#9E;g�kY�3e2u�#���Rw A�zs�g?QЁ'���H�V�<�F������q'��R�܂g�a�f�#8-��<j��G���u�Y�ɠrxRB��L,�yG�Cm�ZYpm��SИ�“�t�(�ɸ�e�/9XR\�y��An�<�e�סZ0�D�F�����)���n���x�����+��,�$G�s�AG���tq��0�.�N'���'Z
CĹ{�{�D�ҧe"������V����8OR�S�MX;����Xv���r�R��$�iUd��g ��D�{2�����"��C�� TK��s�/�!��&�:�%�]b�%�iG�]A>��f%��P�#���5�^C����tU�{��3���� 
�L  !�����U�[��CTB�fH/Ub�_B���8[q�$�|��C��T�c::M�z��8�Y]M�Na=����SH}��C������+�\��o��ն�۶�����XHC�.����cԶi_�V�Ṵ��W"ۮ��u��94��5kd#C��x4�<x�ϴ
b�u<'��vi�>�Ņ��$�y�Yj)���Q���c�~��t�U3m�gW���������n\]�H3�A�԰�