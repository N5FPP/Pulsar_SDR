��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+4ڑxſƆe�Q��fHv+�+Pn_<�x��Ԉ��5H��k�ځ��*����ʻ?Q[vhŜ��yA�B����3P� ��"����
--(a���@�_�#�D�pz�
�n�ˋ��窣��W���^��� #~����'�&�{�c T�%��w�h�&z���-g1U�ۜH1�
�Ѳ��%y�Z@ί�"�K�}�cAE�Kp�K	˰4I8zT�Q�a�Crw����P+7	Y�b��ב	 .IR��Q�a�o������r� e~���i&�qB�y�>W} ;��< ��M�Zh�����K2��*��%>��᫙b������R�y��ߧqSz�c�����j�M��X6����~���2���:}��4r�w訅��^7�����B� .^"�j����w7�~'�x�۽�vKO��ŲZg���S��9���Y=g�� `a7�B��I�yȎEá�0*~żf��_?��a�yH����e&N~�<�`X�I�k{er�z�J?�Ӏ UWÎ���S���	���U��`ʟ�
2�G]K�e:���P荫���Z�_�@P-���5����ϰ�Z���z~q����c���rqM��mZB�����cH'˳˖��Ty��Q���� �W�~8$ b��5�T�G�;�x�!IY����Q�\�g%��FOB%a�0�r���J�U�����SW�ˮȧPo���.�����C1չ�R�Bi�+������K��vuX]Jեj�����.�1!�2�M;�7�DX�v�)7-��eN���FM�z��]n��TO�Zb���N�wƺ.�TC��7��,aV�3��������[�{�G��-K�K{�^8�d��=fv�*E&]��Ed)�a����Da�����OE��HpS
��_;�;�~�e�E�#�����f�&"���L��"�+�mk��`�Br�5�G��G�d W���E�88^#�d�����Հ�@�[GK8�_ Z*�?=����u��4:N�J�61{�x^1��o8��z"Kj�%UH�z�nmtS��F,����C�oԮ8إ�3�=��v��x�2!Þd	�`	ǀ0f��o㩙�}�l�w�b�΀��,�G��͛�عK�eC\��S����L#]_d�	5���*���c
��P�½'�s�r��n7����QE�ӽ�j�֛!m�T󛅆;qp��l�:������f@Ȱ��.�Rd���&��������I�)2��QѾ؛./?7�^����6u�b+W����"�����lXIT�V	J$�c�>�	��4����	!�MG�>|c�;��I�y�.��7�T���ǋ�C��?�~ʯ��w)Kd�Qa^m����N�w�dD��9j��hs�>�k�����)��r��^�����33��@=1����πϵ`4dD�n��\�N��n�ϙRܥ�]4�Ļ�|V5\*��h;�mT��( �[zw����h�?�����l�Nn�$7;�(��KZ�������Z�s�E?	j�+�$������~��piTD:�|0�	�$���O�)}\�a��|�����HE�� H�٤yG��q���߯���pU�K�" �ۀ������3��IȩC�J�x��
�ث��T���<����!'��z� �@{�Q�c �fx#���%����B%��\��Ušg�$���y����QUv�Y5F���聞�a0��B���0}��� *N}���A�ES�ц���-���``�Sg��o2�b���T�]?c$�?L,�T���*6߯�-~_P��T�ȹר>��6��eb�ٍ�MN9ΗEw��#�"E��"*�a��j�F��۰���!�"! 6��sN�U�yŠ��ũ"�����N�=h{)?FP3�E E0���i�����y��[̶L�����O�n?�cU/��DP�2"�߁D5�f��Ǣ���l��Ӻ�޸�H�N�;���$A�Ls���`�Z�Co��79V�p.}���D��#Xcz��%�:�i�A�vڱ��zv���)N�%	u@UT	?,	��p~xc�[j$��wU����u���p�,EW�F�7#:���]�>%l��Buo!��݃�FnN;����m����׾��h��	� ��� 2�s Ը5��