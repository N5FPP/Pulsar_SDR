��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ;l�Fv1�Lژ�O���3��������F����Q?���b�V����Ţ� K��Q�G�D��i�o�Yʫ�|�F�V{:�� �{��LBB���Z��^sӽy/��[����I����k���'_hx\�Ƥ�?���ƫC8�r��j���?�[�b��Gk����s��$E�C���Iv{��Ϗ.��R+!9u@Gf6�e+~�7k>�_3�T�@�@����58fW�o$�T�h,|���z.yhb+�[��>���W��Oѹ/t7y����8�A?X�Xw��J~���k.W�$�'��(��ꉑ'[J��TF�S���o�z󷬓�I�UW���{�|�M�a���@�F�J�Q�tx�tEV��Z��i��lzt����#��I ������T0�=C��'1#"V,���)�r����4p1����Ɠ��LS�d�,BbD�י��)�@/
X����0�9�C�'�8�5��I��*���ŀ�К�;R�g2�9B}������Qj����F�5#,VF5~z�wY@�g�ږ���jbY'��&W���Q��p�>��@牣@N�#���Up��]���ߏ����\c0�4i���jK�tƩ�H-c�����d�@+�FRxY�,��~F��(��y���^�)P݈�k4<�w���Z���?4���E�}��_�á��š�0ޜz/B��Ѽ��#f�݌$��3��z#G �W�fĨ��H+hnؐ�&�,�Ɍ��9�ċ1�(ֱ�{��v�RF�T5r�����F6�}6��2l����Ɯ-pw@���
�O1���3��~1��І6	��v�A���@�e!����� S-����193��n���2aD��T�=��WT8�3�77�+��JK�eF�
���0�-:���%u}��_ǆ���N��� ���*c;��R<`{a{:g�U3���yI�X4*d��Y��˹V5{]����&�,�[a��hw�R����~��v�m���N	��\��^8B��%$>���Sƥ���%���ߘ�skF&F�����+���즀���< ��i��e���Y���%nr_��Z��Q�+2GR=�M�-����Dt���ٴM��d�8ގ�R�M����sM̩H��#*�D"
B���{8��N
�����+�E�S�8�o�M���N�;��<w��U��
���rܸU��zk�� |�T>I�m��F	{st�5��9�Ț_)���O�7��o>_��/��0Ѿ̆�Ly��I�FI�`ǣ���k������Y;)���?����S��-�5��w����_�Cs�MԳiV"��`0��ԧ���$�B��
�q����5u,�|��C7�랝��rh��|�Qa�2�v#�^���lQ�ۦl�O�YW��j�����J?�Zwl�"�Z��L�oؿ��p	d��������a5�"�N�`��*}[�d8C_���O[��0ŧuÛm�ZTtB9�λE�z��<�{�����;�Xz�X<\���f��)�
�1�Xd�B�ޛ��|�3��F啸��i�J!�烵LC����r ��'�Շ�6[�i�=ze�	���r�iR�m�Q�2=����<�,͙L>�LHEqb��V��n#c6��j�_רX�����&��v�+����Egw\��N��<��lƍK���[���LY0-�����臡��uS���	�|�o�6�s�������H7���a�@Z?Z}I=x��ޣ`?W�E��E&O�<
�)d����U��rRD1�Sa%�Ϲ6��'nLD��wEI&s�1���]��U�$]r�$,��2�^� �ҧ�6��R<~.ag 4Ij�5)�䓅�3�=`su�/���+[�o��!�z�9�����9�<�ڇ���ì����҄��K���G�`��M���9���J�N�Y�����E�:G&%@J�XIۃh����%�a�*�"b�ʃǌ������LL����|j��iW]b�h�����n:0b�7t��N��WV�f���]�к:h���)�֤L��%dQ��g�U���ӎ5��i�7�͘�h�T}F�s�&�-=tO�g�I��f����?��SG%�u�?7�3����^���"�J����=���u