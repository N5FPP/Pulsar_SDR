��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O`�3��_��Ժ��T�CFâ��2�{yݦ|���^��BE_k�����hd��B�ۇ]C�k�v�;��r��~�/�^{��pe�M� P����y��N��9��d�1y�w��a�qX+�$뻅}{��~����E���ϯ1ī�d_��|����Nˑ��N� �%\�V1D��8�g)��o��ô&>t�Z0ձ�ȥAO��p*p��wƚd_m��jP о-�z�"tU7�ܙ�-��Zk~�Xّ�C�{���Ge��ΚvO�G��B�z�B&���b��E.\5*�;�HŦ _��V��� �;$��x�Qw�^�_�ÿ����0�S�g>��Nk�9�@A�F��#=9��ǜְw0ɰ1��>�r���i8Ii����7�$�JTO�S����Ȯ)��B���WF���5���)%ݫ�]�Eh��P')nx�rp�#F}4F-�0�O8��3���uy<�[t�03]��Y�����VGW�f?A@�_�x
���'�	��(5��(��V���>"A�����&Tk�-I�.�$�d�`�Q�V��7J��P%�p\�oR�t-O$���[ �/JL4|�Ü��I�k������ȩ¤	��D�k�H'1Ƞ��Zr�:�����y���?������o�a�ǲ��79d���|2��D
h��pva��lǶ�}�Lf����0.�Y��r�x��vX�1U��X ��|��^�t�����k"/?[��愈?�!��#(E��|��6��BW|��W7ز�Y�%~旓p��2���wAU�a��?�#n�@��'����t�"_�du�c��j#}�i�-��=1��}��K)�(�3�+��\�� �R]���x����C☟��0���˰n���y��?eq�Zx}�� 9Ur�ӗ��&��2���/w=�^L��f)ؔ= E%��+!����͈�S�ĩG)�U��w�Uk�c��a��h��V�r��r�EsaLV@K��d�.ZR9\؆��'�����9��^�����E�}?
g���f;�p�)�>]-��˦�Kdo�`U3�'u��[4�õs�,h�¡��?u�znP����|���۷��������`��������5������7Vܙ�����0�c�ƫ� Ϟ���#�v�D�MyO�[�E����\?J%�|2����b���R.�x��w1���0Ct�吱��(�\�{����J�A�U�C	�YQY���|����h_Ҕ1�P�>(F`��a�+����r����Q��cۼ�fW���/r�U�4a~}Kn�>�Zq��w��@������O�ݒ�t�/��&���or'R=�)�^z�u� �(��!&#�]�_>����g� ;m�d�թ�d[Y&��a�jV�?k�[����[K�~z�(�7�.�݁�xLp8��9e��xb�œ���i��u��D=m��c����� �6Z� ��#�ԝ��Ĭ���D���KV:��Ѹ+J�S�8�A����=	8��D�?8��.�k5�M.NB���7'$f�-�ٞՅk�UB�9��|��G��P�cf8|?��_��)�b�.�x����[�Ɨ\b���^w]��u�zo��]����v���w��<11�=���#�r�Mn�����M��_`̽�|�U�Iꪯw�[���y��e4�1À�_�����>�QhW��ձ��1K�x.(F�PyEU
1�<J�~v(4�K� �L���Z�D�6^K�2RQ�R��Ԓ�Ǌ�K��Y���*8����6�*[�Ef�l_0ܖz�豯�]�ք��N��=�gR���2j��p�ʩ>.���E;�.�l����=A��iS�bɫT"?��K��h����5A��6$�ͩ����"X���d����'�y݀��m�T��^|�X��A���N�����1b랷�d�Z"e𙀝���9��V�/��6ߧA�#�D�N��{�W{,%�^ղ4���"�pq+�]E�T0`K��쑾�m���j�7,&,� �b�_��s�V��*ϋ�"����8 �1+|]x�Pn}�_��T|�:'�_D�{�(���j���I�$x�<�:�0�B��m����ݨr��B�q'e�Z��\R"�"�"r�QC�ڷ&�pM���6���L��6�z�Jփ$vw�M����DۣqPD[I!?�+��5/��*e�|�lM2f��/�v�G�*uQY���Kx�S.�7[d��[s�\#�3�z��\��` �,�`��&�WKۖj�h �ނ�:��"+Cy�ѬN�3�o��Y��YQ7exS�"�D�����@�Dr�nvg�&�ހf�H�&9�, �����'E`A�r���Ef���k�׎�@>cQ?c���E�E1�{Σ��Z*���x]q�@�f��s�c��v���\��k��1����|�4����@'���DA��[����k�Q�.�R�7]�-tx�o�{ޣm��ޗ���NM�l�U����zɈ���Ί.�Wp�_�:�BP+����"�Wf�)���0^�f�X��܂�@߄��=�}�6�#�������]*����4F/:�<���];|�����d�c��7ˀ�\�˼���0����y�m�4���wWO����)�r�eu�0莃$܋�`��0[(j�G߫�#�����zI2J����BÛ�Pu�r�%J<M���'�Э����h2!�e3�j�.�ٛĬ�[&�\hc�ֵ��,�c�p�aT���X��^%w�&���u�>t~ %cs�X��Ql����U2�_|�W�����n�d��K6~CD����̓�KD�~�=����l�f�x傔uN+4�oWk����饀$��flc�D6U��֯?��������
)a�ƲCV]o��!�7$}02W���Cn5D�?�9�
_F�����������gY��[�g�ßp|&Z��Q=rZS��f��{O�����&�T��'�����Q>
L��?���O&�ܙdLtvE�m�,H���V/蟰2H�p��m��fC��*;.y�?B%o�&�mEB�k�z=����d&��I��9�7Im�چQ����z	]UxatȗK�rn�JVnV�q��{a-����4�}��������� �/|`�pXM-=^ŴA��3V�����Nv��{���r;�����K����^O�2m\������]VDs\�Z�9=��=��qI�OjA�vۮ�`�fGK����xj��?I�)�M��+���5���Vԋ�vYV���LH��x�Yr�D°3���N��YJ�Fձ#`��%ϳ�Z�DΝLU2�~R�����v�#K�O��ĽX�\�,��}�S��s~��~�Ruf΃m���э�ۈ��Ҁ�V��?���{���5N���&�)�'�;2����ȡH��Wά؞�fs��Qگ�4���>���������l�.��������	�k�i6����<�A�{�פQU�Cx�|��7����QH�������n�;`��z�*��?_�vh��>��%\�]�+�m����OѦ�)W#���X�k�y�)b]�Sy4�,,!=/�F�[:��h�n��"�t���M��B��F7�=Dw����Y�
x�ܖ�Q�)J���>Cyʉx�d�o�(�6W"&Z$�g���jʏ^$p�aY1�L���8}�*�S�F�
�+�Ư���[U��
������
l1��"��t�Z�`y`zҤ��f������L�Fa��^҆G�t6l���I�L�8� )�-[�d*#�vv`��y��T��*C1��䂩�Q�LN§���	��2�6��n!;��?�����טF�H�?�\������{S)���h�,u�2�� þ^�����3��վ�7w<qqБi��U\�^���S����@��Ys���{�I�?(�H�_~B�p��	-O�AF�h�D��+�tE��DR:���q��A�P���s�>�u�KK]���pֺ^��P���ԯ�1~ŀ�����z�æ��9@� �%���7D�9�STPB�� ���߾GP΅��fsս�����%�������-)�����q"���O:�Bw�]�Jsu��UvtY)p
���PRg4Q���Z(p�;������F����#C0�}�Y��@Z�b�:H��a������Mv_�x̶��sD?�������75�'~.��SRФ��n�,EJD�"MWk��{��L��f��	��/U��vx*J�Y�L��m�qJ`"���*u�V;�h�vH�o�M ��(�D���V��Wk��Ke�&��V��G(�#
���b�� �Xa�a�k�pn�+�%X�����S4��bI�|`-`�H�ڞgq�-��D��<����w��kn��(̖�֛�xQ�~�9�x]uS�L�)N3}��Pt�9��;�0��)
�ʬ�99KV2ʂ��3�cQ ��s.NSaZ%I��6$<��e��]f������$����zS���um�埄�n��L���y;ωQџ���?��<��&�.C�83G}B3�y�<xC�%�G�k�hNP�W�����u�)���/GV{����a)#��JaBa)���铉���yB�.Jg�\
UP�g�3#=g�dx�TЫ����O�-�YL���
�4�g�c&�J��㞈k�����a�܏zg����0����c��2��J��x�G�5�H5���N����"��̽[���T羽-���Ն�~ �1���Un��DE��$�P[���$�2W�|:��G��~��	��iZ��ΐߜ����)�=����:�_�v�鱔*��gA����	�i��+8� ����r� �/���ܹ+D��/�Ӣ���`x���4��r��cʸ&�w��D�,�kڟ#���e�@�
C ��,ĕ�LWuU��
3�����B\�����a�0�Z��G��&k��ʸ��M��F��/Xm
u��n
�^����$*�%�ha22jǐ��	�Cd`�G&�����F����u���3<���e���9�-I�|���OB��9�a��۸�P�`��u5.g���K�2��f|�,�R5�5$��"�m� ��s��o�5�y������X�+�W`c�Ȇ���73���ڣJ@@��d�/K.*�z�gl��g}��ZbQ8�j��=8������m`ĊԊ%g��?�۫3�)�$���V(BB�S�)�{Еi��EG��fF[�=6k���рp�f��Us+�ˎ�V���v4[�������������!�����sR�O�g�}w�k٘0���Cӷ��$.ު�|t?j��.��M���u�';�ZHu�?Vl]<��8_z�~�	��]4ih�JY'���;�t���mW��&�%�g�HK�1����Rd,Icl��x��P~��d���	�Z8R��v�#�S�,��\��	�y:���m�� ���]u,�#2���X���#T����uj7`3�]K��m� �e�
ã
�X�m}@�ܜ_�$M�x��a��wϓ����BA�J܎oe�|7"("�$3 E�m
��w鮈Xҩ��*��:��9�(��:��D厂1>D�Xw��p+��@�΋�#�K�v�W�T�?�w�������JÎ�17\#���A�CM;��ev��'҉�ɱ�(�mK�'�P[Z���b��a��1
鲘
�*d��F�3
:�y�T*�'9�A{I'
�ܚ��ٚ]����f1b΄2\�)��[�B��@-�^����a^��~A�9s�tɷ�{ ��r����I���!�aY^����=3�D�Lx��E�̛��G��'����d�+�ӎ��I��>wX ɨp�����ن� �A�C�e�d��r���Ҩ��ݷ�(Q�)�ۃ������O��}�Yىʹ�`�:���%��X>�]Gٍ6B�=c��@m`b�>��1dU1Q8�Q�����:q ,,�2��&/a06(aA���EN����.�,+BN*�������pu��d���@#_2uϋn>=]�Z�R��ea��Pe�\n�Œ�\2GP7󹝿R[�M-����ɷ�7�1Ⱦ��q7D��<�gLy4�I �����%t��@l5���!�U�����q��E�G�r��.b��6,�ͳ�����w$Wc�+�2|�w��ғ�*c��>,�x�i.d,Uv���l�3���m���'�rd���_S)�S�gV�ǔ�G��HΛ
p,m�E�
����C������/��z"g_�~eiX��oe��F|ֲ�D�}���D��'\���y����)���G�p�[�0	svu�6�H�=�v�"�oRC��&��6[��X�ؘ����K�A>�s��S����Q}��q\7*w�{��a�ܧQ2�m�л�i�i� �o?N��+H"��o۸G�Vwh~�Mc�~%D�j����B�Cq��q�M���`� �*u0�iSX�y�<�!6f�*��x1>v��{P_F����`�D�7���ϣV%ٛH�= <��/p�,x<]�|��W����DF��]�;�U
,%�1ؤRX���������.,6y��[8��ra�������n�h���[D|W7���v@JQ�	�%d����V۷�6�#W�CdI�Ah,�5b��������r!���|K�����ŉ�b�U����}��[?���p��L����N"߹�{
3��v��py ��G뒿�H$n��2+Tj�a,�U��z���� �N��\�Ed\��6������6���_�_Y�h��@�.xR�n�������H�|����#��H�zOwW�\��%�>��Κ����D�D1�(�r}C����$�<�gX�����2O�����h�{��?�RH+��O���2�R�z���HXa��(����I�rjڛ�b/r���[-�)�B'[��M^З�~�~�����_}��O�U���� -3gb��顣'�u-����H'BO#O;���
�~�z�E�.��uA�8�8=�RG��BcȞ���
L�e�._TƱ���s�*�R<)�h.��,� z\��D��j�\#	��<�-zQ�U~������ow��S��~Y%:,t=Dvw��(�L��M�a.lJ�NK3�MV���OC�|�0�sbM�v<�9n������%�)���n �o�
_>�L������_�L�3}0!zv�L7r��t��x��l���#K�L%����cc	Wt��U���io�ʫ�#�K 