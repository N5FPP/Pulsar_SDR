��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��e�ik3�������w$����g|��J^]�n��0!+F���;�f�v]yTQ�ţ��{�~������kЌnm1��r�Lm��غ=~ �ŕR�6���q���c��	�Z��+SV�|�+K�V�ס5��� ���+c�sMw��Ru|���h�Tr����)oDA*MX���|vZ|��W�j��"��YO������XS��{G�oZ�����Qz��#�J��i�#�ON,3ŠkG�qB�Nl�N{��TD��f$�U8��(��|<6�	���ұ���-*�]�/�ֳDN:�������,.js��#�0xþ��l�#,?Āw��C�R�`Yc��� {ajD�ke�����|�Ty������/N�3��5� }�
���;�Zb8��Fi�{�����{'�iuہ3|-��,���3p��/�Y`�3S ��Ibri�At-�:�4`�|ܣ��~��_�q���0�P�i�*���Ư�)�I�.*�j֏�]���Q���Pz+�	� ��&R�Alt���eMB��1�:��ɯ�>�L_�mE|q�jġ.�W�v7������_�H=��?�r0V-�_���}ɴ����Ʌ��~Ş;��0u��5�h�{C�(���lR����s ��9tFp�SF-+& -.�Cf�����f{pUoCB߱S���Ez� /�7 $�?�α�"��L��_B���
6�Je�.�x�{N ���V�s�
�D7����{&i0�b�S��ѹ�k�&��2-�S���{��y�9�"D���"�2�َ͗�N���۞�����>�tAK�[�[]�O�����[8e��ə����z��@��*��y���W�>H�8��?�Hpb���,�m�'��U��j��@�ݍ��L��ε�2����O��1NL1'uQS��Ҟ҆{V:��|~�z�����SevE���O'�	�rN8,��Mh�]$�q����Q��~�T7�%�����@�y���9~�[z�|?,�*�4I��W���������޹~�ڢ�CPA�B~�*��]�	e8��ԻQȅ��\��?�W���ֵ8�V�/������N<�yڠ�rӐ^a���g=fL�kH<�b��� �U)%��;<�F�*������Qw�%��������זl����<Ϊ�y-Iҡ�ad�~G��%�2�d�X�#T̠]�������c�����(d\�����B}m?*�S!訪�-��n�4����/�����UO6���2T{�� k�ܞ�n�����d|r��o�2*�U�U�zxр�N������E��'�QV*�Z$�*F?{��;|���Q�&>e�~�0*���/����y��]p�;����Hi��K/���߶^�,����ϫA).�|(f���Bɀ��d�/Nt��Q	`y�8�=0	V��� G�I�-��I�08	v��'��ˇ����%b��8���"dd�M[�V��g�Ed|�LF�ru6��	�+!�ќ�eu
	c,�DZ���M[E��ԇ1��Un��˫�����h,D��a������g9W�^
��Q�_�����tX�ͣ+�1�Yp��E���=0���ܽ��#%T�-z1>Hr>�0��p�|����:�.I[\�Z�Ώ�<d�3S�Ȝ��֖���K@^é�!��!}��e[��ڔ�'���eD�z��u3E飱�P��A�r}�t��˰��\��?Ǳ�^U ~�3��F�6��?��5��,�޸
��>�T��/T�=�|K-���$�:���3�7���Ӫ�(J[�o���X��<�R�*��U?6�vDF�;j�3[Ƒäi?�O�)ɠػ�%�����.��v�庂��]��5w�W�I�a���j� &A���|�֤<��ޘ��<!D�⢐���v�>ih��J����a� �ّh���Q9o{Zn�>�D�9�)��_���'5�ڠOͱy]Eo�M��m�)jh�Y�я��*�mL�L6YP �L�G	��Dk{�v6 Yf	���h���IJ;��8�j�`yeQb���Eq�!Ut�Zv�*o��/��w@%qSm㰮#H�z�E���\u��M`VxIa��$fl4�ib�H��["�Ha>�\�e}�n��U�.g\cN]�8+��ަXޥ���(�5�q�[�=��]� �HW�uLIO���/ \իH!���ׇ��nƥCN��L�&Q��l_���@��B!�.aC�焢�n�f�)T,�����I��2V���7��Q8o͎g�[S
G�6���8�#շ�fDL���>(�~S}T勒����4?�E=�UJ�Lo��r��maa�;��.�(���~v�~�^��D�)t8���Wp-N��Z�F�WkU�#�ڱ�#��vJ��޾����ȧ�V[E��D'l�t����M��U1E���\��Iӣ�{��B#T�	q?���3���ȧ��D r{黟U��6:y�_��h���8�5��?�Y㙱���曊N�������0�p�b�-�s`�6����:��)�q��5f;��m��r&[��K�ͦ���R�=wpP��4�	a~��"��jeFO�n�ϳ��IL�$�Ɏ3b?(��"9�B�r��]�9��� R�)��s����u9q��?�PVX��j�l����b~�*&�=��>7?��G����b������y+R˛hZ?T���N�l����7��D�-���T���ܦ���[��bO�n�5��1��GL���N�꧒5I��l=��$.��>�"��70^↳%��I2*��q�Y�ʅ��}���b1�m��
s���y�� ��#ۨ4&ȃ��tƥ�Yj�i� ���g��z�N1����qJ�3����B��D�?�r�����k|��f����ɢXS�t����R8����;� Zi�L��->^��c�KG7�7W�{�øR�$;q6��Q0Z�Y������x��y�5�Zt�rE�|���Gq�n�FA;�$�+�������R{14.���R��"��n��O'��~Cw������5r^C�m-�(<����{��z�񜤂6��I��B��e���U��<�\�K�h�j��&�on'�{a[�HL�xi�$	i�΍fa9na�K�B���p�����PL�'��,T�S�����1[R����K��).a�7��6�-���Ǜ"D����2�FH��?���v�K���Z��L���y�v����T����3���H"dV���۲	krO�M&��g�����k#�٨�j��-N�Ey������!�>$�lU��H�Aḷ*G4xK��p2'����) jY�n�vP�pRʴ�5�q��A��MZɎ�B�Z0�i���+I����v����\��T	0W�5ak>�4���&�,^Ļ�6�I���C��J��O��nQy{�_:�'�ޔ�h����������ղn��. EԈ���w�x�f�]/{K�Et��f�����@i��D��\�p���%����P��x��#T��y��� �o(�U�� -ley�5C�F��s�"�����`�n�SH ̡��h���k��]t&�نn��cY@0z�׽�H��߀�Q���,N&UsY3���u��f���)�a�?�6g�d��D�2�}H��6���n��i�U?$�b������w[��B|D�/tl�J�o�Iߘ��B,,d�3��jw�86Rj�3�~3,Yc�� �[��2������ ��ϩenY��QW�ݗ�8�/��j�5��P͊c?bkC)>	�~�x�(x���5�7pR��C�CX�.*_�yod&F��t~3ꎵ[��j����ۡ���~hl�v'��Wq��+Ӓ���^�#�R~+��6m�O�C�S>�ɘ"�1xXϺ[;TL��MH��e��Z�������Bw@���N�a	������%�V�v"�0V�D����A�65-/��(l��ʅ�KY*+�J~UQ�u9ݎ���#��<�2_[��N���CE�;�X�>ЫP6Nf���O�)�[�G��J�˓{q�84�NN��@�E��-���2ީ�9������"s�:&�yG�#��  ח0BV��SH��xM৔ZynB����MU���L�^'�"s��G��5y�M��C���{u�����
[R�/��:|�S �d��-#�T�M�w4B�#��^�Y���*�d��]��|q3�bbb�"��SmI�)���Z�m2:}�fDjW��g�H^#9e��;�s�`�)��B��9,U!Z��htB�ǌ_Ư�����q(�.�~�F�?�C��p��I+�W6��%+�uc!I����_��+��]T�������/���5ls��S��p��#�pg�� e9`� �&�� �����:��[�b�W�M����*O�	ɽ�W��;Ѷ��pY<�@�~N]6�
O���2Ќg_J�5���"B��!��y����D�o�iR�N�<�7+څ�]7w�6U"��9�����Ru�6R:�Gs�gW�����:��1MM��y����=���qm�oU�����`�G��R��(��J�OӃ�b_�I��&	��-�.�AC��4'ՓCm��D�ت@6�k��8�1���!QZ卶De� ��1qK&�U�FK��6!�/矃�J@M�'J�ؙ��N㄁Bo�3��wq�̷;�m,Qx�E��tO�;�GZx�T�^�T�� CW�J �	:PUquU���秌H��G��Q/ξ�F
s=����f��:����?�Ex�������F���H��V��wԕ��,�[��X�"�qC�A;�z<^{�Kqϑ��HO�� ��~䧕�y��'�X���ڜ�����|Ls��ᕣ��#5حƾi�)B5^�Qcq�5�`��x�|9՗��r����߰Jtt_G_;��b�Lt/��+�ew=�w��X�D���q��9G{yG9�{Y�z��.&�'�it���3�ˑDo��&e�:��?�M�3�D�u�����b��Sxt��B�y��2t�Y�3Mi3��02q_�*�'�/����"	��\���=��`�J����%��o����WN@��{�&<(TE1�>��~g6��0k�%|F���*��o�~8���/>��*BT�uA3(����1UHWu=ڥ���|�h�I:�~��?��6^�ّ�)ϳN����Җ���y�h��m����I�����<Ι�z �����?�ي�M����Ci�B]7�<�2�߱b��Z#Q�Αk�O�G@/2�'Hlc�坙�G��,��҉�1��D���uSL%?F]h������p��؟��N���0�x��\Ǽ���lMp�6N�����K���rq��JF�G�R~d�
�!zڗ�%���)C9G}~1z6E� ��Mp|k/l���s�;�C?��f�=��s�a.⸅���d4!l��/Iʅg�<2�������hĭd�\�P�~��>�bl}a���S���~��Fr��la��fh�~����_��c���N�
`�>#�������z��.�S�N�),k��? ����*!�+�N�vKw�w��3�N��Wz��*w>�M�7�ȸ���x���M�ʦ� g��K^'r/P�	c�x��)�]��	��͟(*�w�"J4��=w�Q��r_nΦg^��݂$ZV��J�cb;��f��'�`�����]���ݦ�/�c�ڕ ��a�8%�1t��:cc+��}��*O�&��pF�;ZOV�f�@�������k���������{�9����5@�[��sP�r�P�n\��:�t�cj��x�9Av?*���(R*t��y" F�!�F�O)�L~;/��Էq�|��7­q�[��ꕚQ�zϵ-WOg���	�m�B�FpN�O���6�	�����|���Lׇ[��	wl��d���ʞ���3�8W��H��Qʥ����a���V���$F�����,R54�D���a�.V��
�7��.J�d��	�����S_(�%ߦ!�\����	=&���\6vo���!O�`��YfDtu譫�^c�������Q�ٚa|^t�#˜�O�j�r�,��Vv͠�Q<�4���U�6�X�u�6K\Wg�{b �T&EԸY�����_���b�Đd3{1�Ϳ��5���+'������,֊��@��2(7�e��rAR�0��1�S%4���L�y*Q��k����P���bz�
�k:��CK�7{�7��Y!��L����<�V��h�ެ�a�
.��ӧ!�L;Z�v[�s�u��}L���M>����j�*ݬJ�������-}�]��qor� ^O�z�>��{��ˢ ā=?��w4�wIcq��gӸp����k=�)��+��}���b}�8����J:�Eh���ةS �ծU�qO Z�9Z(�Q�N꛼�E:�x85�E\��Je����g�Z���"Պ����l��3c?G����Z�ߚȢ����+��?���{�������"Q��ثgO\D�����
���:28}�1 �+��� �W+ɖR�g��'��Z���\ѷ[[��W^����t+FP�QB�D��` Vl?Ԓ+��Qf��`eޱ��c���c���QE�T-�5s�&C��_}��_�7�	h�ۦ�O{od�>o�������Y�0�hl5�O��j�y���j�9��\���@����=J�p`�&j���k�z��oXP���)�فD��lQRa���F����T�F$�(Y8���o�O�` P��-Ĥ����@[�S��c�VQ5ILr�t%�e�UY����6�8�H���	�2�8 p&��QY��F�t�(f7���#���X*u9)��H��Ye��K�_��X�1f!i�-��Xx�>.�X%�f_���:���:�a�C�]���@����`�6sN��,�}V�3sBOxx)n�7�T7Oؚ�	�nXU���[`y�8�2AH���if	�9�������4�CC����y���!<7 �#�ƕQ3��dg� A�\�v�٠e�,:r�s�}e�#|��֨Lέ!5�B�<u➖f�V�o�йV��
�]zwՠ�%H��҈	񁣪
'�Fw�n�=�X�-W1�� �(�X޷�ʹ�E"Ο�s5)��T�V'���_��/�����"�7���W���75��� �ð�Bʡd4�H�2깱�]�r�V�*x!�O4�8CF?|$`�
�4���Z��UH�1�H~(
:�)H�<��~yk�^�Fv�;@�%Ⱦ4T=S�l1�Y��j�a�Z��0�T�KU��Y�Uݮ����W���n��^w(�mF�+�����[���M�����E0�SFA� �J
ܩTQg�*���6����ێ������O�hi����D�CUπ�����7���@�5��Ybwvjx�1|�:֟�5�p.7�گ�y��c�]��L�ӊaRE�k#������.W(�c8b$�Q�[�wL�Ix���Ϲn5�7+O�*�\���#�Ŗ
=��Y���=�2�H~	��A����e�t�2Y=�mr�;Q-��e�c���^���Jc��8�p����T�;s�F��ج�'y%�<jv(v/�\��li���+h'=�ЋE{4YN�s
&���4��^�^�
7+G����Ή -��]p��u ��܂��7IX٩�$��~�4�t�;å<�v�\'�AΛ����d %�^��$qj1�˻q�=�X�v!��ݚyW���+n���@R��He���,�X��U_=��m�ͳ�> z���|��CM�2b~�k�UBi"�G���@N��֓�������f��B4F�'�n��Þ�RĎg{�$IgN��\�7>/ʰV�Ƶ�Nev�'�/s�O�*���qO9�O��r��)?e��'��z����b?�I�#"�	��{@�W+ ��!)P[�{����L2$|E&-�Ù���(�2G�|��qG�� {���RQ�آ�%RN���_7�~m�@��7��ˈi`����d#�& �{y�s~���fu����~?oi#���B	ڦ�KƁ~�W���@�ς�5���Qi7���>��3�.�K#�����F�������.��|Z�Ȉ�U�܍�i'CE��#	d����sR�.����H�Zg����\����T[�79�>	��N�~J�ix�?��̿�ŀ�/ZO@�u�o���Rj��=�*�㤲P����?�aMFJ�A(u"ɩ�����e��#M�1|��y���� �6�ww�I��2q���6�b�T�o�Q##f3��o�R�<;#Y?sL��x2�e��=>�Z��o�Okta>o�$�	[�#�q]�?�j�] %598��N9L�b�i�a��)����j5`��>'R��O)XkM�� eb*��V#P;�9�׻�iϙ�8X�}�RH�ڕ��E�1�6 �:Z`�R� ���̠�D&e��;����<�C�JzB���f)�!v�mۥ�Aor�:�OM'1��Z��_fm�A�D�����.��E^iZ^��㳮���<xǯ�`�i:6@�	�Q�W���I��e�H�S�sL��j���y���f�n�K��YD�?��wH�Ҳ���Y��zr��^��E�n.��&�8���2&����Yƾ����~���f��]�nw�YE9Z�Ǻ y�r%n#��p@N
�|���%C1��L����+�w�����E*�c���QKR*�^�������׻�p��曙#����kң��~���Ӊ�D�D����FN��{�VxT3���I���J��wņ��Э���_��:��א^=|��
b��19gg�T3�_�<^΍k־ �nв�0��L��%𷈽����n�����*�/i9L�d ���5U��]�?�tWhj��+�1�N���6`�����G��	��O[�!"0�P�w��cVS�'��s�����C�6�j�*V��S�:�L���\�� #����S��Y+{5�c����k{3�f�fp���{���Ns�rvk�Z)�R2��_#GԾ�]#��PYTI�A���k���E."֬�$0W
���"�j���x5�p8��z�0 H�|ԧߞXȽy��]"���(M
�4�cB��
%FƸ�Vs��?���bE
��^��x8I��E%}l����4��!��	��b�v*���y��iɌ�<}S����F
|O���I�\`�WI�y�61��&���*݁�.ǧ/�Ud�
KIWs���0b�=j�'�=��x"H'�a��������wJ��τ�O.*�˱ʪnx�3�ӳ��TJ����3 Y��+�������ۧ�[�S�=�_b�Cغ�@��5�������e�,M8���'�1�&�g���'@���𢫶��n+S�Ld�\EJ)���s�b���°L���Ѝ{�$m-"ӽK�?ԗD	�#������Z�&�9��v���3�t�����le�;��P ʔ�"��a���h�$*��]U�AS�|-�Ƣ�Y7��}�����*N�:n���z���h�_�o���i9��yBkm��P�k:L�ئ�.c�+|: X��n���+B\���o\�&W����ǟ0���n{��_�'�W�*�J��t��:mS�7u�b�X?��FC"��w��w��|f���8��L���e�n��#��=�W���R����!�d�M�˟���%�Z@��Ke�ﱒ�4�hMk��G~K�����|'䟔�>N%��.�Y��9N.�<9�ٺ��?�pd"�A�µy�� WB0K_��)t�X�v������n1�
t����	Fz�Q�7?���
?:���.&�����3�6�^Sc]�2�LNN��H�7�虢����_Lʘȱ�'�x��N�p�9_|�{s�ʌFճ2
�hU	��ZiK�F:���	m�W���B��Z-vtp�՛�����YJ��oL�k)I�ӪI-�|3�,�`Ф��>���G�|��Vt��e
~����Պr��_�f.`S��R&�b�ly���6�R���C�b͇���	����X��Gg�|S��hH���r�1	��y�,���/:�#9�B�oD�Vv��~m�)��_�����hR���9�Ҍf �*FӜ���>$��
���&u���9�U�|�ӌ����G�rc9煐�S�q5�-z%��V_m��Ӣ�~-�|�\@ �������5=����0u�ѻ	p��������NFQ�o�+����_5��w�҈A��Y���YY�y�v1 ����΢x�VK�|�ߔ�j[h�a#������n$��m9I�WMK�F��y6/ dfX��y&�p��P���J[s����'���	�7�e�$����Zu�A�tS���q�e ���w=���xǰ%�:�2sc;X�	��/��snS�t83Z_k�p���0�'��þ��X�m�-���H�rU8iZ�t�w��۴s9���l��B;+
 �K�yN\�˘�<$B�<Y�����4bf�vDYr��|#o��e�����i}+������|���w�J����Or�QA�BUR�i���}�]�
�o萔j�\��Q�'N(3��<���G�F=7��iS�T7�HP����dϯ�`CI������;8�
���%\��*H/;�.�����F�D\�MW��t� L��aLy=Ô?劈T����¼ؒeJ/��R`勫�&n���|�"�j�8�`�E�K7:�R������I���������Aہq'�{�p�����݇�5Ɣ��S�R�V4Y�����9��
��D�%�Eq'�޹V��ֻ�j�{�;{�K�=��E���A�r�TǱ�T1R���� �/ݚ���#};7"�ñ�O'e	ѹ�ޑ|���ċ��wj�,ҖYy�����<�x익�x�-���p=rJJ.y��	gN����&�ƾ���(<�E�׍���Ap��`��ӡ@�������_��<���EN�Bs̬A������(�FK/���e�G0�aAD<���.0�{��6�*�UYz��R��X+#XWD�U���ZP)Lm�����Cپ5�ǯBsHT�%���̚Kb�'@s��@���&��ka�<��	�P=�5�-��V�"�?Z�����Z���Z Y����;j����]Lh�C|�q����	b���Ȕ�'��H��:�Z�_�y�G0�:�~�`�R'2�/���Q|�u㕵����n}:o��#��n����,]����c���QA�Ӓ��1�tCu�)��F�߼6���q+X,V$~�V��]���x$E��������Ԙ����"W��総8���
Io�V�5TjM|ܠ�#��c)����jb�pk|?t/7�kjC��wbG�5;,�Y�#l�+$A�:ɧ�����,( �a�:�p���>}�Yܓ�;oy�>0��ۜIi��W�(c�R�!sh��tJ�D{u)�������K�\H;X�U2������v3�N���^%[P��`�a���s[Kӌ�bE� <����V���&�����(���2n`�:�_���>�s.�>��.��S|ۍ�V�3t��2�Y�1��!�Eqd�N��Ě� H*(���$Y�C���B~\Y(ވߺ�4[X�
�{�K�ʈ��:dR?c��T�8p�
|���	}{�+�4&�B��XQZ$�F�p�bl��F!i^�ov?�t1_�*.Ū��2e��Q��w*!��u���n�g����O��n�xڥ��#��j����ݯ��E��$������w�gI��D���ED̈��,*�3-kj�Y�V���	#�"��@��6��+]�M��{K����@� 
�� =������;!���,{�8��+�
pH��9��TC���5??�
Uԕ �#�[2`1L�jP�l_��m��| X��v��O��i8���b�K �����y��wF� �ǝ�_Ƞ.:���P���r0�q��`h+sů�e]qX����ǢA�(���zi��74rVO�Q/=��MqO�چh�DdW�0Fz� ��L��Ox��?�A��tt���' a��}xF�b���iۏ�SKw�+۪ ]Up��*�'��g3�#�ALЧ<'H��~0���`)����PI��rj&��G��6�W��
j��&�3�	�B
�n,�ob}�/s���#pC�5�1��X
I��=ۓ�"�(�]uѺ�4����9Н���o��:���_���LSg(�{z���B���&S4���Af�f��=be�#�Q׳�����{UF4	���o!�"����Y��_:"]ea�d�ܐJ�f8̔c��ˏ2.�}*E��E���d�2)��=_���c:��EǴ�Ϟ��yzRO��97�W���$�Ō�HU�*)��9��
�,`W�����c]��P��OM�$�L3nj������T2�I�H��29r��ye���R�F�p��n���P����W�KI{*�Z�Ɓ���X��1��rk�^����ʖ�3����p��&V��.�=^����Y�V��C:����<���~yc�:n��\9��0�N'�n����`FK'���:i����g�N��Xrԝ$9q\�J+ ��� ��)�0�e,7�`����3����P;�A�u	h/;?j8��,$+I�Pk�XQ�m�Z��\-�^��jRu8ke�F��<8hoƜ�z����Yc��i�+��J�57��c����S��f�C������]�8\C��4
��^R����&�������"1�J�l���Rw�o�
�z��Z�<�{A��j��ɭ���8�	?ٗ�R�Ӧ"Z���_ d��zM�� �m�b�MJ#�8<lZ���[.�9��/^��+���d��˒a�ϟ�_���f�ǈ��me�>I%��Ky�T�ihѳ��.��U� f݄U|c(�w7�G?f%�=���8Lx�4ֿ�Py8ȗ����ع��]e8��q	6�������{�ko���ܹ $��}ǵ4�Ɣ�bj�_��IX.|ƙ�㢑H��*0�놤��|(Q�u_�q6��rB�+�pOC�|�!˗�M'�u.a��������d�R���`y-�Q�����;�fPk���RL�o`U�)��2Q��h��#W�=�Bl��ڬQ�0!�AI	�i�t�"�*X#������ǲ���Ǧ�f�K�)ڥ�M�4�a�a�D���W3���k�.��t����Y����&�{^�Xi���_3�y�C�s�k�F��1<�E�؃�#���������c OXM(I*	䋪é9	�2��I#�@�¦g��Jh��D�:O��JU2�P�~k�{���W��EzωT�O*�".�3$Ey~e(m��|�
\%MG������@��=-Ԝ�\)�ΡT���'�S`"�*@�+���M��,�2��0?�q-K:5V#�St=۳�M����A����lj��Uh���* ~�����N��Y�����Z�n��	���I�y�[���4%>O+�?V�^��6��`(�^<u7����z�%S�m�֢c�{'���l7���1�P,���*��| �I�P���5r&���M��W���t���
'��K��s��V{��9�G��P�@֏|yq����ŌYXo��	8wiH&�&-�8"�\^���/�3�Z�
�~Q����؀�EĀ996���Ih&Y��9�ef����9655�<�@3�$6�T���C���`�3.A;�Y89B0�u�f9�<�LO�7��-�������\���Lh%������jX�8W��Y�R��J�#'��3�e-R��L��S��k�6v��yB;�+����*���2:�B]��L��g��������w���͈s��H����9�N�FbU:�%`�ѹ-�5���C�Nv�����Z]k��:`5�	���~�.��pZ�q�Ve�\�R�]hXv���Ѻ�ckQ��NҌ㉿$j.�"��{Nة]��MƟ?������bdV���[�x��_��ʇs��Z$��3x�y���.q���Fk��HB���������c��ξ�>��;��YV�(����;�yv���V�!]�P����+	P;`��~��F�Q J\�G��+���c�*$�E�����(��m���:o4e}7D:���4������չ��\C�+�M;S�;�%�{=&n�ş�	�{A��F��.�O�ў���Ê��m�BJg6��u~�t����]~Cbb^9�[;{�Q�릫{*BZsn�y�+����\��ՖB�PX�E��v8�Xk���։��A{��7�M�f�g�62�Gq�,%�F0��������a�mp1-�W;��Y�DM�%FX��2�r+��[�W�cu	�JN���O��^�D�D;T�T��qcV�v�:�s�),�vh�#[��d޹�|Z����O��)�Вΰ�}�?5ƿ���=�?C��lD�^��<�H �=f�g�r��h�Z�����F�� �%��.e�X��.�CPKzn�o!M��n/t�>:`��������xp�%�1��j㈀��c˕�c����ȍ��F*�u�BX9���H|�{�S�5��\m,�L��-z���zLH��9���*��H\!:�[c�}���9���_�\OT'<�К���6<Y���?48q���M�ZG�8W��K�K�cX�]	�lV)�M�0��ݗ��lA���1"*(�3w8mRAw59(W� ���aKq=��@��Y|Bl�}C�na��C ET0��]�K�I����`u$�J�'����>}���V2��E���؏��t{�=p�oGC��⻢!����w0���3��zA�T��Uk��.��{�q�Ř��֢�<�CD��'"��YųE��v��F��:���&�U%������6���5��N�K��p���@���D	�����'�pޡ"y*w�`�i���x���ؠmB
�љWA�kF���̜�1ٍ�h��'���s�x�O���	k��ߐ��]wp��|:�*a�r�&��|C��c$�8[��@�(�޾Ii�P�-��0-R�ө���h���_2��zg1���\nޘ3�+�P(�L�����8�+���з�J���L��I��p��̚%D�����Hb*�<Q��N�;h���៹c���;v�r���p�S��7� nn�^Z��3�q��Z��~��mO"/+O�����q�; �\0�<v�>Y��t��~�?���5�1��;��e�{�c��f�胿����?f���/����SD��"I�8���B&:��Hg�D�'*�%��	J�ˌyz���@p�H^[*����-�K����,������W-��E�����@��[�)�V+s�x�?T��釾I�+N�UH����w��g�mY��b�&g�sH�t�f]��Ϡ�Ƭ�Ϭ�Wc�}�� F��5)���
�_rv{�z^ǹ!�.�&q��< D��L�]}�����{���]�O��5*9��AD�p�H���R�f{���Z@O�,�N��[V΂�@�E�v�s�}�R����A�.0��/���fbl���tr]�&`D�c&�_�7���B~��m��֏��0W[��I=b��*�n��kC\� -!-����
�R5���� >�ta0&ә�:���������׺]�ö���҃��h�p�2ϫ��H(
<	��ݝ�V8���şMX��m���6�d� �K�xa$0�DXΝ�D�B/H�� )+�Y�w׍������izW~��[0=q|�?c��Ӱ�XB4iJG�����z��<�4�t<�0�ꝅ0@�A]pC��ZuL��߶�&���e��
�%²ɱl<x��g"���+l?�v�u���UIR
��ל��{2���$�#a�u��#�FSW\��ߕO�J���`v�Š/D�����C[j{ԭٍ9�D�{�ӻ,�/���-�#�u$=���0N�#R)�ϣMQ:4�na� �}�+p���L��*&	�	�����ը�c�T����P��(�I�
8�����N�y���qH����܎3 Y1���j�ptI��J�B_��q��`n�n�K����[����j�F���j��9s�ښ��]�Z�$�|��;�U�}~ڡ��q�!<􇉘�g�5>�wg��2f��,Atz�Z� �f���h*B�l��T������3�pU)`��!��L�9c?t�ҐGY33ɻ��Ӽg�\�a���Fc��c$�,�����N%nPb�g]m��ro���3u��6!<<��ppm>|rT4�6D.Ēu������C7h`�Ed�h�q�^��U�@�|T.߸����"y߽ѻC�����$-|��e��#��J�����0r�����D'*�&k�]����G�}��<�R3s_�R�1w�-�2VJ��Xsy@����/���[�<zԗBX�z�:��!��+yc��\+3����ap�L��G}l���/�:�4�$NS�Ve�O^�A;97���&`61��|I#M\���u6�(b��&�53p2;f��$"�x߹d�D�f<L�^�m�G�J���ʹuPe����A��j-��r3��0*xcC��L߃�����!,]y��h���#Q�̗�C�_����ԩ����QH�6�S�KP"�H�4�H4>uM$�]��L�w��� ���\��Y��d��2�ͫ�� �4ʺ!���K�C*������"s�<�y���H'�2c?r��S��d�P��|�L>���Ϫ��_������pb~��>���TC�мs���x�[����㉉�C�87�g�+CG���}s���ox�e�d��SN��,Q��繡Ǌ���¢3�Rd�j~��m9��c?1O��p�O��Ï���^�}����k�(eCm��6�"�9��҈~��re~���g��h�A�����9�|{��&���$u{wD��m��������^('�ȥjI�u/v63W2аp�cx����y��)f�/�X{��R���8Gɥ�-��f���u�x0�,t�ة��ތ�b̨w���<�H�ʒ��z��������Y2��	��<��]5��>��� �\��ԃ�lG��o���`�!�,uZ*bӅܩ����%���\�~��T��&#H�ӻ�� 9������͉�|!��R{�2�UY-N�����(k�hb����h'��5��i�J�#�g.�3;� �]�r&����MG���7+��6レc�ڳ]=m{�^qP��|�H��<��Z�>1t�����Н_��?ǙB�<G������脞�)ZM�<�kw�2cd&%�c»�3x#	
Uw
Q�j��+g1t*x�z�V6AEM��A�CG���'�%<����O���)�c)��C�h8Q���/��p!��d*����Py�t
l4^��ȁ�!N��O.O�B0���2o����`Qʁ�%5�����gc��#���CUYu���x�[���r^1�%��7�_������z&v�ѱ�o�P����f�(��uS=Q�|��_��I�+���_����i|�Nd�����t�~ƅK��f/3�Z�_cQ��r<���	e��N�#-g�
�ĢI*O��?�%3;�K�]iP�/�:0�1��m���0dєUP�SC�L�,y��/#nA���d�ny���k��_�vJ{A�N �n?m�2f�j�2�2J"q�?�H���Ӵ,1����c�9���Sm4w~���V�; �>����{���mpص����Y�^���X��i���N�Rbe�DdM� �R����{z��zP�_����i��3���A>��{���Cu�1=��Wn}�9}���q�ٟ�n:7p���q{�@�v�8@�j�Y�6�����{�)Dѱ����n�]�(y�n�3Hܦj^I2��fE(�{#�%��������)mD��y�pɂVDt]82'*F'vr3#|0[�b_�@�d������+O8�_��&��%���oC�;� �A4�<�l@83�a �d%I�d�ĸ�W��,�3�l�^�Q��G#�O̍��Kj�Ni`l���֮��j��ޱdD�Py�u�Ѧ����1/Ba���K֘��=�H��Z�6�����@X��Z�+RG���!{�%ǒ�6�)J�7EW�Ӟ��j�*���6��bB�:ݝ Px�����kd�J��s���;/�[��*��me���f��O�K�ܢ�0G�}��tA�wF~pVf6����'������eX�6�]K�{�,��\K�Jd��	 +��f�-ƚl8%���p��
�͠�������~���aL�~�/J/Ǎ�&�te���p;j�83qI��[bR.a�i���ܗSZ�~d�c����� ��_�9����襠5�P�
���*^����ݱ'KD��5�.	�\6���)<πA���!���YW띾�}Q0�Ѷ�,K5�H}Ld�RC����	�(�oZ�C'm�m ���?�)������2;|p+�)�v0��XA���=f�^P#�򆖢gy��!��
JC�o��s�=��
���]��P4$5���s�.�p��i�\Q곒�Ĵϑ ��.M�}j
��Q��)��@�5��Bjs����/�ÒA�Ѝ�L�`����~ؠ=�~�����/��]�-��H���u�`>�B=�cY�3�>��PD7�)/�j�b�����$�^_��f��P�3��p�I�d��/m�9��:��d��3�Ak.t�j,����P�o�-�ҥ1�89˕,D�.�	~t��o�U��g�L�ylbs����e�O��O����<yL߻�� ���v�&����Uű�'�N���r}������r�����s����/_I��t��϶nlѠ�Ő�nQ�.��t~P�6,�L��gWL�b;�d������.um&ፔ���%�<i��LA$C����,\=�!��t\2�n��Ll�gZ��m�p��O���
XK��.���������f�n�? ң�/�FSu��>���w[dW$`C~���zgވ��7S5�z��`#��`��(�
{%ZbgZ"�
��!V{�P�Q�,�1�l)u�Z���Xq�ʇ:B�~0��R<�huы��ǖI��^N�~;B�B�U��`m�d7][ERh[��6��S�\	)����CS.�q^Q΍w9���f�7/�
�n���rB�}+����(Aa�uW�_������`ۤ�O���~_ǳ���P)Ȫs��5�!�PXl:gt8p�;�>�)��g�F��)Ȕ0����3�����6���i�e��o�`�W̆W�Ț`���n���uRkR��<h�c��j�6�Y�C�f�R#F����5�]ep���1���>���q<�iK�S徏�̙� ���M#� �o��)���,y^\ufS�4<t��,�Z����K�vC��������N�~�X��OI^��MIx �4�E5�ch�x��9-(� ��W�.ר ��7EZ�Q!ⰴ]�SbS���_�C��Va�D(���P���O<��+�N3����%?��\ʹ���K��,4���{�o4	�Ώ�x	s7�q\F��r'����M=t�[Wl�2�K�ͥ���-���v�=��&�ln�MZU��~5�Uz�c��&X�{�%���R^�s�m�B��A�-_����*R�!/�N�PT5H����E�R�z�>V���9#�H�8�ʗ{d�o�Q�
ָ%�R�/�`��.NX�+�����jaj��c����[�t�~�l:��*��u$�}a~���Q�P��غ���"Y�)����Wzz���.��k|�b�Wm�0�}/��ò��ܮ�`g�����WU��ؖa,�M��R�1�T�v?�(�h�hX��+�1�.��3���>�2�D�^
,!dG��3���ͮ$��g�eM�����oL�D�������� /�T8�_u���j͖���ޚH+N͏��a(ڶ˙�A��}�Gnl���2�QJ$��u���
�#'������s`c�'�~@j6\?�x��M���U_�43ϝK���ъ�k�;��媞Va��|2���C�F-����	�cAB�.[�5GY�a��R/������w
q�ۿW����[l�ow"�z �ֺ�睎�A��I=2b�f�2��~��Ƞ���ۼ+p	Zt�<�ifl�O}{x^��-�e��
l������&����Aݪ�U�r�֮��.*=�@����X�h�f������&�9ȲXo�{l��5����\������57%}���Z�q��ŹS2�`4&��ߌp������]h��\ǝ���w�m���'{胇���+�>k�Z�R!g�گ�M��a'1�b���VC;�8Q�*Y|9�0Cؽ�31�c���B8��z��j�Z���}0�j��J� p^�%�W���_�J��u������CTz�(q:��>ߤg����=sP��M�=��y��̸�s�Hu���b�:�9�	w����uMU�p6?�.��@���t��;��]N��ʔNS�q1�ä�!�����>j��f�{�1�5R�aml��#�Q�O�L�����o��%f�ѻ���L�$���*����($��RM��_%4Y;��Pm5��LIώ;kiych��3���]k����e~Ǳ{��ˬ��^�;t�ͥ%��a�^HvR��E+R�|%[���v�^{���A퇯��M/�x���C<�)T|�E��U=��PY Hn~�9�Ork�1��+�A�9 �5�e�(فH�7:'�Ux���!&���oȵ���_��s�e�gҊ(&}�W���V�l��=M�R��b�u\����8��b7D�Y�]�������\i�͎��G�i2Sޏ�(����4�ğ+R�_��'����rj�9&T6U|ڪs�]W�����(95�����3�om���R�E)XW��8+|?K�I�L�����x�����,L� �ϖ��� ��@�'}T����o��k�������)e�%�,�q�lN5��ږ��H�r��+�9׳�{|�^�:s�pv��q/�V�h��Iw��Y�ˌ�l�&�&����9����vp�<�}c��z��R���M�dd��Uy3e5�}[jAn�N�Z�П�P�}h邁���T³
�O����W|�;h�^/����7���üG Q�`��L�z)�*�V�N��x�c\n�6ύV�D�0�Y����d��ʏ�kPY"�}�B�X�����3)��7�!@�i��'�0�$7�e&H�߇{]X���[s'��>ۛ��-*I�)ؼ�!�G�_,
���2�5�fP��v���
턡%��j����>>bX�i�ȑ:'���i�l(�][�l����h���i�H�m�PM&�êc��O&Ty��c4~�~@��:/�$!�MKi<E�'m��̡�+NfC�z�2u�	!�60�6|�!f��0��w̴�5H_?��+�m������o�����e��H���U�,*De�1�r^�x�X���+��w�6��`l�{�M-�����Ϥu(iT�<�{`+�.�}4�I����h����k����0خ���U#����FC5NigF&�œ���;����Ƴ�h��5;Y,��F~#���+B����X�sA
%�*�f��~��+
*�l��S1��1u.J�����I��l�U��������[��%[�2��2����W�HDu�'Z���ʮ�[����	,�;����ۉ�x0%������?\"A	�e�c:�0�ǟ�.N=`=��]�@ew��������ܯ��'/.��%j.�Sq�V|�}�04��¿ӯc��m�00���Vk����Iw�)X��7Lhz���
|~�>Ⱥ"�Ft�>j"3�2hz�-�\�ѓS���+|�=VT�������e��׆�l�j��$�7���l���y�P'UXb������U�������ɬ.*����琜��wr�7d��>a��3]��IUAO�@�I'��3cQ,	 �/�nIE���3���a
I�4�X�c�Y��q����;��'S�r ��Xm����S�C�9p�P��aȕ��10�MH]��V�{�;_��r�;�؜�L62qx�ݵ�����������޺xĬ;x�A��퓂]�|��s8��.9�W~KC��@hEx̬���3'`3d*{�g�<��W�Z���&���Oɫ��Ƽ� ����xG����Q��;D��[�PaȬ�$��W68\a音*L��Ke��tG� ���-��fV _��O�f ��h��V�A|����Ch���dt䜾�ѫ�lj���A�O�X�ޠ���/���_�F���Q�;���f��)�� �?��Xgl�������0_�]�I=�x{�P �!\,��u���It�O��n�;�ݟ�;��g�P��U��w�O����Ș�!%����}N���6v���+���dK�[�\��T8�;�)%�S+�"�C��v���]n��<�\�JV�_r6�A;!�7'6N��!���ΰ�}+���5�\_%{�"r��s@9�r�?f���W��)2Q�Y�h�g2�h%�I���`j%�Ӻ;֒�<�җD��)2Z����(s��"f�9���l��cY~؋�+ �W0���t}�A�E:2-�d˼�<��Y�����kߟ���j�(��~�;�4��Rdú��_�?2�ފU�v@�8o��wPC+�����)R��N)�VCi��~�����09�gί�_��W�BT��Փ%�Y�)�w�K�F^\9��~�n�iGJAy8��B+ޤܧ��떰�t�#��;��������<�xP�fXꭂ�\�|�{L"��6#���P4p���t�����px��HZ��y��+���T1K��:�@7�S7P�(�)����|M=x�����u�:yY�͇o�R�`%�T����_�H|���LV�L�s�Hʴ3kK�o(���՝w!���_��c��|oy�^S�;�Tu��{����韀
t�Dǲ�,ˑ�u"��=D�;��1��n��'�=���Fw���<�mǭZ��w�������+��/JگԴx����f19���{�=��>$�l�f��*�B-uR����A��_�S"C0�)CT&��$w��x e�s����|�8K�P;�mV<�T��D�g�DNw�i0iBM"��lOo��������*,�8���am���kR�~	�"_z��rK�n�!Fzq����t|��DL7��!e���a9&�QJ���}�x��/�hw��Mb@�n8�3�_�����<@]��q�E����0� ]Dѧg��20��A6d�l+cy�)�����(��a>��i3�L�����Z ]SnUt���4��aj�{����$�PfPpd�	�����ǡ���������P᝽�}�՗�\��Z֠��6E�T�d�t��
R�Q䌹�[�PB:n�:
�m��6��fm��	�H�7-�{�lͽ�矴�k
ܦ�ЉE��3|�>�5x�s��g.p����� Vs3!����i_F����㳨�Yqd���"3+rX�1M�ɩ1�Q����e��:�����wwZ�ǁ��5�bi>�_�>H��:���[V����찄M���kT�Y�$2��v�����C��U�c��b��a�B���)w�p��٨���qb'����	I�[�V0r��h��'uV�-mO ����t(�Ju��Y�t�
��`���/g�W���Q#���{Lۀ�,J"0�$J8��7l����c���%m���D<�&=�)G�5y�#�Q�p��n�8�	Z��a,\0��x���[������_x���
u��2i��ea��2<znW.�]��]��/�)~6�4LGU��������1$��1g�j_��iv�@���B�w^ny�G�E>��~W��҉/u3M# L�v�v�\�^�ʷ����w�ww|�x��$�N�sg�Q��R��њUA��|3,6.�['\ԈK�Y5�զGjP��O��x���5ɵ�gȼ�Gh�g�P	4Q�U}��	�U٣.E��WF��t&���	���r�G�Z��p��Y���߄N�~���g`!����o��5RH�бΔu1Q�&����"���iـh�_������1��Eu)��*c��敛=Νc^քԾڰ��a?���>B	��9�|�B�\������2��y��mS�f�kA��)O���<��g�����v�D�;�kz%�kb��׉yv ��!C܄4�U9��?
��>� �y���*\�\M� N�l?��d�mlwq���l��tb�������^2�����2���q�^T��N�E����S��L"ҴW9�C���
{-���HH1A�~�|�ww�����"�V����T�ݝv��J��c�\�,S���խ7s�!3�o�lC�_[����-��;�Z�i7@�F�!D+����S�Q����K�LA��ZC=�;&�����R"n����_��D�ڪ&��Js_�?ρ�|�j���>�� ����OW?.f��U�j'`����L���,������|4�"6��m��j2YK����G^m��F��%>�y���9+�~ ��{`e�oYڙ�E^�	%#��q���YA�s7+���w:y7h��'f<���0�f��K�f�P��)$x��:蘱����%��O9��z�g<;Af$[�%v1��i��5?I�W��hV>��;K�6C/�Hl��0�����&��v,"t�ѡ�/˧#D��1Ͳj���Ln�E9���$SmE��d?�ٽ9��x;o���oo7��u���Y�6��k��!����T`M���cf��� {���FiK��ՔP���䈿�k��9^�ݻ# �`禩X�s��}��N�R����"����� b��1����0�g��t��kY��@2�!"�7�~�,�:@m���nޫ!Ԅ��b�G$�J�T��-�
D��9���Μ�a7V��[E�'_ ��qkZՔ���s�������b/�� �7ۦ~�^~�)�}+b"����
E������12R]��*?����jG����?P���Rb�Wl��C�2Z�S ��ȌQ�2>��<�LZ�YS�a_#�nu_��w1_bm}�45s�G��U�	�z(s��4��9E��R��V�SH��9�r�'��.�k,��i����۪g���]Ak�	I���ûY5ٯ�a	D -��߬6�=N�.J�t�yУ�bs�:�O�}��������䮲���Q�/N�NE?��9cAf�Z�"g.�C�����%��HK��tye�Af.J���.e�z�,l��@1��aV�d��5�Ɋ���/��:���G`A����]�ws<��.6~�e%�S������H�Z���}���5�5��`����	�n|�꟟�9�lAu�����d�ϕ�Z%��j�	Ż^�|��a�vͮX⇂H����3�!:�����v*%��y�ʸ�KC�%��K�$+�JF#��[�w�'��+!�EPâ�ߵC8�w��W�B�K�_@�w����>H������1�#����tnҴ���g�t�:���pW�VV��
��ឃ1�v��[U�U<'	3�&r-���Fq�Rΐ;EC�lr�v�7�'� a@$vAN�{����)��#a�Z)�g�l ��3�v�Խ���,�HL���d�z��s�ϙm"����R�]����;,n��GlA
���GZ� �K�x,wI��#\^ɍ������<p&�C�j���.����9ío�Lj�x
Ј���I@�[r�J�,:�J�����~i��3A=�ams�	���5؝��<��g at$8�� A�߱����J\5CAQ[�q7=W�k�]����;h����+���Z;i���ޜ�>�(�t�k�`�S�.r���S�����%�T	}�{������ZMB>}�׃�C��H�*f:ks���A��x��E��9	���z�g8����K9�ї�;�I^�U~�f4`�i4�8�U#Nyk�Ul����>�(��'�%]�"s�
�h� k�v�;�3 '>���B��`q��GwMc��ݗ�j[8P��8���� ���x����O�ٙD����>�+z���h�qr���Ic��:/�9d��!�b8�Aئ�0�?��ⶫ�K�ߚ���������7�{�c�(ד�7@�K0����E�15.�Z�f��S"^���Q�Ez�.�R�kCX���+����4�E8I�lL]ƫ&�@�᧦e��Ǹ��-<�C�+�W��@�Gw���ȺK��0����h�`"!
�R����9�ꢐ�5��ǹF|p�S2E��o�
�FoP��ʳ���.�i��U�w��k�D�g�檱wζS  ��j�@	�#�v�+�\fbf�yy�QfE���0��Gu�T ��_Ě�>hېu�a��(x���A��:�z����ִ���ٴޯ�`�K�q��8/��0�B�5=�ADZ+����{7z��P/2WF09&#��Z�E��K�"wr������K|��!b�hT�.:0TuMw�
����@)*�|k��:�U(�|n��z�OJq����.����?�w�-9$�xq�1	�k'c��Q=��;.��c�&I����:��o~�M�zYܿ�S�kuj$�m����9�:6�Z����'pZ�(4٪*�j�"Xff�r(R�7Y�S�����/Y~�H���=Tp�(��/A��yϑu?�T^���
c����jSLe�/�<����I��}��G������7л�l� }�r�Xp�C~W��z����w�'(
�,M����^"A)?�q���f���!͚�vNg���J�.2*��s��2������'�rW}w�F@@x��J�c%r
{O��_
^]ܝK
��.0#�V��5�):<��	C=I��Y������Uq@�v�ĩ��ll{�&m!D\�tT�O{�?��䒀�S_D��Z��J`�M{�o⟕�˖��gwyN����\�v#���g3|�L�㒪���3J99*��њ�����Jl��e*���7e�Xܼ�� 1����.�4@���@F���Q�z6���|(`�B\�@���8"�x8dC���������f�9�D�2�iHX��!��Y>���g��}��?'��a5�F#�c~�n$1�,��3eV���Usp�B����L�O=�;0��@jqy�Z�1��mV�W�c"z.��N=%Lor��O�f�(%z dY��Ő���/�3���¶4#;�i�y��r���kM�H/G�K�\��Cjes]�ȩƻ�E�B�P
�Kg���V�/*SҚyZ��q���z�ʔ%1�m2� ��.s�ϔ�26fg����S$Q]�w��U����WT3�����޸��j�{Ƕ��=���W�/E���D�4[gi�7o	i�q�eP�����`��ݵB�N���˞\V����
���Z�����W�~�ٍ�s0Z'�}��m�2����!G�1Λ��B�&�KD�d��3]�e�D���T���H��\{���g� 9B��D�ڱ�-�UD�W�.f�/5��j����|ߗ�إ�� i�ٜ�q��R�'N_[���2XGr����q
�g�j���4á2v�&eM�����bilK!T�%�Ь�:hq����+�����viW'�Cݬ�-+�N��ҙ6|K$V%Ju��a+4���C;�� �-)k��)���9Z�:g�C���j��H&#'�ƅ���&L����a���L�lڻ�zg�OU�%̍�9��%5�Nm�7�l�l9��E���[�O�d`M���[ k������@`f���D� v��<IDf��v:�?�{�W;����(�E�L�Z���1E�|	�Ɲ%�9��D��L��5���@39�p�k���l�	�N*B��Ua���V���D��u�+}R�����H4��NT}���*m��C/\�����L������w(QP��p�'���d:�[�u�G֝�\R�h@�)e��"����I�f��=5)�'� ź���������/6R��<]JLa��H���آ��upԁ_�~��Y�i�A�-�;��6gl���o��������3��~�8y&h���{}'�/w���ax�����p�1H�rB��{��x�4xSΈ�!��X��2('KR�Jda�ˉ�ƅ��3e� C�����b�gD�5��o.f���B�5yͧu
��_ز��(ndX�&��Ǖ72O�谵�n����ԧ���9���ԼR���L�x3 ��ƀ��NQl<���B*�D.� �:1 �2��$G��u�-W^�g��[{\>��M�Q���9!>�}Q��I������ʩt� 2�^W��>Ip^����U�`�ᜪ�A��\���� �3�w]����30!�F��~!2���w�d>�h����`�E�Q�e�jh"��7_�Y�K��8�U_.��@NƜ�.���l6Z2�X*���8,eX�Qe��@��᱃��5f�M)��GP�w��o)���E"�ʵ"�b�� ����+���I>R���F�ߣ�Hh�����N��	�Ĺ����\���5O��-GJO������Yim{bADa��z�K���e�Ҵ!f98���s�W��I�,���Ϻ����qzaeTY��x�5Ƹ/u�Y�CW�zdg�;����'���qtֺ�Ӗ�mD���p���83��~�1̆d��A���bM�d�^�G����x "����U��8�_�1���u5�2���'Lګ{��K Y�
x�>a>9��q��w����˂>(��{��b�aiz�Ï5�{�~�#h�L��81:�&Cr�Sx"-f������R��,�QGB�_�FÂ���+)��,5Ŗ�do�@:y8*��$9B�B�{[�^�?A���"!�kb;��ԋ݂_vŷ\߲,�5V%i'�Z�כ�WY̊=j�'�Rn��C��3̨�A��2>�����ž�"��Ժ�~�
MI?\��Pckh�/c�Kֈ�a�r�����\�3��zݛ��F�������dL����b�7��V��U6����ak�-��0Q+�
�&��>�����G�csP�v�ɩ���!��>��]s��Bf�FM�KW��N��Ō�#� ?-&��\M��5	���$xH4�p����W%��GY1˱3nX�MŪ�k���Ы��(�h��3�*W�h��0�^�9#Ѳ�PṭJ��1+�EHL� ���������N^=�xŗ���	�݁�xN�	��aֹ�js[��S���٪d͓AԔ���$����5�bp�y��6t;@Ѹ���H�b�s#����}���1�0���%4iwz��)L�#ݤ=�X]�@�Wob,����`a��gm�����S���Y,�&����Cw�ӧ���xd;�E��Ӆ��wi��OVK���R*8��0���7D,ǈ
_@� m���RH"7��3�D�\�7JJ}}͹�<5�)dO�Mv��p�����K�GIJ��9�mG�����!����-�J�Yt^�ᤓ���U�>8 �|���z�>+��c|�>�bTb����7�q �I(IU�*Y�'���5^�VT���=!8@M'�+GgR���������ۖ�����%mD��8+�����BjS	 ����䔪IOKB��6'3����=�>��hZ�{���)�ͭ�fKa��]�,oM�:6&����/A��8}�%\K'�����]�rq��(G����o���󾴵js{�V"�c�+?�\۸>&������C)�'�� ��XG�4�+X6�D�p�I	d��ֶ�'];Q֪�Hh�<���Q�g�+,�<u�����2�w"�C�1�:��2>ID4[!�A��$�b�k\��i٬a��J'"��-�3�9�B�/�����ꯞE�2��/����;��t���a1S=�����\;1/���&*��GWU,4���(}�͔��t"L	44�m:�{2#���Vy?!X_�t�i�9Z�ג�<Y B�R.墚�3����&ɪV���2e���렄W6�gΒ&�����w�D�x�T�R��-ibp����!�g��ڊN�DcC`mF�%!JX%RF��G�o`�m!l9[&F�H��b���T�]���:[������<,؍����#�A�%p������z&Y��ku��]�%�g�/*Ǫi7�5����|/b���/�]R;P�����CV��H�_}3\�WL�IYk=�U��s�s�}�{q��讯N�T'��	�ؕfO�
c�6��T<D���K5\�Wm*0nL�lCfi�Ώ�0V�h(I�7)�B^^໶wbqN���3���6c���x��-�S�5�r �}��眝�Ehp ����9|��ś�Z$'�E%�T��[�'�\���V�:�A�=�8m��]��]�;���Ya|�Yƪ�.l!8%{h�Τ�/Lq��F��TDZγ�f�":��|?��q�O1�C��*(jR3P]HN�t���4p��U�M�%���!��%G�)������$�T���D}8�� R�m
����5cx�P7A&n�@��̪�p��-��H	"u�v�V�Q��R'�>`��cq��K���,m�� ِ,�PAb��r!Aa�V#�/�Mn]Kʒ=�I�w�=��{�sq�`�`�Zb��M��[UՇ�w����^�]G=�r�e���=hj~c��I�jض9�Ý��qPn�
���:H�
����C��^Y�%�9�������C�=�ᘳ��d�
��Ec@_�٪�o&h�h)�|��ұ+
B�.Jq�j�t$|���1U��ψ��.-	_B=�{�p����r>�h�U���"�	E=��7Ni�c0��?�Zc�K�?n�3��\T��G�]�z3龢��T�"�+uG~�`E;��W�w٪���o�N\K����� U����׽=�0���FW�������䢶���S�B}/�j�N�n�4Hn��w�'i��'!Կ�.��������,��A����M�L���A�? |��KbZ')�	���"���O�L��?Rl�=�gN����{5��o4��O7��w�e�e��a��S绩������;����Ȭ��IO�~=�G,*��~t��Y�y��$|څ��ڏVm����S��zdP,��4;J	�1D�Ȫ�V��q��.�����[V=��6���=��쫩��F�䍈 ۄ4g��h/�>2�(Zw*��X[v5�`h��!�"�nS��eI����$��/A�)�߮zS�M��uTN�{����چ��+����b�CP�u�o���y��az�k�3y� �U�&P/t��	G��d�Ot������\��a\��]��ϒ!2g�^� ������(�e�C�hV�2���?]��E�3��r�B�� �	����W��� e{�T�v�P+�BL��B����4-p�x �V,H�H���x�Gr*P� ��'����N0��(N�L�Y&M3�#X�i<�*o�|)�n(W�	h�@�Zx*�
�'A6&3�0#��F�r���([xj�I��vga[�a�^��u�[ 9�_�e��/�2f�~|}�x��m/�&���W�Qn�+ԓ-�v�x�fC�O��8j�B�m���շU�.!:u�u&����G0V����j1�)�;�7Pއ����	��ʙ��(��9:Z�����Bn�&��՛����(.-nomz�� ��@�+����뱠�b��-a��Wf����Aި��9>d��	_��?��{���/3��-�Ӄ��+{S~if�4��z�K�+��������{�]&+=��R���#�<��Z_�S���Y�+%tۧ(��s �S����3���	���NUeҀ�=��r{�Zg�q����9X_�$��M�2�� �7+3fCy�oӇPc��=���$u���?�b���X�ܒyt�3�l�9������U>31�j(3&_P�1 '���9W�2Z��8\P�����)y��|�qe>wK��;Y3
���9_���I!C!,rvd�b)��sk��Cu]E�]���LA�[rYz<+
��e�����<&������t@e=�.;����髊!t"�)o8U����QO,�-(l�AՕ#%S�0���&�����/b����˪�ˎ��������&%����f2�0&��,�x-p�>�C��pSL�b+4w���^�����ه���󆷠���q���!W�1����K^����l���[�GϮ��\/���U�\#�|�Ba�HБu'��W6�XFZOwpZ����6ͳd$V�SE'�(=ץ�2ճbյ������Q�<�W"�I��%$_b ټr�UH�2h2�\�ĵ�L�0�Ӊ[R�\�n 4~n���l��e�U�F~�ݛces�B�nv���6vkK�}���c�@u��+'��j9��s��Qo��04B�1�Y��r�RFnCJc���.��ڞgGP���UEڽc[��_�`�rYx'�?�B�� ��?�[��� �t��Z˃�G��^���G�T!���f����vL7����oR�a�W?�l�uU��()gn�Q��7U�a�@㎇fry�>}A`���b��w@�D�ط�!�ȣ6�g�Wp�1}��%U
 `QyQг��e�]/b&,]��O:�EԞߣR)##8����~q`��P��Z�
ʬ����~��u������G��Ny��ޓc�R�-��'����l�������gv�י�oJX�O�.�����<?&�b���Z��?�w�>���d��v�r �	P}Q��E��㰇�����\�ٕV%��gk���o��&�=6�܇#�j�p���q��:`8�h:I�(3�Pth]Px[�N0lH�N��ʒ��x���o�; ���uA�o�C�1;�&�q_�T3����θ����9�KFt\V�@�'�� �h q�D+)Y�[����`"B4�Et��akg�� �iF>��V�`<#����M�i�q�)����d˹�Ff��R�mӥ�>�4��J�|Ԛ��M�����)��4�ԋ���&濇G�u�8�+�Q�=kb��g��ٴ�y�8H�4�+k�I�2v$�t�.ޚ�4*#�t;YD �����-��mV�?�B_EW�'�:Uִ�5�f��*�G"�9��' �Y�Q��B��4T�i�8��|٠��
�E�`��t�Y9አ�j����Qf�r�̑��K���t�:y��:᭴
?�S�cѾ�p�*U��|Ja>�X�� ��Y#]���X�� ��w|N�Ϲ��T��Y�G�s�8��-: � �.�MU�w�t�yN�8��b�骬�A���/��EW6��e��;��:+�N�@�S�i�S�#ٖ�N�yA��S)��]I�F����2f��E�ߝҐ���Fj���H�q����=%"�&:��{[Cj�J���Ͱ���.�w��#�&��BQ����eƐ�������3?;��4n�)
����:^%�������3���$���C������P�H���_o�y@
�?2Q����K/Y�:�b���{�;���&��C�:
R�=� 5�Ȇ�­Z%\D+���O�,`��j��_"�0��O2��n#cU&hc0b4�,@����e��[��p'Q��]t�vh�RP�9E8{|@�q�p�x(���8��܉c
S�)��[�C�S�B���P�s��fs	�67_�|���w �I%�z�Gjc��It�E��5�qv�b#'��hQ���I���5��
��
:�����Һ��y�|K��-�h�1	���f�	mj n�п>ܘ�P�iq�w�_��c�F�a��Q�gI�C𸝜�}�#��Q��o�o҃� �U�����|�e_K� �
2n�h��a�G��Onl�}�j�8�+��Vo�Tv7!:(�"��X�T;���xn���~C�k�����ޯ����E�JT|�tHL����S^Lu���v&t���6��,aAɯRߡ~�l������zJr -�*ԥyd���c�2b�D��V�$���3^��7���di�R�G���O��R� -?D�������I	��7��Ž~2�a�cs*�c��;��WO�����&M�BK�),������3����R]����G g����^��H�g��qc�%���"ݲ��������dK�bHv5�/P�:��@9`�S;cJ�/�J$��VE�~�����98#iE����Y1���wosI0�x�c�\@q<�?����1S����nR*�ݣ����|�N��H�w�̶�~��-���G&c�9Ѩl;�a=�w���" ޳�Z���$B/oT�讔<@�V��a��7D��R6u�Y
ʭ�?�7o��O�����z݃�[�vK�g�4sP)��x4uÿj��W �?J��y�У���L\{����<���M�o�~܆����Z,z�I���p�k�O�P�cD,��E��l���oo�������y�(�iC��r��m����*m��b���!:��|jv�yLV��vW��,��b�����̘_�M�qyz ����b����,E���"!k����(Jw�`
��G��z�`�m��g�L�Z�?L0��՗�����6�L��Y�=ؠ� ���R�]ٙ��"��c��!��mqSX�vS�?<X�E�7l�U���>��V5�i��ۉ-(�)���̼K�e��@=@�h�ϑ�K�.��&�~�g
���;�����^��'�_%�]!1׼����w�3,��8ͱ
z�<�#O����2�zuˢ�4k !�4�ţ6����)Q���Lڂ�wE�nb�zp���d�k��^1�	�r�U6�]��W>�_��T/�j��K򋣒n7�fe)I���\rԻ�Mr⩴����Q�������VY�K�� ,3���F��5��pJ��0��Adr4�Ēi��CL���� ���i��H(�8_Xx�ĹKY^��r`�_�eV+��8��)ME� P��ߒ#HkLJ��o�E��QQUQ��G�ŧ��<7�G����RI5��ru}�:��<��pSO��j��f��&��{(e�7~��)edYT�W�:��M�ɳ��IuR��ȟE*ͣ��Z���F����vG�[����q��m���*�_;���]u�c�Clm�M3�}$����U�ݢ�k�zҍk����P*|�6Z� E��O��@D-y�Mk�Յx���~���v�	�U��!T�-#���u�<��\Cvq���h���7�=��Z'��!�u����)�o�o��g�%�v]�G�L�O�}�;寖v6��2�Y͠~��{T+D�~?�ڈ*��#QJ�)���(3���ۭ���U�4�{���U6��~.�2�@��v�$]}�y�����MQj��)�j��ŉ���5�bd7(�1)�C�>�1�k��#�c{�8zљ��شw#i�q�D�61��d���P�>��l4֜=B��ጧ@#�);��;9�ۅ���j%H�Fǧ�I �r�-�n�/�`k���M ,a�{��q���Č^�&}��!��5+��zU/i����xP�L�)�N�fׁu��tf��ٜ��5��|*�Ti���ޔ�Ǿ���p����if~M9�a�U�#�x���|��|�L�H ��2\v�D�ǆU4U�j�W�#���B3g���4��;i�4}w H,��Xg���}bτ������`�+7��[@j����O�?�x���}��h��js�H7�hЎD��i��
�&R`��_BC�ń�7�����O�����5U{���T�I�`�*P������5$�e�n/_�~A(3�¬tW�С�DQr��3��Y��!�5Yž�	O��xd_Γ�m�Fȿ��Pd�����eG{����$4ӌ�9 .�(����!��܈g/�gM<-#�f�\ҝ薻!�y˭�Dx���j5-�w���b���3�� ��d��D^�'��X.^(w^�/ъ�G}a4��7Ok�K\h�y�j�}w��t!�����e(aC<�I�ߎ����n�pf�p�
-���P�&������)��� Z_�D~P���-b�^�e��=я%~���}��F����|]��8�lf�AUZ5[SD���ף�z��21�`,���S�Y�C+Ľ9���C�Xӥ�p�����'� Jr�(���𶎼��g4Q	'�?�\3�/��U��l���F�n�1(�o���fzI�<�51��&ąR��,��l�n�CS��I]���Ktl!>���.�.ӟ�q��#��9wa߶k��	���@����%�t��-n�F&b��~t�������<���0nJ����x��߉`��
�$A���߉z/qk���uƋzL0L�!k�Bz��A{f��k�ž>�F�O;A��o{�Ϗ�H�|�w�*w����F��<l�����ʁ��V\L�Xe͙�[��	e�KR;q#���PLqC�T[��-�ضO[��@g�U�wt^hR�O;��h�HS1)��܃ムb��e�ކ��7�Û�K�ƺ �^�`��3�['��
1�MM4��(XC�f�0������!�����}�v7Z��t�)��%9͐���`�',��$~��YN�v������cmo��[�� ���@>m�������z�f�E�ۅ5�'c'��\�Jf3q;D@��W��n�PJŁ����{D��.��F��Y��!G�j��A*xZz[�,u��	�7MrC��e5���!M�TK9�R���GC�;``Wu}�jϼ��\�e��r�b'ؠw��ȍ��?+�S5Xn���;|C]���haJ��e�V4�W�r��y�v�\����35�n���V��4bA@3a��<|��+O�BP,�N|S�Ǭ?��i��^�9�#qx1$&x����q�'�ږ�5UP�"=l����1�`�w���>9	����7��d~�:�:���ź�M"��R��&N�"�\��!)� �l_߉��|H%���9|��������$k]�3��'.�(rd��ȣ��c��dUJ�k�i$p���)q�h��ř��{�7N��f�1E����Y�����X
ГmQ��4�qxG�3�Z|�1=Z�=%������S
����.�ak��RԀ�)3���7�j�:��<�# �S��I�&�X�l��q��cT5��2���l�b�k�y��~�rH��P���>���E�W��/�� �Ŗ�J˅=��A��i��Rc��JXW�bU��\'��-!�Y�\a�s���gk��'~^զ,��k8ڠ
�?�$��O���3�Kz̀�7�5ҹlAt��h�ğ���������f2��y𠏒����=�/�l ]�ࡗI�j��'"��A#��M4K)��ЃNm+l ��t��1���#��[Bvu��!�������� bי��Y^	Xg��S >!Z5��������:�����I����Ҁ`���æ`Or�&��z��>���7�"r�m:��A��0f␀O���7b7C^�F�� S���d��C�����V���m�P��tȓ������P���3�����|�� Sfy�cy?� Ŝ�@̼*U6
v��_���L�����>�����b������|�� �3Wy�E;���a9��+z>�a`�����3��8}fT��%�N @��6`?o��@�^��@L�Ҿ��	�Q���_Ůh?@sET_�*��n1Ziz�����ߴ�/���v�&��Xe@�R;S��C���d �727m�Q���I�륁R��;܋<&b�z�Y� $��G|RB�|v�o�6� U`;U�EH��1~;�y�b%�k4��a`�*Lz+�u�=3�-��Q�D�/�Zb��g�>glQ\U-��;(T+�e7��'�����<' � �+/�����k���ғ`�����'A��4l4�#S�n�R�A�*U. �b�x�(z��]Md���u�&�Q�l����d	��hge����L��&���	wEX�7*�+��}�B��m�mB���Wx���<��� ٲ3a���}�Ի]�o#�����ְ2��U���e�xQ�W!���a�t�֕���#���J(�O�;�D��C/�cnR9g@��Ƚ�Z�m7�n��y��5)�t.T;tV�i�H�"�5p��Pb/�J��ĉ
��Ӿ�f�Q�X��"k~L�	�%b�ʬEBU�*�b����1����i��}��j�#e5��Q��;9e�ŷ�wgF����i���u�.�Ɲ���bfG����шQ}���h��Èp7�.�u�@N2j��C1ʹ���T�*P�[dE�d��0zy����O �4y����܀��C�3�~	a��2l�{��ϛ�f���"���&��©U��r%Ց���i�Tu7�
X ԑ"i�x%򕮶--<����F���w�4HH��°��#؁]R�+�鋹���̤���R��^8������>#Xh��a��n�`�z��Be\��C?v-���X�>jsdM�RB�?3a��k�t��Qh�,����w����Џ�7�@ڨ!��'e�+
i�hc��q�ҧ���5q��W�L���ݴ�.��+��2��!�U�7�7����:p���v��à���&v����ɷ=*M��O�Ԇ�����z!�-�7���)=,[�Q�S%�t mSMћ��S�&7��>2�Q�)x^�N��}��u��O������Z��0�b$Ѭ�ᣄ�؝d�p#b�|�"�8���W"XS?J�/ī64����y�jlG��L	��M��ks���W�٣�Q�������u/_j#64ҿAi�Hq��%��DW0l�/�&zg����(P�S�\�@I���@臒�;ƒba��f����#4�Y%�����~0�u�f�2P~ N0{�l��K�����#k�¾ۍ�t�1��ävN�6|��o%��Q���9��w���,�xv����'a/NWՙ�6C�2@�^�5�\����5��A���
�l�=�J�^�m����L%�0��ל�;�Z���J;#Ãj�.�_$RR���_�VnXvcB�#��]��u�Y��/p9��:��
�
��
���A2*h=���q�ݝ��.g��&�I��{�y�.EME�W.>��DpĚ�iS��&'<Ȉ�*��B��ɬ �>K��#� ��A��pH�7x�#���!�1u�m�8�U�m��_ZJ�|��7xʡP�o��Ig���n���I-G	�u�H+�-AR��ru�*���Y8�c�0r�����6��sm7�0E�T�}=ƸX�L�A.#��&�WA=<P����'e>$���XZ�;Q&�����
0
1��gq�{;w�[K��-A+4�ݍ�J�
|��@��W�/��_�K�҉�o���2wB��eb�$�<��6�|�+eͯ�Ehm��5�w���SQrIqa6���z%�f��Z4n�� �d�>���O�}��e^��*����c1���T8	�A{.C��d��>�XSu ����G�Q�e-�%A-Ѯ��ϓ�r��~�t��oI�I
��Jm �&$ePf����<�	���# yZ���HE�4�d��F�Tr�$*�S�$2��?�}�
�{yhX� ��J8%�KR��blј���;s��R�����\�xE�I������P�m�M�4L�RＪ��oB4�Kq�l,{o��T����S�R���rl5�A�.������הv\�Lq���7��@�X��_CNz�,H!�F3�*�g�+O�L-q����W� S��_Yh�N��[��>B*��[h�M<�=���[�m��Y=�q���Fp/e��w�ދ��<�QY�}�#��q\���&0���� ��jR��vܕ��D.uf���Ǭ|Og�yQi�d�R������?�Y�j��ڸ󊖞0}R@#�L@�夃�.�o�x?�#�����#x�[Mf�fΝ�'���0g�]8������q���	�W�Q��v�!p:R�(i�����F��5'���y>?%�KQ"I��wF~��=Ʋc���8�+���9�Z�;��g�u��X	�,��� z�Ԏ]J�:�P�h�����ؠ"؏��,�ʑܛ���I�m�ll�]]��.]#���w&�|�<�u|=.�!������H�`����Tc�x\E����ɾ>�2��+L�ў�vb�;��ZW�4J�{!�	�qI5��R���
XN�]���y�����V؊i'�� �q�d��a�����9�5������3As/�Ӯu����\�Rg���.����I�ɱUAb�P�S䘯�;�d���c<�����>~�Q����F%�eY��h�������O�¨�z�c�X<1���h5�JȜ��k�� XU��;k�S�@�x��F�f7�V��<]L-�jF�i�/x�K-,�m��oG��ݶ��臭g�������B����EIt�j�Z&�9�����\\s(g�9%M��Z�~Mzn�($!���oBͥ�JN>ف���W��?32�ݳz!��|�&�����q�hI5sg���>���E��pO�6�r�D����k�%L&;U� ٵ��=���*{_ܖ��|��f��)o�(V[�t�z��^�q`�\��y/��/Ӑ�uv��yO��f���v�k�C�0���|��Bciw���c
 �t�0ӷ�f �r��,��P�1�����n��f�1�F��*WT�>�kU�[�#���q=���N�?4*��ŹQ���8�h*J�js+B(�mRP+1/�=��$aJ)i�mŔ���O�}����h��X���N�V]4�r �,;bd��?I�����Q;Ƴ�o>T����]��,�:E��zT�����z�n�CIu�Y��s����4[���wkߡ�������2w�k���	Օx�u��}W�XF�:FC[E���s�F0!A�
r�,�`mzO0D�^[.�8\3��h�ѯ�`�0���.��FsR��%�#��/�����~W@�z(勛6��CU����8C�q���i��7�+�E#��������8҇h��P<_�@@�#�A��
�n�S5���ꈫ0V#�4�c���i2��C���rW`������*a�PǺ/��#kL�U������nԓ2*�����r/�-�������1	~���~�kfby��]�Y?��v��A/�.��`֨�@�՟��@%ֽX��*�N�Ϸ�D4Ғ�d� �D���&2��ؓ���-Y� �z�$�x�Ӆ��ώ+�E(:Sk9?:>U��q(;Nu�dW���r�)�x&��c*%�'��ƅ44��o"V<��o �8���)uV���$4�RA2��'�T�n��j�(��P ep^�ٴ�չ�5[^ B��"�!��8a�Id�m2Q�� ��	s�A"6�o7lNX��q[��iTKs&�0�G��+ǳ�"k�(�y5��V��jVIlJ7�k�נdgD�Ȑ�|I+��y��ϧk�P��o?�q��F1���.��.��8>�{�l�B�G�[�cЅc�HQsq?��Z� ��g����U��{����0�M �������5Z�ZBSV2fU�9����Yo��^	���#=��~�%p���u���n�IR���zJ��J�U�<�}ǉ� *m�����2��������H�}���ٛ{�/?�������d�eLc\j��DU	�=�nF�)�7ț(���H�T����^=���4���@X��a�_�$'!�b��I5}g�d� ��w���T��i�F�M��V4L�e����U���0e2ym�H喟,��8�/P)�顒�
/�_Fm����}q���L֚��sEX8@���?HlBb��̔8ڃK���GϏt�n��tk?�&U�8MUZ���mu]7SCT <_��G�VנE>�cw,�#����A��¥��tk/���v)$���R�����St��r_�j�%���� �"IgNn�FE���5Al��W���ˇ2lN*%YZ= ���I��A�m{X���V��i CX����{8�M[���؃qey���^B�D_	Fw���\]�����[�	�WD[E$q0�&���x���������7t Ca�V������˫��[J������_E&y#���H*��V��ˈj�����d#����z�T6\�b�W$6�Q!k5e]k ��n`T����jR�X�AL.��,v�_�����4�Fx�04��*�ar�؆�$3Μ��#J����e�'�ۧ<�vA_��>�{��e�����
Ba@p[�$���\
�Ko�uN�,�����+H҉��-��o�-hf��l"���ɲ�e��5�fA�A�bdD��1$��콀�:�p$^[��D�΁[����Y̙�L��l��&�Xv	��.��ЄU��&����JT
���AW�5R�J��`�q]��@�Nf	$-�M��fZ�>{ƃ�-7�p4�ܨ���QtX�fT7B�L��),n|���5���q���gV�!V���>�=�ܴ��lv�&�)�D�)�Q7E�܈����xh���0]�f�v�K�ߌ�%)(�����R:�[��,]��"v����h�������?� ��)���kН�B�^)/�C%�k�>1�&����M�!}�M��� b��l�r`�G���Q������w�]8ܱ.Ѐ�D\J�����oK7a�� �js���I�$JͲ�o�ҁ�� -��y�c�`�P	�|qR��h�D����@Z���jr7:�{�r�m�=X��ܮS��d^��A�h�^��k	�����{eo駬�13��d��:�%6-���B��у��%�[���	'�g;��N��TMi�
�Tv�v�3���}��
�mK�sP.>j�Fٲ���,`��v�]��~�@���$��M�61�Pc ��7��2�e����@�՜��C��Eh�0B������ v�l0� �L;H���|�,�4����L&O'� ��)�f�'�H>���ܡU���&�
B'�)~H
G]ҦB�����7s?�8*g�1����PU�K�����<I3��R�Im8��wc�Y��2���>h}t��Y� ���M���k]��VF�|�҆nD6�{
�cF�ްk|d,#ԑʀ�}\�xI�K�.��1����쫹d�󆹌F�K}����DO��+	��Km|!�,r?Z�)�D�P�E�
Y�,��)8�% P+�c*򏲅�sq�\����C��?\�Y`/����`�L�f�I-��l͌L�'����BX���'̲�8�&;Ňf���H���I��6a�������zE����ww�?�Y�f�V�nF~��RN�-g�l��S��h��6�<�ւ�`iu|g����M�p$tb�s��ξ��p�c�嗷�Ff���.��wx��rk�]v��>�M�%�y)���BL,h {b���V���Y�io��r�ut�"�\-�攛o�B���7;�6��A!�c�R-��u�>�I�����?�D�-0��c�.�95{�DZ��xnV҄r�������"��W)k�46\ܲ��Mܮf��20�Ξ��P�hCb�2����(��Q����F�nc�6.Zh�;Pݎ9���W� �;��Ľ�5ٺ~Q�}-&�' bpb/b���%@T|=�7�H�J,�%Q�ǜ
Ԑ���UD� �8|3"s}ܓ��Y��5]�e��V[�m�@7@JHi��v&'R�w�T� hvB1k���[�KN���*$�z�7Ÿ�Q	I�g=v�x�3b�H�����A���T��ᷜ�a��M�t�{ ���]z�N[��7��Q���V��[�ًᕋ�\	��tX��Ir�[�e�l-��ԩ�m����-?�Y���S�OAo)�����:��@�;��g���ays��?��FiOZ;{���/����:�9�4X��5_�
�	'z��q��2g���o��w�s� tY���
���~[�%]����6p�9i�m��{t�3�N	U�ۓpu?h�P�G��rlB���&��+���O���Nm���mj�m\?�����s�Br��<t��0�:�N��~V!�l`���I��}9P��1��9��iZV@��R�O�ml$�A ��ѽ[ ҷ�[�˕X,�c&�����BD:y�<g�V�����Mg�;�7\ԏs�>:�?v�o]�x��C癓��ݬP#��Ѱ��):p�a|�������� �����;F&n���_����lҝ�"�UV�*:N+�lKO���Q�=aC��C��������'X�(U�w���0.C�"�rR���WP�B��6z�ՠ�%��Z��n�c�	�tSk6Jk0ż�ҙJ.����3�����8fDtj����z��3�\�E���x`1��ZIx=�NH�ao���+>�i��}�R+Iz��F|4�g�ި���w��I�h����;T�v���B�3[L�9���䑍?�@�RTA�hk��Ӊ�X�&�!_�ESV�]~+?�EKͳB�:�B�>Ą���1qN1U�Ǌ����2\�\?�xuS#BK��;����r��xY�9�q�x7�r�A��MED�R�P�p������JYj� 	a]Ԯ���0U�� ɚG�l���c�� �Ǟ�ݺ����N�Գ�+yZ܏8O��|�q����=N����t�U�f��R~��U�KF�9�3</TW���Q�:4�%�"ܫIw�<i�0�r������7�m+a3����dÄ��r7I$#�@ޤZ�K��Ԇ0N&4 Ie^/Ty��=�N���ں^o�V,D��<��C�T�̯�4u�=�Z�X�NͰ�}k47'}#���ə�!�w[�y]HF��b�J���9�~p�8�G���탹���(�X�"�[~�ǡu94C9�qrT�m�����۩�!(Pu��G`'^u��V�+�<���lo����]͓�}�-�5�nV >����c%IT���v/�r�!V��]�t�k��`�6�@��M>��,iOl�i�U�ȡ
�
%zm�XN��c��[��qu�PR+��t�q��9քe��2~ڒU�s�<P�A�Ro�X��
$�9��^��sMvL��{�Wt��ɸ�;-�)��7l����~H8t+޿yd�\)tk.BƨK��̮�E�,���,����b���(q�#���Ώg5��?v�F��0�Z�[Ò)�ծ���?��7(���'
��c���}�+	��k^�*�C%ͅ=�E5�ϯ���'῍�D�*8W��y�>�D�������w+�Ɛz�{n$�>����(*w.��@"�q��0SZb6R�w&����ݭ�k
�e/]�������>v�p�Jq�32{?�9�!!�
��C}Q������u�F�_�%,��P?����׼2>��{ٍ��?�q���y�!�h�����1(�&�~1E�����k��l\Y"����<�)n���]��0��v>���S6t9�<�ן]��B�ӳq��b�z�\�H:��);Z��4Bk����b)�t�����[]v#ԠaJA��l�yFR�S�6��jk��ar
 �"^%n��Ɓ�i(� ��ȏ͡뭷���D'�N�ڏ��Q��`g�F~�i&�Q^�0��?3Y�M3�h�q�1Z3��WG\�~jgl���!P��֯��'
qf:x���x��)���Z� ��i{�М����:+>�K��u��r��2��0�WeVc���2��`�����@<3Ll��uv����'���/y��_���H�v�@<_g��g�� ��w�LG�FG���M���!�*�6y�?�����i5=�Eof9"�K1P~ޖMɨ��j�u�H[v���*:9���M�/~�\0�R��-|��/]X�-��q����sy���(&�)�EY#���D�o�`[�\����F
@\`���̲���G�R�� |��0��TUi�O��L2�h�@jk�����2�J��> H��F�*�'��&�MEDӒ�m���GX>�d������p|/$zf4�B����(�*��q�4"��Eg,�,��+��� H����.���:��B}S���Ⱦm��U%M��ro<t�P�u��l3E�e�ڒa��	��a�M3�L�TJ�;ә�'���Gx9�-W-���pF�I�|{{�`�>��dY�!�0\�pqba�ͫc�گ@��X�7m��M��MLR'�	��ƅ�_Q���l0S�}���\_���G=�'��<��6o�h��VL,���S�
BZw{���D�w�DT���Z�r�l����8��Yx�t|�����^`g7�����b��쩕3<XA�c�/�)ej�v������/�yd@�q��xIκ>��l_�m����x��߉n���=uh&�v�鳠�&���o`B��C�q&^���!��3.�}�(����h+Aw�z��}Q�R���=7-#�tY�awc1N�EV+�ޫ�Ѵ,B�ћP(� ELZ7\ �eHJ`irh����&:4�SKC���}G2��c�&$?I����*p��<����:!�u�jя��%�t��?Y�vh�	�*����ǽ�L�$�Ѡa6u8MúD@�E�����v�z4�a�!������1
U�dz�!����e(}������9]I?���i#K�a�	��.����7Y�Q��e!5~�O��\ќsI��H/�`v���z�7�H���=dƨ?C�Mf��؊D������2d�4o��X�a��`5Q?bF�޴1�X����Dӷ��6�pxj��G�iW�߇(҅r��o����*ud��6(uP-u��$��r�if'\��ٓߺ���V`�cn�s����/��,����v�B�Ġy̊6�����	N1��h�u|+53���B��cc�(����:����YiU���n~)�b7�1����	F�HR���o�^#z�H�1m;fv,ֵ��K$�)64N:c2i&��\��̧7w�8Z9!�^0��!;��]���F`0�4���`�	 Y�g{�m[ hTaEXc�D�	����*qf��'����DgGR�u�1F=*�r)�����P��v����~�$���j�%g�=2F:*'��j�4W���oM����Vv~	�1�Ѕ�"���Kk��|�::�n��U���ܢJ\��Y���[�\_ ����-�������XHU?�v�1�S�X�-������:+2��)E^��ɒt�����������N�K!z��y���#�E殐��8�׃��ޙ�����`�[���';�=S� �O2oP ���>�&W��ޣE��"��d�("�Z�7����4��V�F�������Ќ����]���ecM��r��>+s��R��#ag�Z>Z�F)ܘ���r����ژYZT�z��y�V�{qZ}��U�4N� ����&�'�}{aޒ[�|�ob�ubL,�;-)�ʬ&zGT��U�J�0� �����K"/Gut/v�ܩ�)d��
NE� ��KT���t�2>��{P�s��,J[�5֦DE��8|]ǋ�/��C���m|9V��9��;�~|��K�2�?�	6�a�׸����?�bQ/ܣ�fC`^��u���z=��ʬ2(Tǳ��c񎠩\�%�d-5�Z�!z���*ٽ�λ��Y�pWq��ز�z��"~����8��f��:�7�HVfv��U�����G��}�ݚ:��P_�j�G(	��&J(p g��yT%�z[|F��^+nGtk\9g,�.��s�HK\N�����G��3���i��j��Ue�hOf���`�`n����/�>i�<ً��b��	U�r���93�/�Gu�ѳ����d�N���+�e�j,�H1�[g��^.K=B2�L�ӴeRs���k|�?�����ϰBo�<'-Ph�Hb_�K�����d��Uiڣ#v��)|FW�l�]�p[���v�'���
�g��B��d7�(lBR�o\����Ͼu��x��6L$��f��}3D�Br���t�F�N]"k`����b�t`�����3�d��I�p�R�Ɗu1����,��\G�O@�TЋ�^�#������>����fx7k�Q�%6�&Wu�%�[�K.��&�`^�g�Wq,	~-�ۇؒTI]ݼg�V:1>���[y*3t
�w�艘VRBcu��@�Z�$aW*]��j���]脋��%b$���r�;��O�:�Hl	�+��<T.}F�����WI!�$���T����T��޿@�fY��u��M h��djN�g����K2^$��0�X�U��?�݄&ne&�l_�]�9J,	�qW�c(�{���T��%�'q|"�|W#��!BE�-�gOU�CR�o�;��w��R^����;��(UG1y<�wR�H�C�,�q�ќJnX���.Kc)P����U�伔�أT4��5z�߲V
�{Kی<�Q��Pk�s�~aY=s�eZU:.�%�_)�~�;pL��ȶ��'^�)�yk�������'�9�F���ۡ�)�]j���U�V}JI����Ŭ�M�*ʄˌЗ:g��F�Vg�8���<�)�}3� j�>�����x�yU?C�Nc"J�Q������3Bo�GLf����X�K���4�<!���J�y]nN��!:Q�[p����}�!P��@^4���.�ܽ�.W�S2�r��S"��}Wut�(�ҧ}*9L<,���J�\-����5�t�[g�g������9^2GY0��Ba�QE׶2�|����zi[�hO�9#����l-9(�n�1�^b�l0����v]���J��~9�{��hT\����T%��x�~m�D�T����/�i�BǳC�|&b�b~��{�6�j{�*�z��;�p8����W 쌔�	d���GB+�Aޟ���@�͇(��<xp�K���Ԅ@8�d˞��WYCS�zzF��{^����ڈ2+�fG7i;z���
7fN7��w�Մgר����!�_�(��� �!�#��Y6�鏶��R��HUj�3��I|�' �2�� �PLʳ'G,�&��7_-���b?�B^�b7.:6i�tPCTIw8/͡ԍ<Χ�ؾz4�b|>�T�	�K��=@\��
�t�n0!�}�Z=�g�.i��Ǿ���e1bWۿ�@���ڡ��*���[��ӆ�xSE����"�t��0.����nh-a�PK}�yk?�Q�j�}
"��1t�������O�!F&��o�=Xy֜-T�m�)M8l\^����j��`�0��<��4ad�+\��%����dЯ��3P�-�#�'	%6��d`ʚL� A.�~0��kD�`�E�6!�\����~J��sLֹ���-��pvҭp�m��K_��E��}X�[A��pQ���U(u�2�M�G�1)�UAM?!�P�=���n�������E1�c�/��/��XY��役Ý(+6CܔS� ���u>�a*�WA�ӻ6��.�������`䞸�+I�GhD.�u�yж�� Y*��9�ٳXn���kg�dJ�>�^3	�î�He�C~@�gK��85�g�J��(h������M��ii�%��E���+��Rdp�W�7�w��52}%hU��L�Ŧ-��;800�$��8�d�rQ�*�8����hݴ�p�(NG��د�$�r�Dd~�Zz�VLwӍ�2���;"�}�a����(���X�_������﬚r��A
�T@�]L}����1S���A�@�e�m�-�ǝ�\�s?�7�[�o�D�^�3@�c}�CW:,c�r�M����;�N�W:��~J�Փ������v��e��/��`\|l�Ϸ<��F_`��f=���aPo�Ӎ�F`H�X���{���'��iWg1i{� ���8�!ako]�>\��GL�x����!�Wi�J�{�l�Z��TP�^�͠��LKt\���z��E�����#(�ȉ��|h��S���*�=�*X�/�E�t��l��?j�ٵ�l������xulK(��-1�:�πz4A�QC>VcbLwA��%�?��mM}虄5M�Q����W\�IT�n���&�8�uٷ\����l.��Xd|�La�LGK�Q6��˝�t+���߁��aS&)_J�~Ʋ`ks6����_i��������+��S :�y�>\�l�?��G�X�2>w�ߴqt]w�2�F@��Q�y^��%y�d�=
S��J?b�yn ������b_�uֶ`� ����'[VbV��R�@.��X����Ě)��=��\�б�R�J�&�h
%ܵ�����Ka&�f0P��ܧ͞����\��;l�`�����`���`����r���1����/�fLQz$��,��ZDr�����)l�W�����W�w㑣p49�G�(@)���)��DVj�&R��s���ّ����0���})�@Fd�%"�av�.^f;V��rݤB�5�	�ME&]�l��0���J;) �p׫c������__H��6�' �g���m���fI�n�v��
�`S.��Uu��9��	0�WL/=B�:2e<F�1��,EQU4f�<p��N3"�U�i_�x�J��V��Л�ʻ7��-.��0����l^��%�Y�s�8˚mE�j;�VA-O�a%��d@��=3�+K�u�O ,is�ɺD ���Z{d��c�K�\��)���?8�<p�=� ��+\�?��hɷ�a�291[����:�H���O�K<t�����\2�j�c���}�k�G?��Y�)غ�?���Z��M� �~F�������&����:~��1�b
�J��%V���{F�a�jܭ�ݶԭ�l���@�����j��8ցaM��Ao���US�`�S+�� ��`���a[�A���9�Чr��2טP������j���9BM�A����-�C]�k���u	��Lf�f�Qr��̄|��Ďd5�:���Ʊ�}���{Fl(��A��O�3�hB}f�J��7�2C&ɇ�]Bu�: &��h�x���_�ð�f~�]N<	�t2ڒ$�s��vL��7��23ͬ�e�(�� ��6�gJ�:�_~1�ؿ,��&$č"'v8�i�R��5�P*O����O���eր��C[^)<��V��Sbj�}J�5��թ��!T!�A,d?��� �*We3�\&#��3]���UՋ簑	m��ř�N�ںM��j��յ�zz��|T%���Ud��ū/��2�-���������Ī����.�h�j_1	���o����uň[W1`c8K(cO�u��NuqSV�YF��3v�|�]i�E��|@�m9L*��*ADP<+�yX�U�9�	�]}��F��X?���@f0<2���W��ge�}�&g�ZД����$>?�\�l%;v[P�e�h�aŉ8�"0ʫ\�_��ɻ��8��:�Jn�%��`�X��\5�=pt�ĥ'��,����B6��������q�~�C��q%��%Vh�NX�����/��.Y�N)F;	9#*��=�5u�Q�>��rJT��D�u2�9�S�1l��p��MӑbDܽq���=(�s��8�)Qe��0�'h�cY<8.�݈����2�桐Cɳ�b��ސ��a�+X=&�_40�&��u
� ��F���S�}���B@B��J�?Q�����^X��]C�;�f\����\)���Ց��R�w�ol��Y��6+�����VY�;Ա.Ɨ�-'[�����N��g_$,�_�j��[B���}���C۹�jr�����D�K���<���{��9Po��V�v�a��?�c�t;��7)����m����<9u����:Z�'�To��TɭWg�m��+��Z�i�=�-�d�WF���H3�&�0V�R#��\T��v����~y�*IM[�CmB\N����Khf%!�Uý��dBtG8ֆ�l�r�2l/0��Nߦp��H���o<��,7����cL��(�> ����k��]c��T%�8�@�t/�19N4�E�pM+��4E(�)��;/��o�lL�F/�\771�0�V
t�t�����>��g3.�	$c�%\S�~���G�a���5���ѣQp$�d&�_���о��|��*#�����K7d���p{B&���߭�ȥqUZ���)i��k�yla
���J̽(��S`#�T}���9�u*O*ޭoEb�aғ����B��c�f��7�8�c���Z�s��){���+����/P��]11����ir�V����BS1܉ĉ}�XJa���CFǳ��Dc_�)�X%�'�-�����a�A���8�q������Ь-���4�*TS|���7��%w��z��)�Ƶ`��i4H�My�K9*YD$��zF��l�M=��u'3��A�0k`,�,*��.��S����O=����7�v���j5 +�1{U�W/���+�6����t��UY+V�����\�� ��-˒�sAB#	-�A��!���YI��.B�i����O����+�O}���G�����F��f��O�2��8�8�ئ���E�+;xϬ�5��}�;��񗭡�؉\�H�	�ʳA�"�ΛZG��
^�ih*W��w����_6m�.�����v,@TG���S��:�L��Λ��$���[ӮM�����ze�Eg�d��A�Y�^�3�WH���65ׂv%.�#柈��xR~ˇ�0.���KGݦ�vqSm�V��մ(�t��쟵g�n��&��h y���ٞ�	Fm.� I���%K�e�(l�Dm��R)�8�䊺_�c���@m��#�H��}��_N��"�4[vs.*;�s����%ͳY0�x�2{��<�L�N_ʄ�{R	�@�-/��`�I�{K���_ ��ҋ�h��&�c��\m���d@>���4�0=�w�p�{�T���� �� H@:�\]3]�/�k=BeR�������+����fH�6+U',��׵	jp_AhqT��7|8Q�+{[H��-���j�}�c
��<�s�`��a'�}�L�9�m|��Ff�w�D]� ��+On�ܯ3���d���JO���V�w���f�}���<9�s8sc���qZ���+�Fc�7�C�@����/�C���� ��F��!>�l3M>\_k����@G�MR1�����ѓ��"O~��%�f�'���4�Q|錰'�ܰb��σ%{"wk	EwX��C�Nӱ��a��=�;�M0�i�h&c	���Sjئ�� y�a}���x�
јJ	K]Kh��]��k�K!ES��P���+2D㧖�'�[�Q�Xk9Lb2 ���(��Xe5 N���<��(�`����4��P%�#�6�a��NB
JH�� Q2����	ۂ��ȇ5)~�R:-2�o��4�\�W��mJ�:��y���u�^\���������q��Ёz-c>5R��L]v��i�.�s���D��򡅝;��k���伱�d��n�SZʞR�Q�j���̇�0]T��ڥj]>		���τ|�{zI�%ŧ���a'���F����"F�k5��J��Tf�o��?�4"��=�4!C]���$����żۇ����<H�&`�~���+�F�X]��n�{��Ɖ���F�Cυ��<��_y���bĐ�p{���������N#ϥ�O�]�2�$ ���^C���(52��> �i�����R7�k �4��C��ӦD��uҎ�A.\�K�s�]���KJ�?����q�Զ�����
C���:�Z��JM� 9m�V/����)���m��%�G`��ǝ�f�<����
}C(ݘ�xH��7���H�if>��yv�E��|��q�f˒���_�����c���iZ	Fё�$��ZyĎs��
�ˮ�(�`�oux���̯��l�=u�/ ��0ڍ��e����n0��_X�X��5 ̨$aG��
���"]x�Zq0ff���*k�$�oݧ� ޼��7̕U /92��b���iu�)�F�*3�o���Y��bNj�}C)�����_���L�s�~�# w�]D�t�\C����>�ģ���p<@
��-A=[K�(�KZO�5)�/���	���|'�7�9���Q�q��H^��Fp��$�����dc��*������ה�6d�{�)5��z�90�.#p���2ՑU#�#�R�l��!n%�[iÇ�v ����g��"�J9X�P<�?�¦����Gi�DL�NS�g�7�����R�stb�JM ��z��Es~0��[7�H�1UQ��<���d�-}l9Vd�D+~L4I�Mړ����b�A�#t�����丝�
��<t�1��Gg��}|��)=�m-�� �ŏ����䈔��-����Cj��3�����F/�� H�v���Y}g���o �y�����z���S_@�l.��W[eRv5���I�G��J���܊�1������y*W��6�+)��L�?�r�!sI`�����ݻ&3�k#��	#��	呏ʄ�ۍ=@K�p������b�a�u����5\��q~��+��~�ͨ��LS��(r�Sܔ�aΗ����XԨ�7'��N�tg���RH�e]��U2�pd��D��!U%p���,�0ߩ9��4j.5�&`����c�n�Hd�������;�[R��g��<�������=0擌�@YxH����x啍��0A�4��v�<�y���	���Ί�C���G��8t!�A��a2j2C}�3c;GZ5�h)��jC`-���4BnM��E$뀥��B�f���0@=�ح�T�y�WFdֈB����-��8`ki��_�2oFM�����:I��88@��D #�5������a-��O�M�}nl�;*��ǩ}Y�J�Kĥђ.�����G��T� ~$��������E��m�5�F�q.�?@�o��%�ggX>���\,'{�V5N|�$c�gf>k~Ԝ�cEۡiEC������ �A ��aȯ��y��fV�#���O�4����e܏��Vo��*sm|R���:0,u_�F|�5q�r�^;!����F�j�S��)�;mO����3��ߏ����ϑ�ܓ:��A�T�>�6����֦0_�0�.6��;f�4羡���*G��٢���;^ְ�&r��@���ޗlU�仛*щ�g���v4���a�a.G@ط_�8�N�adӶ[�L�o��?�7[`��cK:�
R
����j;4J��#��X�]6~D�`P^��Z�}>9aMH�������I��v͎�-�%R�)�#�⑝�x���[�^�F�WB_; �a�H������}	ǳ��cƔ���8�E�Ang0~.��F��y���[f�եh���.�ji�B�cJFP����_���hHJ�Ѹ�d�5�,`"La�%���T��[x`�ax!A�z�E�")e
���C��R������E�Fe�q�
��w�kN���?�x \����\)F�yFȹ���҅sOA��8���ͼ�V�%�X��/�)E�E$�� �� �:��rs76� �g�b�hĲ�U�{g�GS��!�.�����Yb����
z�dL�$O�qU>��c7��h���J�KE��?����ǲ:�LK{������?��KˑV��PxOk|k����Axɉ߾��V��|����4��2�jo�3����'@�l��,Q-���bn3ޒ	/�@SZ���љ%;4��V�
���5��~�ai\��n���R��� ��ʡ�wU]:é�CW�K�}0�!xw磲:%�ڟ����~.���(�\�@o, ��*�^�p[8<o��/+�b�ɄSnh_{�'��a���R�E {,-��
o�$s lR�$m~��Zs	u���q���w3�mܸt*-$�r��
ڸ���G"�o��]�HZ��=�q���b=$�L���(S8���Ԣ��$�v��|���=���!�+���["�`ч2]�3[�т*_w�h�f?�!�]TW+7,��Nռu2�-L�И���\�����0��j�� ;~^b��^�F-���2�Қ��oa�����0f	�߹F,2Ìm\��հ�|7��1�m��pC5:7�ӣΏ����q�Nڢc�@#ab��!���<CA_ɧ|ټ �O����zF27/�+�/MZv���L��2}���+%,KB.�(]v�@�}������3�h:E�ڴ�>����ԟ�(�#:H�U�c�\G0Q�E�Q,��Z��v� ��-�Bc�0���4wy'>a��W���ɸ��3%SN����)�����W�^ߍ\�ڱ���3�yaki�[B������S_-O��F^�E�atW�S���[�˟!rUE�&��w/Ē����^��i��y���VN����ͪ�Bv"7e���sp�O]�xyBt��>�z�.l�ڪ�y�V�a�������m�59c��`����VPl�!����l�)"�IcR�hY���:�6��\� �c�l��]�M׭�T��5�W/7l��[��0�������������-��%���H��X�
wK�Ѻe�R�a�&+P���O7���岬�v�5�"B��mUp#ۻ�+{W\vǫ�?�
VpY�S@ǈ�/��aw��.Z�ND���fq�22��q�M�s���0��~�����Lcv�Ռ�Rc6�ʄ�;��ZE�~���h��4�&-��i��� ��&k.��z[ 5��V���"O�$�P��h?M���u��$Nc�e��ls���$S�g2�j��3Kx��4*n�YY�o�������g�����O���3�ECK�A	X�?�T3\xΖ�39,ve�5}pK7��B��� \}UQ��ò�]]nC��B�F�	4i�"}�E�Ui�=�l@����a����L4�8�N��~=����q[1F�>y�1;�^��	�Ɛ+��zr�����<�=d�1(�qh�m7X0��P�0dj�$Se3�-��e<_֬�qqPH����1�,�|zЂ 8��Q/��˦�r��-�avɸS>�1�͜��H�|ˈ��Ǉߝ*}�c�?̚�Ş��a\�G�D[��t��X�H���>�ɺ]|�j��ﺝ@X5a���ٶ�k�Z�l_�Ui��i兔���T�c�lb�K�ߚ�)��'AQ6�$����N�-^H���Y�u�+si����K�~�Zk�<L�3P�v[-~�l����|��1�V|t/	�F9�����ﭤ��0�ښ�i��w��2�Lū�g��wq�ƙp*��}TDw�A�ʖ�Մ`�g��'-�pt�0��R�*~� �fϕ4��J��TΉ�u�m&�d��F��B&��
g5QY)?��O�Z��E�w�>�M��rG��er�e^D�+%�.[C��3
��A�el}����5�*�\o2�����Lwz�p{H&.IO=	%M>>xF��&�¯E���J�����"@

�H�65�ǻ3q:�ah7a-lpc�ݮ�LU����hN�ؓ�t��j�� S��2�H~�36�Uc+�:��[^�C�0!����8)�,�b�	|��q�b)R}�zې�)i���)j%�M�u��BR�ʔ^���H�)�$�Y�M�ݗu�EpC��O��[O�jZy��W�l@�fY8!�?��~
��n;�f��js���l�	�����́�:�n��33����+7���}r�z�7�J�y��s���S����6]~�w��w�w��r&Ϳ�(��+�ś�g��͖�Z~k�D8�����TM���?|.��ToM�o�/c�th�-��)Չ�+����/�b7�-�S*��~<�MO�"���PE�
4J���G᥮UmU9����𲛒8Ž��x�	��/���f�53�
�N<�v�id���V�}����|TDx�����i���S%O� �������S�˺;�ܒ�Iܴ@þ�8Z9�O��%96���9:�v�)��ӿ�c�d}_���|:R0D�Pk��ޢ&d�%�tSY[I6�KT:*�[G'oÍ�D�l���4���3�Z��b(�k):2r��L��H�,	?����L��aj�8�|/��FWQ�u�![b�fTip�ϷPL
��ݿ�(�>�_S� BD�I��uP�g��rX|��z�?���-���P��("�D�5W�#��-�W�6)���]�$@�Y&����ˠ:.���Z��Y�� n�B�]�ht`z/܉h�
�s���Ԑ%e⤕lbagOw뢷��0��ny��M#��Y��Yf�/s��i�Y|s����]�:��1�\���ɨ�S�g��^��n��_��4OC�����vc��4i��wI`�u��7���prb� ��H�Y��d�;��S]iy�T,�G�a���d��-�M���j2&����s<&��e�c~���C�Y[��\�M��|�[�� �5h����\����W*��͞ �����6�A8%3^�QM��E뗱�������Z�J/n"����>�~�-�dM�<_���v���fv΄)��g������
QY�����u����o:�C�͒F\/�
t
��㨔|�<���@j�_\�0�#+�Շ�>�sO��%�hW�u�g�j��`v��e���hȉ���b�]B��s0!#��2�xj�J+=/C.���N2"�=��ʤ�>�}7c����|���∩���u�$�dlsJ��,
BCį��yCGb[�ۓ�?�;,�H��et����Nkf^�L�B�sAm\�9�v�%�,&����R�DtNpd%A������f���甝���Vkɤ�`��0��"ˍi�����AN��'�k8��(>[�}�edc��>;;�G���b���2yѦ���){�4�]�|�]��F�9K��!��X��s�T��&!���A�=F�$�`�0x	V���3�N��hZ$����Ə՚D�k-�4[��3!|�sHسUD�4�I����4����/�!-�M)F���LH�/)�Ǥ�^v"
W,QJ��H�����N�,%g�^�P�|}�9��fkSh#�C�𝕰�7�k� Z�G(4��+6
��w�e;m{�u6E�M���:;wH���󻷉��^h'1L�]�W����ەf1����GU V�m��Z�C��J��e�.���LM"��Z�b";���ל(H�I��v:e�S:m���[�����r�H%o��vN�߾�� ��q1]-���8����ݷFhY��WK[%���?�b�J�JT]�I�t���K�'��v���<هW�n[+X/{@�6�ɬ恬��a��j4�2fo���}�OD>�֝�:�4G��e� /�~���U�-��ٶG��y��,�ʢ5](� R�Z��@Y��y��_�F)�9#���<��̚��fL�^��x�}�U۴5z����v�G���n�����,(�Gx�7(/��
���j���{���ɝ��K��-��_Ө߄L�ywh�[-)�ߍJFr�[D��a5���z��}T-atŗ��5)�ҩ�K���ǚ%�qL?��6�`j��׏�@���t9�m`h-k��Ư&t�$�Z�=E-W�b A�^���-�Ytv���Z��wxz^�E4ȳ��O�k�%Xn�آ ���g4��Sb�C�e#�AY�B�uyi�!m���n��r�+�x�'t�4�%���琝`N׎9�o������p�{ͨN���-�����9I%�FQ����Y<�囎�dd��Zϗ�T2�~-(PsV�s�.�����%��e��F�G��<g�+f��F���8;!�\�EW�FLn�y�����	�'�`1_+!~�|	��dV���IJ�vA���a\UsxҘ��}d���ș���~g�g�̛�U��[6����G.ۢ��vk�`��t]u:j�$HgI�Q~V�)�*��_���G%Y&K"Ӎ�Cc�6��v!�a��ʵ"&�1���=��Y��e�
��y�����������'�.�$���Є�%u���x/�̟�R�V/V�D\U�$U@�k�Ƶ�����{>�F�d���#�����#|%��Y���U\mW���3Ty5��}����X+�t�w�<���7k$�Vt�X��5��`]2�?�c��wh�l�wks��*��Q�%�0AV�`���h��<0��8R=]�-�F�I,��� �@Pa���Y�"P�ic_�ʥ)W�2�`t�h?��Ȯ�-�?N�3�TA�3�w6�����]^�@�c�+�B�@W�t4��Tzx�����}wܠt��WK|wksm�����c�K�J ��}�kr����tVZ�2��U�sJc�+1ا,y��q?S]�k�� #�����4j�v�o4���� �U�_��i���6A E��G{����9E�aP�܂�kF�	��G$���&嚜$�w�3l����q��Y1�����?*�P���'$ʣ/�2[�7�f̕B����e�T�(>'ljF�e�5�h�\G�L���4�<0��n�îC)������u�F�[A�K,�:��&6�ւ-��,U���<�����L�7�\(�oj蝣''��%~���۴&l��+|h��P�#I�@5�����ց1���X��睇�4��j�&m��ͧnK�	�?�<⩹G�f���~��1��
��͔C.|��u���ӵ=��AGa%��@è[ޜB5*���l�>��$Co��Q5��yߓ�̵���'ʉ+2��jH�C�r)N�*W����y4r�fu7�c��<�e�`WO=
�ק;���W��X/:b�טӑAm����s�7`z�ҙj�]FbW�׃&Wegb�ܭ�X<V�Z��YC~���\ ܎(�0���g�S`b�J\Mr:x�I��|5yQx�����KO�������'�������z����pYXI��h� cO�Ycǣ��h�̵�:Q�+�������@w�S��݈2��]���OM-�L��kd�AŰ�4Bz�7A��YRW��V�*H�"�D�oY�q�V���c�B����;���N̈�@H�l,���f� �(FPD�Ɂ�����q�v�m8��qze�ܓ80�����c�>��tX���Y��-4XnD�6~L���Wjv�����]l#��6
�60�z��M>e�6�;�t[B&<��_c�;Fe*փ.�ԡ)�EdFs���"b���|�*��~�4f^X2�nawv�$�bzD�)Xt��ݝ-�!Gz��B!,b��u߶*�+��Q7�Y�x�N������r#�g��p�y��!a=�K��+�<��w�<��}.�q�TWhw3��MYN�`~m�0��VC�4Rt}4d�r�G���s�E:'!���2��~���,��L�6�2�0l�w?+�a��S�cREj(�v���H�aː<�B��(_�rQNHͅ��h3y�XÂ��������pr�,4'�
,����u��\�Hε��מ�Ln��k0[$6���c쟬T���sυ#JY��J���As%e-Ι"�B�]T�'v�X���e�W8����y�א'�*�v�h�0	Y5U����<_3㽵	�x����>�&��3��]��v���nI���DS��Ei*Z'�*�k#�o�N\A�h6J�WK�����x�c��೮t@��3��&>���RI"��hO�kRL�.�vJڋX�Pn�'�Zx,	=1L�3��˟V{t{Ҧߦ-`�4}R��[uS+G��J݇�8Av�)x(����C,&a`/��I�I���<uer�N.8�^��~іGX�0�,����3B2h(c��l�{	^�R޵��@��KO"�;K�@ӹI�`~����Fb�|��U%W8l����C�+7u�6$_�����ҹ����t6Z��y��Œ�:�{]��H�i~o @m3lk	\&:��s}�!���CNLs���������M?�H]#��Q��t�� >ܢ�3\#��\��4$�*�E'Յ֙��v.Ym{��,�mݟ�:�e��V��D�����f ݫf��a�50nV�����=���Ȫ�j�hH�}����K�k�s�Z�"��]�T�'�[k�\���kk���pD�c�mȞu���ov��=:}DO0�����ӓ�oͣ$-D�M��Y���})[5=L��P��%}T>�z��N1����aI���odSya�Ʊ-�7��_6�k:�$��]�3�{��*xb{�!9����]%Mi��(�U40�?��|p��,h�+�m���� /���VgX�����v���!�DyU�h���*��[�@�L�NV�u�imz�ƔjŖ�d�� �����B�[����S�[*16�s��B�S_
�%Rh��˼�4�K5�3�,[�ċ��(ϮZʐC4��A����md�&CB2цG��*�\�\�Kf��z� �=���2�T/=��5P�j������9ɥ�l���#7�+B��G@�N�t�2�I��|�,VD?�F��Vk��o%�"�e����.u���bF�.5mk����^Eȼ)4J<}��rRZ�7"�.ܘ�E���G�w	!eE����J pz��,MBMئ�y�k�ϩ�����Oi�=�nǏYj]�M�V̐�f�F��~�p�����UG�y���]e��|��eQ����+&���M"�gZ���E3mQ���K?@���P�W��ߚ�+?����u�;
q^��;�CgŌ�qio1�I�&q��xX��yzߠ�*f�����ο*:h5s_g���qp��]�X�˳BvHZx�s�q�a�x3 ګQ�	�q�o�B�L,�T���"-�<�Pl�]:�l��Vh40~��I6�o�O:����p����jH���'�~�_��lkP�k�ub��s���M����{C���B+�+_��B_v#�	W�m��wb�3���[H0�a����Š��9�����v�NQ��s0��n
c��{��Uv�Og1�"�@?n�]�q��)��-ě��t�
"Ѧ��c�Z��<AW�ғG?1���,�����܉
b��������W�o�����&c�Y*���%4+�>莠�a�̔$���_�~��#KA;X���[|��D����E b�/"�/��i��iiO1��[�cb�I-!cg�}f����a��f�c��*�V@�3�P�w�(5��Z{���/F'��Ԓӓ�D=$	�C�̱@���M��̬۹�ܿ�;����yt:m�� ��>J�I���A"���@ȕ�S�&a�G��*ނ��)M�����/��'��]�ގ<T\�yk/�6-(�}s���hݐ�.-1!����+�6��=0MxAJX�SWL��׉B���׊�����Q����	e��_�X��u���i���?��G��bT��Q��7Y��c���Yh�/��v(��F���n5�B+̷m"�p5�&��Q��ġr��\�Z���d���#�3��N"D\�nXm�dޅV�s��/Pr��SAm�e����1�t	�OJ� W��@�����P-���Y����(��" g[���٣����;���и�ɡn�/����6� �Cv������3`ך�w;  -@M�,}�����lK��~�߭�D��T��ǌ��fx�M��yl�\p����>%��es(��U�� �>'�_[��m~@�����+�>7s�!�~V(�v�|���~���B�;� )"��=|�ͫV$�B��0�p��γPR��!6��I��c̆��b����TcU%��nt"�a��FD�,q�����x��Љ�	5E;��L��M�NX�B���� "lB��� ��a���g��1�o�/��4���*L��@�/5A����
a=��i�ci�5����"#)�Ę�q{��Pa���)��"�QP�ʸ��x=$����~>hj�q�|�R���FG��t����򏴻���w��x?���܋�|f���vV�3�3t����h�A!g�!b��^$��ਫ਼.(q'?���mn�O�G�7�k@v�y�;��P;TH�e�4�3�*z�����y�,F��wS-�f���$hR�9�3S=!��ſS#��_Ȝ������@=q���aL�
9���ܓ�A�ǂ](!"��|Vt�8�9�\����H�χ?'#p;`h�p�	��xd�ug��y��*I;�vg>�
;8�L3#�]b��c6_��+���D5��1X-8ƌ�w �j3 �%J!Z�����^H�l/�w�N��D2 �wc��y*��Ǝ�x\]1��b�
ol�9�]��)�����48�E�O��Fu�rjy�;��^2-�6�*0�.B瓐P�Բԝ�#!���Ͳ�[�]8��pYI�D,�%� J���/)HrL2r(˽~'�֚ZH�
}.��FC������t}42=P��i�׊��~��n��ٰ�zG>�ѷ�9�o�גV����Uv���oZ*ta����j�U;I���(`�Gjto�����#�^�ko�Zl�ҡ�1�O�D7þ�!N�㲉Ӹ��J�oC.0gqKk�v��ǋe�� �vu�����c.�%r:��,��,���x�c�K�C�| �o�Z�fOG|��I|�y 3SqA*�@�;ω���+��J&��Rz����%�2�.{��`uO��~(�C�kHl��s$�S�驕��c �����3ӽxP�p��`ലB�ܹx��[#�#k6t1v��'^����ͯ�� �(�$���]���K�`��#��Ǩ�U�@/��[>�ܜR�����l->�G	����ɇBFkβ��J�}�m6��	��� ��3�<nضkPݔI��%u^pPKp}_D�ͺ��%�� �H}��j)�*[�l���}U�/$�;�4�.�H�K̃��������q,���S��e�<*ſ�?���q�c =���L���`~jO?RGH����7�S�mR?e�.b{�6��Ȯ�mr/��������5��]��w����`���z4�2���̂�Bx��W'lz��ؼ��D@*��l���kːh)-���"
�'a��m팒 �u�F��CՐ޲�];+��~z���<�Eu
`
��3P�x�\�a�-�����I��n�IY*��s��Iw�T�J$N6	 �p�~�ߑq�?�p@��rI��&ԝ�R�qƤ���e��y����zzy�� n-�����-�̹Ů���ݡ8B<-!��gQ��%�>�s� [��gc ��ʯT�U%�kn$@!pĶj��v���c�Yj2���_d ����w{��j��~؋�@=��]Ɩ*r�ػ�p���G�+ą�"�/ߚ��3���d_���|�;-iE���R��"�i�s�����Wٲhc�f�õ%i,����v�$�K�O�*�����!�(>����of��.��J+cˑk�(D�6 ��[[��B>��-tm��#똾� �=� r�����0��K��]�|۪	B�S�:.��}��\�ȶT�f�]����|�י��d��ˁ3��z�������;.=i��k��V_ԝ���|!�AG�ɕƮ���ޓ�-��
Eҿ5��g�K9腅F���N�.��Q�q#�����\��w��,�C����r$��t̡O�x�:�c��8g9���6��b^�����	�Ⱦf�d��W_�WM�i�<����i�f5zmW�����:c���&=a{(_R b��:�>��$�7�P����y�\z��W�>Myut�N�ClN��p<�����^ǘĴ ��=��)�A�y8�U��2�Z����:�4��ۤ�\n��a47��J<��ٟ��h@�������WތLh��0�H2���(���Y=A�v�h�F�.��\�K��!���l��;S����7_5Q7�����i�z�6ɼ�<���5�r;ҧN���;`;1N%z��í.Ot�(�hN��	��]��f|۳��hwp�L���M�p��F�����o�B�k�x��,ILg%Zy�̇�_��`�㹇٤�p��vM����
�Őqr:��q�@��o��LCϨ��5�;��;�p'*��.������2v޶���S9ڿ�yRt*l��@D�-�ؓ���s
��V]���{y��+��1$��٤2)�F�i��8�
ヌ ϟ�*�7�K���%4�,��`V-X�m�m\s�!����ٛ���u�3��^�[mcC�c~kgU�I�^�a~�m��T�A�2������hRQ'<X���<{���e�b6�P��U��-�#����s�08b�oh?~�8�bSƀ�je\�r�2
I�޳w,/3يS �@��ϖ[Hq�h����I����dh�n�qL%6`�^P�cV�� ӥD�K�ob��ꄺ��/�HAߧS�w�G�esb3$h��c��c�DE��9�R^�z�	�nyYH�%
�}�IG��6�"�+���'����o���ț��p栋W��	%����̑]�$W���5]t��8JDG�9�E%>��{l|����\UA�N�Ƥ?a�-��'4���uK���0�ToMM'������ؘ�%�pX(�Dx���#���P��Nj1`	�ْg&�>,I�m|���/�V��$�v|�X9Ą��N��vuc
]F7�&8�)p`��yG'�C��U�"f��rm�v?`ieaB�f��>��P���CF�E�~�@͜#�9��ho�\ܷn5ht.QJ����c��cӗ���`�W£s���٩KG{X�)QQ~N�S�u��ƹ��E�Rr\t"����m*/�^&�A(\�WSTʡ�4��L
˷ȹԄ$@1�+�I��-�T͝�m��֡�~8�5�@��� ,�|��W�"�|�w)���hO�a�4�l��L&{�3_i����8��tSh�Z����Vo)0�U|B"0T��dEܤ]T9&�=�?gH��4NCce5��������sYsaS�7#��_�M�8�Q�`�y��-��!�����n��w�T.�,J
X�������Yr���s�Pp����vM��ED��3�)�i�xV�IT��:�:@�v�O�Ũ���`�hh<#�>������2�|Dq��(0}db�a8.������Yy��R�mMHؘ-73O��m7i^�W� �>��ɀ�V%�G��ۇ�O�VZ&�jԅ0��\�¾�_�6���vΝp�&Ҍ����
L�p3VT&M5��d���D>Ʈ�Tr�&V�b��A��U*g�4D!r���5I�5BB�Y6dwDِ��*J��|_eek"tK��xҷ�N].�mK�_e
9�7:������<�Zͱ�A�c�@������h���X�	�dg�����]���k�}��@|��󎮢��'ORuf�V�w .�^ݗ�����	.
r�v+�~y�=Dn�c�Z3O��`I����S6b�v\Aƫ��ީ4Е(/]%�N*��M�<�f	W��B��F̔���vu�\�F�j���1^���Dt��=}�3 q�P�h��؅_p��
GPT#=�N�֛~�O|�]g O�<(b� �)���)�=$w����x�!��Ʒ5Z��{�}΍�˚��eǲ�HrQ��`��Q�?��GGQ���,ЗUiz,m�c��Ff�4���Gmbs�����P�RU�%,�������#��}RmXC���Y��r�*r9�Ј��������(��D�6��n����6��k�O�D����KՇs���3�"��,�:uS�>��3��P�w��*L�������j^y31@Q� �
���t(c�2d�`��s�A|��%T+v�����`*\���-|k:��_Tn�d���>NY}���*�4���F'x��	����oN\eX�&ox�z��%r�t���e��5Ժ����:W+"��9�BǓ�{����i}�)���!l0_� �g�c(�"���wN~,��X!8֮�hND��ط�XҴPy���Xc�X�������~����uv5�b�׏5Z����|ܮ0H&%I��GMPQ�~F>����p�wSB{Zĉ���4	5�V[1d��~�L*����D��l�K'X��t��e���[B��[�/}rh�n��s�
�"�(��gѿ��;�#Q����gsA�K������~�����چ'���_ fs���\�����#s���0J�(�����lu�y���J<�SK˨V&Y����(
�!�#���K�	~�����qVYC����?n��s�4K+=
�3��:�� �&T%l��o%��L�t"���ݡ����_�}$���T)����j`��3�O��(��(����U��s%��i��ajɛj��}�W2f"~����'���p��#6��ؑ��k=P$��;[p`���Q2�pǍ�d}���CB{��z
"��욪����)O`�;R����h�����K�]���'c�l��=��h�Bʞ�z(
G�o?:�`�T�5��:ț@�����Ά��ie����+�%��uc#�ZnS�n$6!�,�֚�g;b�=)���D�-�%�T#�^�Oo�@����\��'Ϧ4��Qt�����u����!y�VoY�s�zű,r��/��7��4/ac���h�7���� [���->��,�`��<�Y��D��e�?Ln�.9�0oĆP3��B�:o�&�%}>h��/�I:� fx���c�k*+Sխ��c��l���%��DxE��5lc�k���xB�P�b�W2{|�a�!�%/�r"U��~)EmA_�a���KJ
���k;����| "ˏ_4� �����3|!���MS)�s�0�u{��Kq��˻�?�US�V\��fZ,����Д�����8�I���x �3��E�� �,��p���.�ok�9����<���S�J�H�Yk	Ь���D��ؐWD�u�6}���H`�[�ѥ�=\��,���CP����g��"b+g��U�kP��hҁ�D<���Rq�{��Y7닶q���-~�Rv��8���)��h��V5��2��Ҹ������%�3$�|�^ƅ�(�.e[s����rI�T}ܞ��l� %�imݫ<�o_�o�*����
�Z�&K�.:m>���	fdV�'%V�<[�5p-ESO��X<Qm�v�.ɕՀ�K�����2�k�ǎZ]�N�C!�B�-��	�fRh3ȼT�|�^��x^���m�@'�����Q�A����à[��{,S��Fkq��z�����7sw@���E&���~͟���LL���=��zs����pB}�ʇM%�܀hw�K�[Yw�?��+��0Ga�z�ë��;�mt=��XbvF�'
S���\W���F��l{��3��$
����\��-�0< �G"��z4�S5Ȥ$��X,�]Mqf�W�ހw��6���Z�b|��d��x�[���%2s���p�&��k5N���&S���s�<[Hmq�.?1>�HM[z.�04p�/H#>Y?��-�dh�VGF�!���U(s)�/��a��߬ѯWA��u���Nq�iuƤ�3ں��� 
»!���n�۷�"�=`
�� *U�"�b���m��=�r��랧�h$�P���4%�p��'2z�rlW���<�k���_�l���Н��9����x�J�2>�$��ib[ޠ��\<���5ѷ	/�A�g�&t_�'ҩi�qt���d����8}�������1��V�@7s��8�����{X;�@�F��o�-�a��ҋ��ܰ�|5P�����a�r���\��N��݆�$ܭΦ5�coDw��J�.�=��l�J���5vk�� �k^��_�>LK�目�t�Y��2��eU���:�i��p�%��b-���|�ͣ|�Db0�}#Z'NM݅��M��q�gb=��)�L�	E��a�<�	/ßՏ�_y�X��|$��Rt=����Dw��������0r��ob�%�2�n��ҿL�{s���So�UE��'-w��	ku��z�t����:g��,=��ݳ��b�����u�x��p��3ki�M��(�$B8Ur�Z�?PF�N���Ĝ���NS�mJ������s���"R>�Β
0��H�8�}`]�	 ��/P"_I-��ے8{�;��;��QrY$6���l'�>�}�
��*^�w���5��a^�R�J"is�р�Ϩ�~��Y���ƣ�ᫎ�=����#3�+S<K�OY
e\k��ο�E���5�#�f�D���{	�Z]]9����l�s�[t���"����G���B:�K���HE���`omҦ=`R=��<M[�d�r�k���vD�G�`�T�[��t0�O�2�DH����ѝ?	".�B<��񠧃�[�_�����L(Îr�Gg�ֿ������1�UZ�5aP�x�-�/��N��0δ��Q��0��p�C��I�k1��5�t�X"�y)��W(�Z��?a������I+���ߧo;��U*���2�ۍ��LE�-o�鵒>������<<�Z槽�Hh��3O��
�͟~��K�����)���J�/sw=&\�j�T�M����O�h@���3����mӧ��Bq1{g�5N����ͮ��#�|�`�ef�.��ꙏƲA�G ��cd�^J�aO�|���Vg_9{~�L��Ԩ���pS>Y���VMR@b8��~T4sN���op!���#�:oB>��> ���7�!�T�0�x0Wsn:�_���Z ���#�k_0�c�I�t���@+���\nj��?���N2��~�9!C<Ԁٰ��|(#��4/�)�.ʃ0��wS�*;㼉pp�M��<�w��9K�s�81.W�g������|�-�&�W��Tv��v�3o0�}w����:�������`^f��!�!F��j��3K�hӫQ.�bӠC1##�Nr�rn���"��Wb���F'��JG۸���m�CE|>y]q�rP�?�] �� , �c"�7KGP�엷=';�%����KL��)�����y�D�p�����8��7.��J��Է'�����b-�ڞݣEuˈ�4+@ i:��-��9�V?�V?�1!01ܿH�"��ׯOIͼ����|Q�m���j��HH�<z�Ꮩv�H������ŞM֒�0����_v�o���8���lX���E��4�qY����f���gt���D�N�<zbMJC��)�^(�ԃ�)�g���S����7�;D_�_�hc{S��zR�z«p���]�q�|�=��R��?��>K�ݯu]f7˥,���X��	�pK�o���{�t�:0w��ݢ�!�$A�V�l��U�������h�
���OUhN���%��Qyrpp��b9;�]w/���H�+�XD���n�l�иz�.��ն��Q��$S�+��$�z�-x�!�������_�1�yG��]�gO�D��z���i߀���XbD�>�c��{A���P� �ŋ{�-"�/)�{��.����zF����0��.�?�ɯ�Ž����M�}8�J�J��Vk}�߲�k8��0�;��uW/�},�9�	��7XR��ȏ;���4�YVUkiyJ�����а�u}��
�8J�����[��a|B]��4�n��y��ٵ�JlAK}+x�P�k��=)���[�.pE"b���=�8��}k��̚�XjR�9�݀)�\@nu��d�J)h�Ԝե:4iƦC���`vČ�\Rzs�Y�b��>�<�5�Aк���P"+��
P����"o�-C�^�sTn��O���u(=(;����4���A���;Ӯ�D���\���(M��Vo��Ηxg�Sa.��p��c��yw\���Kwb/�����9.u"[��&Te������3:A	eŞ�x~?���D>���HI~Lqi�9!��\ǄQ>x�?>�D�ک��\;1;�K��j��*슰ކ����O��2V#���
e�� g��r:L=>c�ݓ�{�Kʳ�m�G�;u�ş���
�aZ���;�qI��-�]!UU�祡��]���S-�SG�r��W/h��kB�5�X����P\ �iݮ����O.s?w� �a/ݹ�;�1�\4�C��K��Z�U~��I��������Nz�iq�0#�-��rp����J	���9�'��$���ڔmJI�ы-��_
ݬ�kĘۢ�f�<0����"ğ���e���R:+���'��G��\�y�l pr �_��Ԯ�GUu�^Er�S/]\x}�Q�<�wp�9
�6,�^���b0� f�?E���|��q����"�#R�}B'�r�҇�F��	?��n�Iw"�_�	�~"ST*��z�_��R��3�,O��	]��6�J�N#AOڌ����j�o���5��R�kU��6��gZ
��'��p#��sʫG'���ծ��%��/����>Х�!�[���'yײa"�f^F	��
�+���s��
�8��a��F��H��Y��
���І�o�&�4���, �ݳ3BS(MKҙ���&�{Uac��D$C��6o��8�A����`���x�ϩ1�9�<,6Hȑ�!�S$ު{8&�F��,��T�W�R4ҳ�|&5��,�5�0B��k�~��Nj��/�� |�#M�����?��z��wy���h�?R���>��yhO''T���2�|��D���<�׭3�Ũ���3�X�n��n���+)�O��pOA �E��j�Ů�W�h�����"��X9eR�o^�c U�HU]g�Pn��D	*),����Ħ���ԗ�P���$ۗ>�p���tϧ����Gj���u�债UE ���n��Q���7KJ7m�8�9��Ve����!t��f�'�+Ԃ�J��x��D�C��,;̅r:8Q�9�������g����y\^�_eX���1ǹ�Ӵ�_U�E��cnщ��G��<[Y�~?Ъ!��1���7�\���2t���|�dtYKT�@#���#�֤6�� M�r|�o@7��1����j�������R�����q")���(k-s�c��������.[wZ@W:�$Ӛ�w��#��K���-f�9�s����?���_�	EN_�s���{�`��_'�Gb�-�˞���~�\��S�>��k��V����)]eA��.��G�	s3IW�O��؆���E?��+"�w�����U`�e҄<Y���3���EW���-��S�G/�W#/�*��K4C���0�fBϢK����7O���*}�!4eS`�])"�5���I ����r�uSsol�*1��ll��\�@�A�������=�\V3
 �?�(�ϕb7�r��gF$'x�Lފ��(q8z �N���8��\h��>IY�%n
�l���)�S��{2[�%�p�|\�@vִ����X��4C�)�$J��4Cl�<���&�l#B�����l�o`�5-�R��%w([� -�bR�P##k�H�����6�Bkb`��(����`���я�=E�J>Z��o@����7|֏~���uk�|g���7QE)eƛ^�	�>����9���� &��}��3��O���BO��B�����:���"rC�7vZq��U�:���On�F��j��$��DZ� _t+p�VR�e�l��2��:,�{�a��)F�?zk�~��xP�p�~p��]����!���� W�E���4�=��&���k�O|hlI�7�vTL`C��@hKHy����.��A����ԪQ+��^�/w����P^ȵ7[�F�iM+�0.�k��d���<�~��?�_���4���򣗥'Ŧ�����ԏ�r�������6�
�HeǑ+��o\�q,���o9�}�^Yd���'���C� a%��,9x��j6(�=�}�*j/��o��q)����)1o�`FICh���_��A>����{�wB�`?�h���C'����������CS��ȓH5X籼;ss��z�˳�e[�
L�<��~.�z��)�L)��[rP��:˄ sw ��<lߺ+�z����F���u0/�
�����&� ��if�t�s7>!����(���q�E���-l!Hg B�4'�����/eQjĹEo�^�r������8�-^���Z�{��zܙ��^6�Ԩw�t�6�$��G�oPeֲ��+�/����'5�,='��D�ύ+Z���"'�}�"��kϸB�3n�-Sb+�wݲ'���tMR{����~Hk��&��I�;�~ �*�-a���� #6���l��'6��ɣ���PUC)���vLr�IC�}dKT9�R�MK;ٰ��k�6�]�o؉�/a8��m����^{
����>�#kϘ�Gz���v��Az�v4�~�E&�	�wd�%�/�� �ZBLSƄ��"d(u�J����ݦ���?z=��@�k���s�C�4)��p3H�-�Zg�ܪ�#��ŭ�pM0z��nG,�f�j��$����J��m���ˋ4l�i���" ��TbT� n��3���:��Ue�`�Q���oő�H�\�ͽQ�Q.Aq�,m^�_�г3�~�7��0��a����n��񿓯��7)ސ���R�N�\q�(�`3}�g�:xa�H�@r�Duo!��nO���. ��r;Z��8���ݞӿ�y��Q��������:{�C~��x�M�&���������i���������㘌;u�ulb����9�5��z����*�Fx��RC���0vXf<�$SU�j�x��f����y������ho͒90�g�F
F��:�d���H�V$bC����}���ɦEV+8׫,ӡ��KS�k��u�:�|�|�Vj��������
�����H��'��u��|�ca��h�Î�с��ڢ�y�-v��=U�	C���b^>�Oߞ�%�G)�W�J+�Y�y�5�?���P��œd�� ���0�*fM�j�ZFf��m}�[]��ӿ�]�����Ը_��C��j��Y�4���l�����k��+�p1�D���E���h!��a�¦v��U��UB�0qf�O`�����ʻ��r^(48 
���)�(�UL�v�~p�ۨ���[�A���G�
?Z �������z�b
3O��'2e�c���>�y �V�F})�]�T\.���Z��wc{�Z�ݒÔ���p6�/;j�V����y�YiK7.��i->Nare#vE�8�����[k�zo1�o�G 4��
c�j:Usc���F��Ukb�m�O���������X\�p�\W}"(+O:��z���}�	�%����՘�3<,�b�z}��@t��r���B#�(xb\�6�w�׵;n:ʐ����(�K��%F-�{t.4-Њ1������������\#�����<�����nsZK��;��~g��2K`YS�1	��<�@L����4$1&���%!	��%��Rf�uZ`AtN9��Z"z����:�^�aM�����;�f��	��5�f{�Ь%�a�g3{�=/9v� 
���]���o�� !1�� B�&��P�VAXIS*�y�'�{�|L�,l��;3S�M�}��3�k�hJ��2��J����l�"ŕF�ds�;c�Yl|q��I�ߠ�Z,�k�������C4rI��S��*��10�C[I��W(>�?EG�X�
��
(PJ酿b������%��g�q����XР�m94�>��iBHC�����'�{ҡ�m���L�e�ζ&/	03�E��EC��2�ZeCYO���Dl�)U�M�����e�4�(���S��kᙷF��tX�8��3e-w9͠��KI1l]G6��!wŞ	(��M��䎻�t�� O��4�VILB�cB�����:S(�k�~eoh�T�x�}NI�4E+�p��_{<p�X@��U���"�ھ�Y2��t�_�D��`�p�os?�3	6Y	�������O�e�8�u (_���x)�;̬�[����4R���;��ƭ���EE�ET��{��,L�p�aig�`a>����d*N3���r�u��F�tPǞE���o����й �Z�i� �"8�� ���H��29q�&��>�C_�� |���A�c�>8`�a��2l�? ���	��Z<'n��X��?�����|�w��f&��_�#
z����u�l���;��Ӭ�ʪ��H�4�hfk����/����d�����LS7�f��|j��T��U�B�Y���}�^8?�Q��yZ���D�@�`��9�ʒ�h��i�DR�[��D�~��u\����L��	�#m.�Vz�%M�$C��}i�)�|��v��H��N�j���h����A��m�tN[1��O@a����/�+��)�eu4Ċ��]6�{��S��),���J�<��\��n���Hr��[]�u/�Ν3P�j� ��:^�����f��V2��J�LR�K}�1|���S+�0g�/���U�HT�� �&�����6b�s�چ+��&��+م��&,��U5��7��`���M� ��+1�-�ο���p	L�y�����:�.���	w�.��Gvnfi��0�o�I���K��u*ݳ�e�y�\G�-���柇��,�;�n)M�Ț��6�<
�K��;��b_k/9�=(�rBe����eK�-2��5���p���5�}u��1�>����ك��1p������S�{�كW����*R$�B���Z�Jm�����,���p�L��F�/�V@v��k������	<x� �,4.�!0-�ٵ�<����m��-���3}�|�rPCUz��5|�O�a�O���(r@�꒰��b,ˀ1.�'�̵h�č�\'%�N@k����y:�:��nH]����z���=z�"j)�@��
����Á��{��#(�#�*��*S�$a�l� Sb������B_x@Κ�p�~<��8����{�a��,��?����c�O���38�@�Nx
�`��|+��B$��Z^�fp���52-~�m0�,�gz6��{�N�&� O]��m1���y�@:��c<<�iI�q7�h�h�S��q���_KW����z@�Jv�Zt�̳A�^�>��D$�9E����o��Z�/tw�]9X��\��z{%�[���VT�J���yɄq���~���R�� ?8�[�M�Q�qA^v�7�䪩5�T瀴Fo=a�0O.�u.f�xtyvs8��M�ꑆ�F��=����T���LP�2�A���)��bh�%�0f��6�ᅚ	Wz���&������sI	9$�@DR�C�u�m�ˍG��~1+��:�&��tE���6G����K�'R��w�J�ϥ�S�7 (e���*��a��&nj�.�l����Z�$YK���X誟�/�`x~Fsu�+t��B��ӎ�f���C�ʵ��lrO��t�2�#ſ�p_[v)-�o8��&���jVAÃЗ���<;��@�R99z��
��yV���|R}���t3S�P{jP�|���v�zځ�����SZ��H.�8��f����W�Q,�/�mzY��<�i��2��xR���1,�j����m?2�+)����U�o���	��7�Ja�&�[�zQ���~�$�i"�̅���:�=F�F��jiS(ߴ(��&�5�u�M��-�qi2�a(�3�H�����\T�@�@��Bs%Z�Tچ���J�Q�M*>���\�{�fXo
�ӂ�e}�U���L�S^�����~����n&�:���HYf(��P��^#����/Z�~���p���xݘ]��*ʵm���Q,�����)D&X���&,�S���Z,8��C�C��gڜ��Ma'��E��ba�����o8�Ux\��4��Qf#�:�Fay �x=�XeZv�F�Λ�`Ej4�g�Ѝ�e�� �r[�S��|��I��#�HU8o$��7:)�b�#���/�hrO-F��u��V�J�'	E�� C�W��J��$��u�a��qɗ;'�79�$�.�����1�����#�xX��6��طЦ����Z��ޏ�6|�Nl�{�Dn���t�~G���x�Z���[�c
���y��OG���bV�r9|o[�m	�A&V37'4P�c�����4�Gx"�v���\��q��O��|�;�rMt�1нS�+�q��?�'���3�)�r��o׶�ݏ�t�:>�`-&�Q��?у����AJ��9���.�0[~�!ӮL�P$�/�rf�ї܈!���&CC�JSK)�R��>\R+��yGw`P���7�!Fr�ä)�.�Β��Fo��	�W����Mu {�_�5ӄ�� �F5fܫD��(�W���vvDk⧶�%�?�)0��]�S{�5#��+;>ǵ'�J�2�
��ѩp�0��dE.!�`ʳE�����7��r�O`Rt��㋏Y��M�m����Z`�¢��ߤ�iͦ�2�V�-�cF��>���BB;<"ޥ�Z���/C>օ���_�=~��ܗP����\���a�I%�v;�`U������*K�˥�䃴VP��Uw0�
;5�׵�
��+K>v�:����ʅ0$�
o�35�����J䱁K��۴�^�(خ�:�xF�sױH)�g{�-�ps���	�?�b �B&����<��02ߤ��1�C�����w��IB���wtoM�m?�+BڥI���:��a�t�aI�sK��GЈPć���H�ݰ��%\��F�bs�����boe�!���j���})A$n�v��X�����N<���w����#5J���ۗ�J3f��^�'�~r�7E��lr����˹ϰ��NL���:wYb<�n.w,�����yY�+��'K{�w�w*/�|�r�G��L�.�p�~%U	ۜy:��W�QM�KSkf�X���Wi�*I�̙���DJI���l��g��D���X�"m|��BoB�F۠�a�{�[��J�s�d���DqQڅ-�Nm�B���?
�'�
C�8`�>��N��m�a+�;A��&��Cs���f\N�og�B�(>ы6oM.�=}Ѐ����dV2^mqd�I*�Y�����4��!i�S�HQ���l��.H��U����s�۩��/͸@��tg�q�g��8^��=^Bc��}G;N�i�/����D�U档�t0t3'a{�E�E���U�Jwz�_�<.F�0 `��b��n�Q�"��M��O����{��$��y��I�;Y�1<"]������ӱ�;�KS��Go�����Ez��¤��v������4"�+�:cW���~}s.c!��}T�����i4i������d�Tڟ>\�ݢ�;�����#�g2~*\��N:��)E<~�T��A�+�m�|�߶R٘7]��fW�aՠ�4L��	�6j[5�L���l�E'��^��xP�跨��%�)��2�ϴ�����>�ⲫooY�I��%���:�8��p�  Dw����N7������!�8��eI�_��E��{��L{C�71(��I@��w�:�>[�B빻ʄ=(!d�n;�`a��)���W��ma�>��y6��Å�n�<���$3)��Vd�u��V���u�e^;I)��zy*)MI��E�xBP���-�}/�"C�
|�5$#�=�cr�Ke�k<`:4�"R�iE�GߕԬ5��)1O*{�Y�B@<sm"L�t������ �w�	r��;���;;��`ʾ�⪘�������OD�ی��^L۔qAv��L)���7Sb�vj�Ĝr]0��q/��fq|�DW�d3�����	8�d�U��=f�H���n�����A��uZɈ���Hۛ�;�Au���Q����!�j�2h�y�]�Zo �!��H9N*ơ���h�\[��B���{Diw؀�5)��_�D�:�&�\6���ƶ>#�7��ѯu1x���8$�m2=���}#��eX��ڵJ��,�Ĺ�g/���P�Μ=��c7c��ԁ��ce=EK�@���U�;�P<��[T7����\r7)We�E>P�>�����q]]�∶&�n�������>�fx�Oȝs�ep()��9�u13u���C�hw�������7S�V<+�*[M�m��2��*�ʸ>����:��Y�����1g}y� V��h�͌�hp rp0�!���ь?�;��}�op�111#����pEA��e�kb.=o�'@���r����=J�'�f�a���Bm=?���ƥw���.���k��X���0"ʂ�=2>u�ZA�>�qn��(H�Y�-gUu^�N��������;Y��V�*k�gd~��OCij�t'@����A	���1c�q�"\Ve�ѩ5�*�p1A!��\���^��J0���9C(�c�*�KW<��n#���ʔ	Y��x j�7o(J`hYLC,Q��ѥ���I~yר*
O��q#������j���><��m7�*��������j�ce�����{��Ie.�1�9��`+׽�*�:����Y0Q���F�R3k�!|�)�~�.}(�.��f���d��/�Y2�!j�}z�mY����-CMQ<���亓k�q�4���$ʁx.rܶ�6f:߾�ƥ��h��8�`>+��^�_1,W����Lw��HIགd-�b��u�L���~~��E�G�ǰN\���ϗ�;��G��k:�>Y�m�?���+7q�B��~��k�̳bd lv���o��y�k���'	�\�Y|ɑ��rv���;b�E"DqK��~�i;j�\#2M�U�_�B�����?�0IĪ�(�;�6A�c�Ʌ�]���y���e�nl`��dԾ������ �fߊt=�,et��~S֥y�j&�I��^��!��#��b��}(|���'aա1�\�[�}f�+)��6D0��#�i�A!y�̰���� �,p����գ��YZ�& :��7��;"d�Ws)i�vFS&��S��Z�/[�y,g��`?���?	~��~F.���f�"�eVH`h���}�!{��&�|=TCF�Jŝ�� 9�����+a2�$�r��ZT;c�� �f�l�u�=qZ�X��ۋf�R"ror��%��h�LO�b�l�k���)~`�E�|�0��ֹ�e� ��Ѫ�G:�c��s(&L�~��uj���/��$N^cdA���(�ĝ��.4����%5����iY[�qEFP���sW�W����߈���}�\r�}ǟ���|�ť�hO#�`�p��~߰�l�3�~�V}�B��h<���!��^�|˭��v��
������%���3` |�g�@:M�#9%����T��4���!� ׸�
�L�R;��׷R�*(�#S�ɂ}\�x߃�]9�zޖ�Ӧ�A��)��ջ�l��׮	R�$S		?L/kJ�'�z�$귵���k^!��ZFj{F[n���y\��ӖT,��r�H-�W�u ��9�Q�hHFȫ1x���z�3������!Y�-1��0����]ϊ�=�G���b��~ʩ�t��g;�h��+��M.��y���"Y� ����u��Y�-Dc����(��+�֛}��erV�y_P�c,=�p��(t\��kQ/C{jc���&�|M�R�G��gw�VW���.�wI#'�B�0�G�4�����n��4S/�
�T��!�^�YބRS ���S�W �$��s��Ē�A�n/�1�$*ޡ��d���|�����Z[��pD�Htp�J��Cr`~��J���maLX>DķB�=!Y
�B�bF���h�̓�V�[ͮ<��	<�X��̜���� �x'�4���ӣ��3�+|�
Sg�Z�bD4c�%@�$t����{��=[���`�KP��ֺ�0B�n_ o��h6"��Kց�����Ͳ5أ�߷��OK��#���o�|#-bk�zf&��N���W�cJi<��P2��
���&�)Y���36$=<�V}#�T��%�(��X�f�Rc"�R�VP݂\H�P`w������G���A��7^$0֡���Dx�n�,�(�_��E�:3y��{��]f%�J�~D�'�V��ml	$�P�����oU�E�R|��c)��:B�3�HqS�#��r��V���&pn�!���A8.A�_gs��T�.	9�\/�pPE�����C'N�������#5�,����;1��+�7�v�D���x��wc�UO5w_}5��!^P�M����-�f���4�_f1��q��yi�N��5�Zpb]�d�y��ܚ
Q���PЫieY���8^츳C}��uE��U�pq^_V�Ž��[^����jR��6�	j�����.�L��0�)��d�
�A ��y4���K�c,���\�؋��
�G�b�5{�_휞x<�VR��N�/B�9a�n
=��o+?�y���zt��E��dbXuB�VRƧ�V�ȕ���Uf��w�_���� �W,��z�9f�������)NE���~�SIӓ��q�Y���i<�4I�K|����^�����~��c'�d��p��#���1���R�(U~C~`���	� � WR�+���$e2J��y%�3���vY�m�ʶ<Io.�=�7���ZW��~��m�A8��)y��ql�{�&G�w����I���X]�g0;��hP��;7F
��k�+�W:���2��<�D�*�&]Wl�r9׉^�`��Gs�T��'�W��ځ�:�fwP4��.gμ��N5�6�s��ho4��w?g��?���1>ir����䃃��`��B��(�- �1��I��2A#�*i�gr�c1,��1W}���L��=k��Ȯ�{�����%�qTd(>\��[�s���2Y���yh�y�j��v�W�sv��jy���_��/E���0ޒ�O2�<�t��0=hC��$�3;-V��Ê������F��/{��g(��*��k%� [�v1�~���G���f����YB���E�õ����_�A3�ܧ]�H�H�UWGC����z����/�nQ��������$�Nk�kq��J�&@ �p��K�p��@�A�~F�n(����D7�~�30�d�b~���6C�uh_-�a�������"n6c6���);���N!}X������(.��RQ$T�����VIy��6#ɐ/�H�Ɋ	>�������䬁՜d�Z��^�JL']� oM)��Y:�mk>[�4,�������H�C����HIN\S���{��i�G�c[Ϙ{�ȇmm���O;�kK��JW�3���<lf�O@p��T0.�� $:��?�͝���,8��(g�
�`��{�ac�<1.���\h?[Zf�V�yhTWb0U��}=�yJ56T4w�"�J�s���S,jUP0�1d�%E����aW��ԯ<ҝ�>�Yo�牝uă��%x�K;�7�t�4DQ<����{��J{�7��F`T�>;�nO�zO��(!�6!�/�B}Okv��
^
���\M��`�}TB�W������pSȸ�ڢ��Fӥ�����?�����@�j�F`^u�9{g��v�hM��5ӓuN� �ڸ�"rev�G^ƾs��©
���c��bU�J��JD[�1�1�g�J�mխp�@xT�\B�W�Q��e�6[�zt��ͪ���@�X^?c֪]�&�����4}:*�M+cϦ�sz&F��Q���0��\F�"y�?f�.`�&�-W���t��02��T�V�9>�5���E���q�	0 lU�:��Ýf��
m���`M<�P���@E�L�����x��hį��j[69�]�m	���;1�x�H�
y���K�f�W4vtU�
���pb.�����I1΍2N1�3����5�w�D%tW=KE�G�a��{�<̈U왻K�N$�fW�},r��;N��rW��k|G�;d��}���$1ߔ��4��*uv��[����^��(���0����w$�r���O�r�-_���m�9J�S$���sXBJ�:rS\�H4�|q��Ձ0i��ή��#.@�;�X�6�8�L���<Q�5�6ya�҄.d2�4�
m���|���w�M �ŋ�l�5H�vI7s���A�]�[���{A'b���gn��W288˿�|�QE���EMi�����t1���FD��
t�T�����ߐ�(i���?��\�R����7���}��.�f�<�F?4��)��c��ʡ}���o_g��!�zu �)Q�JD?����g���1�7�J,�U{Qz��O�m�L^bNWR�5�-w���~Y�Ķ(�p�v3޶�����h)���iQ]�r�.������7<�;�z9D��3j���G?!|d0F]�_��_�v=�d��k^%c/���O��&��p�b�[���oH���@n[q��D�gX�*q�4?\"�F���T�w���g���1!�0y�T0I8/A9`(��mU�%�[c����g�u ++\� ��$��owY�F��I���4l�C-�q�
>�Nz7�EЅü�R�E ��P�4�`�L��,�����O�B&3"c-�Tֵj>;����p::(DHTy���a-��24����.�A��w���h�u�K�N+��YY�}�Rz���C(�`_p�Њ|Xe�e|�K�[R�!9$�U��q�_u�7Q;L?��M�N�W�͍��
ʛ a� E\�-^��/���@˱����#m(������RT�~	��S�pk����"�[S�:H�G]�}�q�̲� ��2`ϴ�F1xj��;�2�,sV`�X�/4-�}�vy�b_�:.�1�O�$�n����0�|ں@6�۠K>"����3,�vԙK�8�d.�Ϻ���tF����8M/NTڸں�z;4�@�m��jDǞ�F�z�s���%ed:U���0lJ�� Z��i�_�Z��6�t��,Vp�e�6��H�b"*��t����pU,�(,�Q�F^*����ڒ%G��((���3�e
yĬE�����t�'9H�L��2L� ������=B���q�FV*��_��W�˔�ȭX���\����^�ƘC��i�\[�^��N^ԀX� �]D�^���\e�� ���=�b)�����Z�"C������'���'�n����1�;N$�B<<.���]vi����H0܏E���ЃX#�#�_d�c��nPi5y%�~OD���=,�kӄ�)���<�ʒ(�C�����N4�jK�U�mW��O���[���X����`�"� ���n���j����R T����x����Y�-TSG9���f�g��Р�ԉ��s/Ѷ��%b���΁��r�2*I��jwm�R��^�F%�k��0�}��f/~r�"�;���czs����?%�Nz�����:\0N�R���JnP	d��[�F�ׇw��&'m�$n>��N��=D|GG�f�R8.���	��ew�lD�A��Y-�0�/H\g��b���I��7l����I惐��4�L��)�9�Tp�EϜ��]��;��8�6���Q�}��fh�v��0�=5[�}mM��9��{c9m�?��%�#s��t&�w�.���0P�X��Ua��nA�vL�3O<�܍(���m��ށ츸;)O�#<,DM����iL���ϯ���0Q"����|ƃ�P�V5e����������;���{�99a�M��66�d�e,�1ļ} ��d;���Ҷ�y�|Y
��Y�k������]�7T��g1c��)p��uۗ^U0�fR����<5���7��r��	m�1��H
兢���_Қ-c�I�G|e.?�O@9�U����#��HU
������4e��ܼh�O��P��V!��d��0�ĪvH�+���Go����8�~����,���jj"��d�nq�֨�7ӓo�^����B���J�L��X�c��Vp奱���&_��m ���U��9W��>��I;����j�`�G+7�Ŏ����+�P6X�=�@[��cs�)a{�KF����Z	����h��&�qO�3�#�+ﵻ�}��p�%��.i�7� |�LI��r��X
?#f�y��� �c�t����*���+
�M}$�Ft5��D��v*���� yq�TY5�n([�[�6h�_)L���w�>�ͤ�q���D}�i�EL	�^\�����s��|\�H�������/��'쁂�@�mDH�Z���\������i��s�`���Z�wN���D�d�mIa9�m��g�r��KD���<n����ז��#AV���'��avc�}�Z��g�ڦ����e�X�4��wv�|�N].������i���3{"]�w�&��˴%��z>EW�a36ARB�d���l�������+,QI
\����iP���B�s�G*1)�����Q���������'��{N�~�Z'�:�(��[�����YI�4
�jQ����Z ��prj5;SJ����l��D=&1�N�<ɽ��#jCǸ/�r���r��-���![o:�:(��>Q�^v�^�rR �W.��G���.,�~�G���ib�;�f���(\�^��͚В��Ӡ3 L��_�Urr�Z����hF^E%uhT�Ϡ)������d香�����oX����+93���u�m��Śa�.0�L��W.���0#�B,�	'R�D�C� ���'�kO뮇(�=��E[>��{���sl\l�v��d�E�IV��� �_r�tu���E���ߐFG��}x�1FђB/�+�֡���<�/�(*S"rn9ㄩ�Ant��.�(�,G��2��;��E��hB8p���-0Y��)��Wj�.�n�����[(k�1�z�O�4=�n�f��l	�ɇnZ�;F<u'D������u�2Q����1�b�JL��BXǋ�(��� �#��zt8���"�ª<z�[C�*�n ��5������f�T�N��˙��-��������ROa��@��86*��<�م�צ6�e3��('���.�N�?�n���R����a���`�B�G6���VH,൏�V����M?s�T��4�X����*�gy�ݫ��� '���<a��5|#n�$R?W��ʃ�ִO��A9j�nG�V��3�+�2oW/)|�$ 2!h�y�K���]��5��*���^#�2/v���T��s'��{�=���c	��8�H y��AH/9��bڟ�O����5��CקU��5vD�m��ȳ)p��N�q&2ע�K��2|+�R �2%bѰ�{8��Ǒ^$��M>{{zc�d��L�*���W|N�[c�?��+z�	��SR,+5-r�u�������N��/1�R�~{�̕#j�$.Õ�7��q�ҕ9#�.�f�I�m~|�����q�� ٸ��$�lXyX�V#�3nA��s!����I�	��DD�� A"������8b�ɰ���{K�7��PuBp�;���*]J�~IWwR�=�-��"9�1	�7u`�X[TO=I�����
����)�D�Gj>8�T`ͦ�[�#�}�lu,%��!�ޜ%l'1�k;<?�,w*�x-�=�?٢�F�n݊	zO�ɑժmVPF�ۮ�u�j:	�I����
]l!�p��;(��B$�����ѴFjHAv=�87��V�m=��S ��n~�Ǚ �sY�����}�k@�6�)xeU�
 Yx��G�*�e��FcHU��_eFEUό�-}��{���f�ܽ��?PZ_Iy^�3��D�)I{e�E�s���n�k㼏�x4J#L���`T��^K�k�ֻ򃒱����G���[�6����8�O�~��s����I��`6��L�\��S �xҶ��FC��,��4�# ��5.	�Z�)��6�7������+����GI�������6`#M�I~f�r7�'�G�ϐ�eݞ�E�����-4��F��ڍle��=>��#�q�lME����ִ�>fZ�!�8M��)g�a�J�͛U����Ɏ��ZY>~���˰��i4�po���"gj���8������	����ל��k�䦃�5��L����l3Զa�ng{���M��w�����ui��:n(�y�L�Ł"�:���,����XS���\NV9�jn#`93��&�C��.��owI����t�5�j��=��3=���A����O��4��Nx�g����Z綣��C��v-:��)�  �b���b�RO:%+r��BF�VjB��Yǯ�扊�1�(
%z"K�c�����nZB�nT����p��q��(B��P9�Q�O-�'�����=>�C�:�'��ji�c�|'�9�#���\S!h�z��f���<D��|��Q�@XjNI=�O��kB?���>HG奱T�� �Pk���(��ئտb�Y���u�(��LGa�m��	H�ǫK������ۛ&t۳��s}|Xo��Za;m3m�2 �=��M�-���4��J@^X:���w_�2�-���u��&f;,��Y��͗�0���w�2`'ɐ��1{\LU�\?ܽ���z�O>���B�	�6rNN�*t5��H��m&N���Rt�<8��K�b)�#�cZ����o����d���S Ȟ�c��X��Jj�I;���<�7;
ň���0̬43g��vˢ_�����t����Mc�7jW�J�s56;iun#�%@�;�i���lk3$ꎃ����V��(x�����������u�ppd:D��0Ȯ��-����qJ�l���f�?*���;t���I��U�e�^��[�K��<�1����[ o��R���(fø����-TL�8���	����|W/U4���	�OC��t�]��@�H!��n�ߟ�����Yx�=��S�7,>�,3e����2{��|���4~��}Q!.,>ԲA+�g��v�b�e9D:������t����J�"j�e��c���89�3��(���6��p��}��t�^��"�ЃR=�[E���0A&w�n�3S����� �v�#c�����R'nX��@�����\[`Xf5z�%�Y���H[B�U�@���p ����-,�G�I)�!Q��$
�pGn2�*N?���Dl�;�z�M��Xt
�C��]"QO�4$�	� m ݈R���va=O���hrU*����{O+\+�P�5WԐF���4ӯ^,���*�_�3jB�/Ẩ�ĉ�l���q�F�R:��S؟��v3ٟE�R�<��_�Ց+��3LC9J��>��1��/� )q���xB�r<� ҩ�~����od�r��,N`MK"�sh�<֔�W
�� 3��W�)}n�\&aY���A������M���{�����|h�� ��g�߽�x���Z�V��*�=���R}���oVR���Q�c���4�a.ڢ��"��'oѝ:y�r"F���r����j�KT9�)�M(ש"'�=��h{�r
k���-7 0:�v�6��r
p���X#m���S} j��ȸ�w�:�wΑ�o/�2}���_�3���h�gD������Ͽ}<�E9�t��mj2��{,�u����.Rco�')s���]�U,����+��',�ڞ<#�(\�k���;UK!�
Pw��AM>Xθ�,�x�[�T��CmuHn֓�l��ֺ�@{��O���@��;�Sԥ��|M�'��?�;�Xc��ڤ��0a�w��"m����0�`(s`ҽ,�Mܙ�x�����M�G��W�]u�yl�V�3J�RpFO��*��=3Ԕ.&^�C;��k��k
 U�$�#�P"j���0����B0����G��T���јXX6�_�H�{�����y4Y���?���]�;X]a-7P�Q�>�Q��9��Ya��XJF��_�^�O�ơ�:8S�;�-����`&�/�\b��L���l�0x��� �1dg.�@J3ݬ�q��z��Q��"�N+/v�W��2V�(Zck��1Q��~���Q�fM*\�Xd��!��ϯ=�IwD��pY/���E٪5�LP�O�N���2����hH�:!u�f���H����e���o�>Tt0��"����;��������
~nZ�i�[e�#�^j;H���A���m&-�W�q�^�]\_AN)�B�8��C�g�i�7i�!f_N�?R���z����8��븧)�\iĨ�G�ǽ�"��;����
x����s2%���7+v��=f�m:j���#���Vn�V^t~�+��M�Z�%�3��l� 6Q��#�����E׵������^+^g� -�U������Trb��� �j��ל.U�\��Ӣ�cQ�(�^�i4��ٓ��u^�U0N:�IxcJT4A+���e�P���gcY��ͻ~O�؆H�����w�cS#.B��MP��$؃�q|@�� �AM���2�
g��ӇZ,��N0oA�>�j�ݥ������ϸW�z����}jW��w�8�D����;�o���S�����X�S��Ϳy.��զ�_y�Ϧ�]�nP[�IfJ�1T�N�����������
׷�\�\���i�A�]�#K��g�f�L���l�lOL]�o\,)�8�
�]�#�l��rnk�J{8;��EM�J�*��7���R��mJ6su�M����B`�9@_s���l�.�ɏ�ܕ���k�̌���U���t�b�'��`��=�Y1���n!�M���闰�,��K	7�L��qRx�pLP*�s���B@����3�A�94{��g���M�G���$D�s�Z�?���ʀ���\҄�؎M���AH������e�����X��q K����� �W��o��aG��hh�9LffΔ�o:@� y(q�����D�K���D9�|O6:9�����l`P�L�׃J���l���������!���W T��=����ɽ�yֿ.G�!���ʎe[i����Nq�Hy�?Wڇ��d���n�C;?�[��ې� � o��s����Q3���k
��_�,:[-ऒZ��wK��}K�}GY��C4y�~���'2ߛ��;��2�`F����>��/�WoGHm�ŎuZ��� ��6TFFE���ݳ��]���쥹�\i,=�n�~Grr��mK��l�k�Mh��4��uat;��HC���$�}Ym�`�9>W�2��*[�����Iue�&��� �.#���3a����z4��x���D���S9MP��m���DsM����0�0�V:r�d���V�YY�Z�j���HNx�`&'rx5w 0����2�j��(<�0�	�Sw�f�5��k2�fM��O0��ƒ٫5ȩ'�8ҟ_A="�ltCi Ve�?���M���@4A�0�s#cI#�!j6ړ�:}r�D�Ȫ�Va�K�W����ʊ��n��U0&Zt݌����P���R0�+�$ef�u�p?������k��`�w�n���&�[ͱW�Tj���q1P�yy��d���Dި��mĜ����~�?� �U;�H�P�pM[ dy�&���$��h���]�'�+~�MhT��7��R\���'��$b}�w(���DŔb?mȂ�5����|����r��@�3*��zt��(�F33���a�'�<K�ʷ�U�_�X,��!(�8�|��X�>:�o) �t�����W���t1ʩs���ˋ9�c>�mz)ݪ�d�*���
�=yy~����يH�,�o�I����tt%����L�g���Q�1����̠�Cj��S�S��W�^A�>�u��T)�h�j�"�;V��*�Ij�*��� i�1ǷC�(��{�U��6:,�G}��Edi�Qq�n�\�qer�Y�\���5 $?�{�ػ	���y�f?���^I��J^N�{�JФ@:�s�n�b�f$+�>�����\w��J�������(.qf7\�J/z��[ݶ�i��+G����Ŗ��������gˋo����Em\��X��Jhu��s��K[!��N)��A�`��,���u�q��C/^��]	�&��c��-�� w�u�Fη���ؗ�'�����a#����z����(���*�a�	�#�O*�~
�ǅ�l�I�dҨ�4�<#�v�w��Gk�1R"�>|��^%KDt�c#�o���&���?N�+Cs��ǀ�e�e�.��-�b�b�y�c��C� 70i+,$��64��8����x�Ɏ�<+����-V0c �J�Yx�@�3޾�!�&I�p�N�3)xL�`d��m��	���Ә�yK�Z�n�MM'|�����=y�C��ErYg���m�9�k1w���B�yny#�i�ha��}Ϟ.��v]53�v5��ǟ�Q����Đb�5=���8�D�-L���Yx�jģ��q�(��^\�)*�� C�>����uF�_�)�*ܙ���*8meF�L�M�>��2�R)OK6��V�ⱇ|��	��`;o7�N�g!h�?�2��o�M(C�:gL����N)tV�'ù]:*��#�r�]�0ߕ�^��Az���9�1� �Z�D,̬�|J��x^86�6�W �Y13��>��5�hahj(*��!n�ݚox�]Db��#�gN%�o��9.r �ᵉ1�	B�\�ݿx�
�����K����vX@���F�x7�J�O��.
36��r�6B�F4w�^���Nj��@m���X:a�>�^N��F��({�	D����7����2G=H��6/1��cq��:��:B������V��K�='�\��]D�G��q�o[W�cZ$�hZ5Q�� �Ԃ%��w>%��sߚ�DQ�6/�F�E��iVPn�	�ʝX��_�d�/�q��l����eI��'q=[�?X�A�Q����]�����S[;@I!� ����r�
��$�9~�fׅ�,�rJy�T����1j$=�Q#9���i��_TO�9D����!WA�/�A�����2�b�c,���e���KrR-�8C��@mI�e��M�^&v�b�������w_$nZ� ���~�C��������dsp���R�.袱jt�X�F6Q�_#*�+mi��0���I�_I;,c�U�I���<Fj~Egm9G��t�\aPiP:�(�7�C%[��<����|VD���/W^��n�j��Ű��L�����\��o��Th�M�7@�ɿN*Ç�h��x���ЬYx�b�@�y��&z��f���b��׸Qdv`�'�N�B}���d43(���\X��ʬz:�:�1�-��Ea'Ĝ�}��3*[c�'�ޕe�0(�k{��ݥ?�����>-�xޞ�[3Rl�yG=>A� ��n���tA��'��U��A0"Z���s�:?�~	R<壮4(~�{��1�8&r
�V8Ә�!�b8�$��}%X�������|�I᭦�S�7T�^�!܏(���۬d��kM��T������e��̘��o]N\���hƄ7 G`����g#���@�g�Z��*�Rz_��V�0cEx�IJ�v:�WOMbX�g=�#�r
�C�"o��v>�}H�`a�\�o�[ϐÖ��pj���7o�M�JF�-V�p��|�r���a�;�JN&p3�zŏ1��<��]��;3��:�-4�b1u�J(?)��z*L{�I�M�G�;�0-�������x�ʞ��붙IF6�|�q�7���"����EC����$����mE�C�1��f��f'Xo���+� ��}2��m�7���.�LY�f�ԗ"�P Q�RYz{۬��C#�VUi� ��[�T�_nMw[��.�BVL������ ���J��;T��5�G$Y�~�[y\'6��>(��y�K��`b��+�����41�8|���d�=s5Fe�D�9I��k���O�f7����B�vQ��ٜu^��f���'j}���
����:0hnW��S_O{�ȶ?>8����m �,�*�j��Ŷz�~�:jJ�&lW*�o%���c9��y���[$�kVN���G�(�0>3��5N�k-!>�~E��/��\Kbk̕B�A�V�����1̴�T������M/�m�L4��d�ZG��8џNDy�Y?���D�I����%��S1.~��uI_wRl���=�������M�	FuI֜O���ueG*����4=�L�フ�ðJͩ�8�@�o@wj�rXNǂ5�R��6 sE� ��s��^;����_�L��;��=���e��v�}�6gN^�cF�~O4��������(:��V�]�c�A��^ �I��������-1�]"=��'[gȝ���	�̷Z��^C>��lAشE�I
R`��:��|�V��w���sXú���A�ɕd���:�S�!3�gݳ'��W�)5���O=���VI�C�*m�<G��-�����ZU��7 �&��v�h����6��٤��޳A%%�e>9�G$�|��꽄��-�R��l���U�z��BR;`ߩ�����Q<�r�1&TZ��Cl8���	��X2!��T s��+$�O�/��Y������V%ڟYd;{)�6���jEFy/�Cy�e ��~�^3����9TUg��(��?�cJ���:��V���5�����vb�F�nҭ�����k�����X�~=\t�#��Mф�sC���J��[E#Z`��?�eq�
Zg]t�����	�������P0���N�nl�"]q#��(�ƆZH ��H�Y��R�c��s�������	LQm�S�9n�g��&�*Ԃ��a\���j7�هW�U��֦���݃α����`���[��nDg�_�PT���.�2 �A�8M��.�x�czK��k�)���A��a�*�u~l�����YR�!f�I)�{#'���BOϙ��ReUr�4:����ն�|�sګ�g(h�(zR�^�6��������t�%|��(;��a��v/��UJ��)�݂�,P9S-<l"�B�b)�e(i���#e���B?}ΐL�%vѰ��E¢����l�l%ɼ��% s]�c��.��y]���'MY4�U��,���e��q��V��i��!۔Kmg1�,���gD��-F�6���4H��C)�a�i��^
���/e�w��I��_�g�}��v����-�Y�t����������Ϋ��m8�|&j�`C�i��c۵9	��8C�m���s��U��`~�٬�P^�~ID��;�R��J~�=�uys�R��� �M��϶�aŨ�Ｘ����E��������F����_��8O,����W�@�4r��åi	Fu\�/���( ��=���.����0��F��Q����F,����C�ȩ��H�CknЅ��&Λ��Y1D��pp>�ς�?��N<���*��1@�$�)��5;��Y6�˯'����F��Yf�r�G�!����Lha]�͂G�ó*7C�X}����p"�ٿ��+��m�4\a�������g�A����6�kk�|���4��X��α�e�F��j�ڰR�`�Z�K�Z��#�v>�\,�3�P��l�S����!ě��?�r����B$�N��s\\2�8T���#�@?�0���^ß�s��gأR��|do�潠!�R*rF.��%�1Rqԍmr���R��2���`&s-CV�ꗍ�K��{l���[��DU*����C=� �m
�]�[
���\�k]�$�8����,�#)3}�5�Nفa��
�u�I���׭�n����.qdU9��s�ϔ�کm{W��@�~����I7Ʌ+��"ȵ0�[��#�>��Ό̩	�X� 	76�9�7�������e��ݾ'	>�dg�ɸd%�:�w�뤟�ODۭ���(�B⇸�������ǥ)�~k	I�%w�o��u��~3�ޗ��Z*a��� DZҲ3�$����ߔ�P�Fia����i�~A�6�������*a��IUd~�sQ.�M}���CЁ��5.�*j\A�Ûg(V�<9�?����h�hV�t(e1
P���8��ܰ�xB�ý�X{�C����Bj��|����ݬ��R�	3��� �t���\#���a��/ރ���QQx㞔8��x�Y5M��m��.�0g��( hZym꒼Giۚ{Ri�	�$�o>'���+��������֭�u�sW��j�Q2ޤ=B2EfLtO�O�^�u"e�/�N���`��.�P��]|����X��5`�)������T�ts�]�I��:���o�į�^5��6�L����`2����z�D������|�y,�;2Q��-����w�؄��'�V����5=��Р����_�@�h.ɾ�v+��<HNJ�R����U�5܃��G��`V��P��9�-D^+���L�Ǘ���RAk[�L]z+��`O����
u@��A���=��.b�"
)��W��M��F)���xPą��p�x ���<���A�b;��9tJ��#���3��|N��>�,hy�^��A��0���򰟅�i����8p�0RO`�ZW�mh�y9�� ��ܷ�����;1�"$�H
s3��q��颱�2˽�2Ky��^ �)+}iĥ:�j���q�H�b�Y��˚ᅔ�xǧ�N��~�7֢`u+���2	���ʭ��aWp$�P�������D�M)�=d��(�6��Ln�_�ܼ,L�Z	�f	U��|���QF@�@&v�O���8�A'�߬�� �X2x��1_ ok�x��|�o�w3�f�RF�(]7v��/��H���DG�M4�[,�#�Ҟ���i��(@�VM {)b��W�Lף��_+��w�t(���H�� �ѽ ���]����IfMPsh�B V]T�.�ɉ9O��)M�׋�ǚ�g��ɡ�Q�&"?�oН��`vyUo{p���zE���� �o�������J[:�ⳡ�HTvԢ=hQd$�p�����c���*�e��>���E1 �m�X�hm�ۮJ~'жJ�7�B^��0�N,8�0M������o�ɐ9B����
39Ϊ���"�m�z���4LE7�=��C}B� �2�i������y� 6���>@�i-�!Xc��Ӡ}&c{������2oƾ>e�'c��\A��o�X���1%S��"�$�I5�9J�O��n�^�����X�=d��3�O�*�po�ST�"e����U�t,F<w�2�̒j�
L�|��q1R�P�U(���B�if���#���4�:��n����ur�'^��(�2�O�?e�D��=0��-F��~� ~<W�ʵ���/E}p��k�]�5�ؽǏV��k@
O�>t�N�mzk�h+��Jx�ݛ>3aJ Hˍ���IzD�+
��Ƚ��4�q{#;N	@���/4���l�{���"�Z��#X��"u�o�I��N&eA�<�꩒��[ͳ ��Xگv�������ѧ�0	�~襝K��N0��
�w+d<Ό�Q�z^8X(zHl��Er�T,R��v�xd�?��`Ad ��IҸ��yt���0�)6����/��L�(��6K��:�H���v*�:#ze�
' V+�� �
]��<�=����=US�4MB�\+����`�r��>r�]Vr��D�Ag����WF�@o��j�a��.bQ�x�X ~{tɬV�"�$�GF�Or�j�h)4_nQ������U�Oڝ�Z�(>N:�_�+�H��9 �Ƴo8�3�X��.�=����~�+�	��Y���5"N%hl+�����%��� 앧� 8[�@�4+gaR,�Ƕ;12]&�B��%#�[/C��^Z&�З���'n)0`&bi�##��4����ׇXȸ�h�$sCA��!Br�ɭ�-��rnDC�CCt0�^� �%fhwhF��=qэ��J��LۏxAya�b̺�Wa�5�?9-��]k`b�B:H\`�G��yY�ް ��B�&�.�}�<���h ��h!�I=�諊ɚ	k�{J=DM{�!T%�l�;��3|�C~�Q\�N�ʒ�i���]������v+�tb��~�EFQ�`Ϳ����*�_��B��xt�ٚ��/��S�������ߔ��.?�I^]��;�~���A����fq�j:ۣC���p�*����@y�!�Y����2�;�P��|eX/c�C]��:;���k���h|�<5��$�!���z�Bb��5���i��iD�J��Ӯ�.v?�����8Xd֢˴7m��(ϻ�Ìb	�k���rҋZCK=;�me��!&g)R�Q�	g�S共\�f�	�K�gBo	Jm+�<�#��c��7�}O��+�
����r�KD���� �T��{�z2�aLx�^X�bGa%E$���ҝ������K�ַ=����v+Z>��2��+l�o����4%]Ő�Uj�G��>-|_�ǝ��P�� �%w��(�7�z%B��������;����W��S.}�'��x�LRϳu��9�e�� א����}`�O��J��?�*�X����Q���S5�l�B��9r�EFE�=y��:���P��+�z(V.c
[f:@Ap���}p/��k�)�!la2����iuU 6����4��l\���Q����*5c����g���!a����@	<�'�i�����No����O��en����x�zG%����u�KX��}���O>q֛T���ñ&�ڔ%!�]uݹK2���i���O�\j8*Mv"��U�}|%��^�+�2�*�t�z�Ǐo7x!�H{I�
D�L��� 8�����>�.0�3����R�d\y�.=��x���sh���|���u/�p�[c4$.���u��n��Lu����Ba%�)�/��	!}[M����c�(@�y#�u��Z�57Sv��?�ӓY�='�X[�m���Mq�a��������*�\B�K�|�d}R�o-�y�<󤏶�&���&��� k�ˋN���,� �����X� uE�Z:uE��6B��q�Fr��!%�O��w�};�"��~j/}+&���d#]p ��A��[�<"2�m�E|/��0"H6Y�I�q&F����L�I�y���	��$?1ʊ`X�G\㏚,��wm>�?���g;�-�֎�+�y8�I��{�Af*�Jb�vr}�Ħ6���K��L*���

�1Y7H	%�n�|��*}g7�U3q�ݥ��H�?������(#��.x���ҷ�R�o�������\X�hL��Ǡ��Q!�;G�m6VFKI1R����R����a��Ճ)�l���;��*��C0jiom�y\�����Ly��f�J���oK����]8&+@U��D]t�@�٩��E�pU���P��dDnṡ�D'q��I�}磂a+7���*�Q�o��y=U�?W0K��k
�~iE�/�z��,\aH�z��6"��-���MD!�b�Iq�,l���܋. �A��P�r�A�q�|V١0�wC5�X�6)9m�G�!r�D�=Ώg��~e�(|���1FwDb�� ��}�SϚ��
=���Q��?i�o���k��6G?ٜg��m�1���$D +�W�I�DL��L��.��Gt���)��O�����WG���cQq_ؚ'���B� ����V��[��� �6?ߜf~���Pg�Q�v��^�j�t{e(���a�0�OM�j��6� ^4��6�LezY�����Mm�5��\�L�V�Y�\C�ǌG�|���08jEi^TB!vgcT%� ��:6I�y"�����c"���^���Kh�ɕe���U�
�l]�>D��"�O)��D�p�^�g��r��t��Ő��Ͳ+F�(�-[�$�y<A���m6y��N+�ڸԎ��)�Z��W�-c��N\�>���m�
7���฻�hϻ^�4@F��/�S`N���7�F�[�L�gR�^��x�U�$���UuZ֗�����$�+�w#�����3���V�t�V�l0t��cZa����b�tN�F��}+��B͋|c�v�u�Y���Mh��٢7Ϭ�j��)E�t�b��<���J�˦E�p�'O����V|�m���[s��~�1Vn�Z���)v�n2���	���G��c#��Wy�E7Kv� �p��:�hRXꞓ��z�o�m.�K[�h`ke����FFm}H(<�A6�y=��@�p��f�v�*l8�޸�7N1b�����p��XB��Z����
fܨ�lq΢�:����&e�\���:���i�ER���R�~-�'q�h�=���R^��48c��EY�'�wv��oj�V���� {�(�۔���[}�B�����VF@%g]k�lm�� W��^U�YZ>��A��������7�����"D++�����=����`͆�TE�%_�4����E�]���'S��TWL$	���5Mfj<�e�ܠx�M�;�
�a�4��5�]^B�h�rf/�sT�N��p�C���� fnնI��[��8�
:�0lq��nj�4��n2�eC��K�%��˸�Oh˫F�q��]�t��^��q�m���U,օ�GJ�Xpb'�@��O��,��ۍ���O���t*�KK��,��!�5��e��'c�`F�Ӛ�qN$-U��w�n7�hN�'G��<�(ba��oǝ��tP5n��W��Ig�$�買♫3��˒~A�I�رB}XQ�n
���iya藛��{����X��O4B��r��~z�4�J��,O7�9BP���: K,&K�6;tU�&�wY�h�'w���av�����ha>����쫟'7�d��H���=��^)�B�=������WtfvO��?�� M�[���X?�
ys0�7k{� �7��j�������̕�S��i��!��=�$"��o:�f��WѾ4���^�tgP�~�E�cm�>�{a�F��{�UI� �qq��7I��:��,#"��5����7��<�����Բ�$پ̃*F�/cw�v��}Lx�:�>G�#����,�Dhŝ�o"s�{�&�`�Зg���`EI?�s�Tu�Q(�И�z ��;�G���E:V�N�%���JB����|=~S0
�V��;0��!�i0�v{�8г�z� [�_�gr�W�y��Q<��r��<�#��K�����B����2��PGD�uê�O�PVƳ`���B_�"ZB���Ί$��}�*��䇧-��Ʈ-�N�����fkct������}z�����>qV����e23�Dd�{�]���s�a"�|q@��l�5��V�}O�P���O)H����_d��r�r,�77��8�1 ��b��"|��&�
n��Oղ��˷�;��[/�4J���Us͂&	T�~~����`�R�7/o�Q0VV�)�,a��}�qɐ��9�
����_K���h/��,�c���X���$1K;L���xG��>f��@P�Ӏ�Q�fIS���1�t�+G6R�ә�����v�@�C\��[��8:��1$EM�-�_%�w07������!�MrG^�j��<��T�	�����a�C�:��/��)d#���O-������޴�E��ˤs��E^W�N�)r(����˖]�{y���NQ0�F�|��:�i�IQ�	ݖ�j�bqB�\�q�I�حm�%�����b�Ud��9@`�O� ��b
w��& ���x��o���A�m�0�!!����C	&1�X'.U�H���~��j��BD���m�t?�J��u����֍D°��͈c�w�2����ㄏL<c5#�tg�������p&��$5!@�ΛQ �?��i���o�9D��w��a�Y:C&{�r�^�F�t��O�����sz���T���H
��6���g,����ZI��(����o?�@/����l��-1�lmY�Bb�v�;p��n��>;lP�o҆��wǻ9�r��e�C4DI{��+\������+�`��&y���s��2p2�T7��s'N�"�%|<
S�)[�#�)����i>�U/��#�:��,R���4�3��ʉjU�|
�/�p�[A��Y��pu� �@Q<)��p�f.�D�{�����j*�I9��{�%= ��w㓰�g�����'����=�gU����s�Nۢ;�j�o̐���Px�җ��.������/�%t��Y�I%���
%�~��"�B|�~r�>/��[�9m@��5�#8|k���(4$�ӡ�kv�'�X�#b3<�	�Z��9���'���a2%�2�d�޻�̍����wԲ�+մ��s���J�@��o�g��u���Vb�^��6�R��Q�v��S���40U���w9o��Y�q0�����O���Rn5w(���$-��,�։��}~Ɯ;�V�z5w��^
V6A�W,����t&�{��j����	�G�V��� ��8� ����r�X�B���Pz-�.��9ǘ��u���|� h���N9��YҵY'���:2+Gz�|�_8���"c�Y�_���h/�:�H��K��#��Ra~݀�0De�EtEN�����g��)]9�_��
�p
�@V��I.N~jgR����\"m4Oz�t&��]�;�}�=�Á�Ր����#J��1F��5��U�FEC�6��F���Cː�gQ<�n��$*QL�rPk&�Q��|Ú�<��sU��5�~�L7�9P)<[b���\މNӶ�lYk�]��!ɧ���\��9�:B���j3��`�o�ּ?��v�ڹ�6�>�0��"�=���e Fe�Ơ�6��Go��s
K�>�����6H[J�_��-y��Է�|�z�Wh�P�,�SkT�p)qЖL�a�~�@�8\Y��2֊��ɵ��Bg�i��<�w�Ml�0Sǟ^�ƾ��٥�&(e����]Y(<9�r��	�9_��{���d��=y�V�:��#B��|���u޽����'���m���>�6�U�|	�h�x/�!\%f�������%�r�
����������E�@VǆH���r\2�n5�c��ĸ��P�5�g��r�F��K懬��?��vm�	���@�_L�cD��d�yUv�'iLϣO�}R�z$��6�;�Hq���9L׸��~ˈ�t�`�섇^���`u����AW�z��&���uM��Z8*������[�M��;��g��Tw�42������y�`��V7j;�<����}����q���ْ�4�JiE�-k�s�:�j�^D�ë,rXQdGd�4@~tˆ�����dP��g) �o�I�
�֪����~��&D�g����a�?�L�Y%�oj��:w�-�= ���5(Π?�Cp:��7 �ӿuҒ�Z�İy�=��w$;z_dD��}��rN<-T�}N2w���G{T~w��0q�����o�+�lDڮ���u-���7n���n���/�ʹer��p�'5DsH�\�	�{�מ�TC���4o /��|^�$�Шߛ��Qa�n�7�`�-�5v׬3��TH�v2�pN;E���0 ��a����� Yd-�%���S=;c[*W���N,�Q=%FiUݮu��Qo&
��U�T��Ӕ߄��+��6jΣ�;+8b��ZF�f�f)&r��[��;i-ʤ�=������G�5��?3�'���n��&�{m�� �V��]���J�$i�;RP�F�/~�{ ��џ�YN����� q��P��L������R���}�˪u"W������*K��/�u�X���
���{��8�GP8Q�ؤ\�=V)�	s���$��hh��}�5������1���}���TxD5S�ʗJ������4��F|���y�h y�+|J�c��[�.x��l� ��۴�ܺE�����p�DtF�A B�H��[�J�u���H���jsX~cr|?������	߉�f�sS�z�c��	����:Y��E��]�@g�B�����י�E/�I|��ᵧ�
��b��g@�sV���7wm�ե��i�$ϥL���b*߄��*������Z�<~����%���5��r��������G�jR��b���H=1�ͤ�%2����k�yr@D(�;�Rj�+�������wwn�/��@5S�Q�Qj���2���ve2y	f�Fߞ��p"h5���]L������Xa�!� �=�Q��,����"4�]l�=���@��Z�F��~�K��:�O��_U<��C�Vj�E7#�{Y5����Ǆ�yS.�:�Ṕo��G̤���\��*�� 45�-tY��UI��ݛ��j�͡r��_��?��:t��6�Ɍ7���0�y��ߑm>@&�3�cUbλj�7_m�
Cg�$0М�ц�㛵�B��9}�>*c��$��Ԣ��]�5����<�e�v &mB'�}�ا��p�>��a���ϼ"~��fҀ��%�/�3����N� �N,l���}~re�V<SfE%86zp'�@뾗`��p��}�ו���jsȼ���=0���Z�o���-�����!r�%b� 0�-��`]-#�Є�n�7�vt��}f��?���t�m3�����Z����F��/��������������2�\:8O��ڀAWKz;%������Y�z�A����z�-���4@����ۆ�mT�Å���)�~X'6>�qIt}Cђ�m~ㄟIW�`��3k�`r�{��������bOuXG��.M��~HΩ��?A1���(�&�"Ei��1y�O�2�	D��K"@�M+����8�%z���r I䒁�ǹl)\��Σ�����o,y%{����k%�)*	 So�[w̌P��`�s1��\��u��Kz�K��*Z�V0��BK�w-i��<�\���0��7��=|��}^r�s?Ꮶ�W���Q�����{�=s��ш��R�b���XmNg�ub��C���dm�@�������iHcx�M�]��".�`M�����4�PFt�Q�ޟl����YR�@����l���й4��N�~N�_8\��]������r�l�di��?Mǀ]��݊��I��.8v���I���w�����@I���A��ݘ �E�D��{���P�p(��B!��$��:�R��h)]/��s�7�[o=����w�� fa�'�v����PN����*��q`���Up5:i��uD���j:pJ�Ӟ��*���D�6z��`�gD���'?��U�gI��C�ۉ�+��䘠6n���K�%��i���` b�}���.�H0���i��o�ʢ:�c�g��߫�P�ν3g�6�q����;i,��={���s|�IEa�l�=T���Ϝ��w�4�	^l�;ܾ@+�=�����8�a��(��/�B�#.MB�k�&1�o3\��Cqp�]MD���'@+�_ҕ˱M6%��x������*%��~�'�?�f�X�P25����қ�͔+>�0�KDL8%���Q�P�K���O�*�'ee�r�h�8Ⳟ��}�a�s*Q}�/�H���ھ�2�?�UcM�P/i�HD��(u��V\�ӊ�K1c�&����
��\�@6��I�alM9���{P ��<��¯x����x��x`�:�@�{��!�,���<�ϳ�e��XZ�BUP�:I���-�0��d��in��R/��@6��[��@܊�]��l*�s< �Цhq�=�">���G��v���d���~*�Yt��+[��ᰖ�zۻ�+�����T�+�˜2�!2E>lr��pV ɼ��V��J�<h�T��WsL�1R�)���$r�PCAygOQ��^�t�qy3�Na�Ն@-����<�g����^�0�
5<�@��6C�D�4,�&[��J�ALYO��V*�׵%��F��K{��<��`1D8�\S
@*;଻����k~(q.L�ag�n�K|찏�!���[�m,���մ۳>Yt��u	��*z��Fg�̀��p1�e0ٜs���S���yl�k��k�Q�l�΃�d�j�C�#�l�X
dC�m}6�ץ������cj����\�tӻ��^�b=mYHI�E�2xӋٲ@����0�:n�"~���bi����H�W+����}���e�����H����{܃�N�J�/obr�K�܌j;q���ki�%��r���ߣ��Ӎ����l��Z�q̲6g ]hZ$��o��ӊ �m7pX0TB��լ���A�z�T� �A�YLGڪ+?���1�=b��K���P	z���+�`+d�GX��'�h�kl5����F�E�����"�rv(�D�
�yԲ��;ρ��w��`�β�թW�M�r����,��wc��"��\s�A��m��d�D���1R�-/3.�����n����ĎvA��5$��5ߵn���tx��ނ$�_b��Y1��*5���K�(���R�RX*߂؝�$~k��2�o�^��Ǉ�	N�^�LZ�/+?1Q�J��$䛘�HXQa�^߲Gb��V�@�*!*ȫ��/׺r��p���M��BC��#y`,/6k^8RX�1�mPxH�t"�'ax:{�������R0%rSn*��� 8�![V�٥c�h�{�3�z�T�S]�I�cA]������8z7��[�<[&�F�+9��	Ԅ��K��o��K��2���/���YO��N�M�ƌ3��F�`�p�x��E�(�n���������U���a\����Q��Hb���8�m:"�0H���Í2�:J�a�M�r�Ųc��b�/h���!bG�Ɲ�m�#�w�Sj̩���~nk��`�k0���µ���Y��&����qi���9�g
��Lی���U̎a٘g�t�{�&���׉9���_ݑ,��\�]���E9L��Ӹ���L@��2������/=h ���S��4���g>y��@��m,�����8(Gċ���90��؅���.�.��»�� +J��J3�^��Dúau0Y�v;	��.�g#ydmx֩<P�u�	.��ڏhu&
8��~��U�Z�����p�tN_ж[A�������:��C<2��#�x�
y��pkd���FBj�CMv���{�� ��T鄤�&�B��_�$���_���.n�C��%$@>���[��x8�YeoL����	�qwC�$Y���I;�<(Я�B��]M����ق�]���%����2y)W��k{"���Q�C���<��J�)�ZgQ�y`�֕@�8M#���$���=&P���v� {�]jUO�i���^�����'���8��dQاqڎ���:X�`9��|�+������6�H�P�aҘ࿦�^����?z~��Wm�'jX6���Ucga��)�_JS��k�DI��@8�pk"}����� ��pv;�P�?����Y'gHr���T!��e�o�l��]��^�kt?���c�kx�_�C�����#�3�ϣ��`JZd�ō(���`źf��HV&����̨����K�1�g k�)aW�]#��*$ޯe �̿n �i�;���;Jiu{�2�^6J�,%��N<���4�^̊WB�Ǒ��w�)4�����T�g����5deg�q=9���2]��]�����`��Pyġ��NZ�b�����d�{i[ʯ���a���sd�"�/���ѱ���EǙ˱�b�6P��}[%Ľ�)`A�������Q�&���8a�8��MȪ����K��~E٬�fu#I��?gc$?l>�W�\k�����.�"�m�w����2M$�~��ً�h*<�^����W���A�#�\4u����X�6���BM�����~@2A��+�U�����җ!�"#j�GE�EQ7�ҥ��7c	�z�*r�XD$T
љbr\}��@��*�|��'�pG�WL?�D�σQ��(�n���h��˼�����a,�@�)ݡ�x���9t�g� �G�|E�S*X(H���z���:<�u6@�����(�������K��Pȶ[�a��d���&��1�=�}���Be�e���d�n8��SҸW�Ƥ���s�������W�=/UM� G�,k����xQ�o]رdY%���i`-��U�<���{az���6K��N��"N�BX�#��2�mrb�xq]{���d:��`�$�K]�iA\s`�d~����1�A�D���*!�����'LPHl�P�I����Vy���!�p�I����Y�sѮ�[�A�c��%WHfB(x վ}p��}�Sl�X���Y�=FX�%�J%,6^���` �?�\	B��.�_t
u+�U�W�4��iԐ81��R�&�@������W�Dl+�v�"��q����`*<�*pz��O���� �'(`�-��{#�KyB�~(�ǆ�}1��˱"���fZ���9�u�
[H�]+�s{��P�3�h�쾺�3x��J=�&kz5��.E?��ն�վ�������
7M��^.���0v�7-�F����^j4MF��eg"�w�>Sݬ�*fc�1�$Mw̼d�G�T�du�@n3��rz��K�s?�7j�$6_<єo)�<�<�_(�m�>=��Jwn��m�>k�і��z%���2�y�9y�FTj#;�*�$7�HB͊s���wa��d-iE��2�<>��{�|�%R�X��x#��~ݙy�B�6�"G�\��)�?݇��������
��1X�~Y�W�����+���H������ eR|<WL{O_�/gIܿ�skpj���-ߕ��:_�=�ErCrt���e8�H'�C��o�i!#u�3IǞ�jC�YiR��Z�o�ˋ�(�~2չ{@�-xe�Ve� ݚ���r/㜳���z��n�6y��+^+�W��'M���w_��w�=&u&ys�bs@Hh@�8�K�����_ �d]�N�uo,r,���*(�VKj?Ak3e���ŽE5:�DG�w���W���m�_0۷}�N����Le� ��މ5�A*���ݖ8ڼ.Â�K�����e����T����bՑ�O��]7�$��h��D�Ik]�ʹ\�fT��y���,��WQ~��H�i���k��"���װm#(2?X�α��ZcshӠX���-�fz;�zX���I�KE�dhݓ`*�}��?��_�Ģ��C^C�W�~sQ�+��!��T0�o�T6Iz���c��~䯽W���?:��մ�5�%�:䷵J��f,�*r���.Y�rԹ޳s1O�e�׀a�x�HB���0|wV��jЧ<��p�X������cĨ�ףm��Q_�7E���̙nE&��B�Nk�B	�Ŵ��V�Mn	�Z@h�A-����١�=d�g�Ћ�*�������'��c��]t�	�_�1L�7���a:4�X�=��R7�}0>N�Yi���ͅ���u�t�z�&�ۻͥ�`Va���ΐvC����.�3�k"f~�=V��Dx��(��V��~l0n&���A��_���),��[��]��k��N��,t�Ȍ�i�f���ar��g�y�w�ᕍ��X����>
�ݮ��Oy¯�;W9��Ĩj���R�Ć� b��}&��0�)f^V��Zji����/�Lɖ��m�*�N�0uQL�ڃx	iB_/r+���H@�ɰ�O>aOk�6l�U�[ָ�"*����$���%�+H�M�~Pu	�	���t�2v�\^��^��r�}�e/�GU@jx@��Ӣ;�*h�8�I�u�A*�B����S#-�<��<�1�Ӥ�?�^w��������u�x9;%��Wu�!����-7ͽ>2�����n�L-O�翝 �ܜn�XBO�a*���!ف��S���_��#��x�����g��3k��+z�(Aɑ�sc[S+�S����2���x��wO2Dhċ�Ds��E�E���=:s�;�?߹Qkc�F��8���m<�vG-R*��"ĺ=oRi*��p��	���!b"x\�_��;��L�����	;��E�ej��"��|U���4���d��A���`l���u���y,99&�����ϔW`;�(��Z�s�i'��å�O0�%y|� ln�2&~�mrܖ�襃�p䂜��h[	mzk?�bfFf�[�˩3���"x�5<� =�t[�˖�i��vk@Ds�L�Q����7k�{s|\���8f
�?����@���A����9I8!�*�6rb��A��`(�P�5��w���������UPk��\�@@f��Z@ �G�qƽ3�5U8��*��^�Dܝ��}�A�
�I8?ۊ<$|��>�F񣝤+��X4�y�����6����{���<ɘ%$��lj����+�pw��f�ֻ�JD���gC�oV8W s,��x'�~�$�-ȥ�I��軷��G�t�ܦ�N�����A��̈́���郚(s�X�G�c�OՏ��l/570�X���J}�F:�KI:b��ޯ�����"!.�*^����{�w���@��v�[��5�"bf����H��P��P
�� ���~x$�$�g��9�=��+��~�E�]+�3Q�\>%��ڼ7h�n�X��U@�V���8��G޽{���������4q���,s���r���;�;m��rA�n#�ZT��
`4�{..����=pZ>�I�i�������ґ�Oߡ�"�ɯA�*P�HI���0�驡%Rx���%X��/G�$~m�u����o�`|E�kbE|�H,�6�-�/͓˫�����jQ���/������Fy[���e� 6��Yu���⥌m�c�Hs�;�yR�sG��HY�ŐtV�����=�dN(�'��+�������p;	��y�����9ix����8��g�9��^��ר6�w�:}^O
��n���=�~�^�~T'z��6Z~��^�Q��8����e�#K(�d&TfP�ӎ�[��\<�x��ׂer�A����$P�Pa����m���şp��49_�W�&2����ޔ("� Ԉ-�+�O�{_UK�(t�3���(�Įl�eĩ���q$M�#�۝y	G���`����G��%xCUk�"������A��/;m�3c���-�CK\w�X�.�!e�����5M��Ut��Ɏ�� C�$iO�b�L��D���q���4���_� ��n����0��rs�%�l'�^����bu�J��m��9�w���,f�r�=ȿ
y�h���w�.�+�h�#G�䇭�FP{Qt���rF�������`џ\�+��هa�BVl�e���&�^.�D���]��\�$��yA4r=<�-�����8N��
}���o���D�>s2��]��}<����0��a��@YaAc��D�-~��e�������Z�+,0�|!j��<cD�<�j-���{5Ye���Z����8�i͋P�����w;;�7[�#ܐ�����_j���/���@@�j`ƙ��Ֆ� )^8V�@JO�E�/!��?��@+��������bOm�<����*�[���b��'Om��"~�i�I�H|����)J S�c��L���?¹�[[si,jQmNk�hK��ǜ'�����d�eS|&�"��yg����on��F�~zs����$�"��u�ޔ�Ÿ���~����J�"!6��bo!$]�o^�:4�z�S�vh�ޡ}�P�(��u3�����>���w#D �Q,�.�Cz���s�*�ԦrŜi?1̥����UP,Q����ZPfȳ�|�Г,*���X�j��.99�ߑP:��8±;��R�u��	�b���Ǻ�$$��*�sH�������0u��~_d3�5@��k���IY�e��s]�(汍l�����bn��1�1�wl�]��� ���1ff�3�W3g���R�Uм���z�r��ڱ���q6����G��TRنK��>�8,�	�'r˂�;��޾�!�Uk��	�W>���$"u�:�|5�9��k"���_�L�p��a�BM�{�s�w�O.�e��W��-Ie��<%���(�o�������.|"�ʜ���nA�$w�6��f|�z��P3]@Nm���s�f�8�b/�:�x�o
q��'s�����6Q��JPƙ(�)3�{ ���i���]���
M[�������}25610�eR�˺5[��cc��q��~w�Gn`s`$�z��'[��b7�����KL$���	O剆=P�B�����	M Te���-ީ��=�]<��8 �O�	�͑�Hٟ�^�����?��;�Ы���_J:�γ�]=��L�PZ��5�'t��!���m,5�o907&���F�jQ��W����)"��<a!��3�����2Nz�;�D���T:w����2��3o���º2�KZ%l@[m�R�A�e��+�!�g��#�w���͔Ru�j��}Y���"�kY� �M=j��4l��͔Bpk|�oj�����v��kMԂ!|��U�~�GP�0��#~�u?�¨����p=�I�#v�А��P��Xg�����k<��k��,���Bց�b��{���x*��7�r{7ʶҒN�@RD���I`S�{-յy�!�Q�{;�����(=�!�D�&u0���m�n�nZ$RL��Յ��AU���G���R�����|����z�:ӥ~8qzDa
S05�4��5񨺵����܌��Aw��U� �u;�$O=��}�ɕ��A�nY�|��q �Q�;Xd
,�z�$��a���X8\�j�ۻ�����m*zV�K=�+vS�����F'L���E��jq���:�\g�������wf:�<���Wm=hꀡ�]x b�ƥ�����"MO���G�'i &G�b�mť%NL���va��Mĥ��9�v4p��*k�D6����bU,׼����|��0�MC�ZYr>[P��$�a_�%��:�h�䪊ME�M���"�
�ߓ}��j���O�	�f�8���"���B��ę�b��M�lMl�A��ex���6��낚?*�hy��� �>I;�\6�����Aq�(.x��ğ|� =M�Wt�y�+=f�M)L�*�?M�!�� 
��Y�OJE�������T��a_�S���c~���sZ��ؗ ���� 8�"%���;D+������v�L�gk�imA�<�5wګ&;�7��%z ��\�.�N).�d�[���9�re�+�����R�(Ul�Z�:p� ��eq�?|w�?5H���J=�#�T?��P8�1 ��HCZ�J��^�U����"��y�ȡH�D?C�4sn����F6V�^�@�Y�8���3����N�Xu��+�ϥʠ�wUq�&|��c�^���7$��aa�J�P�٨�˖�[���C�'���h|�:t��t���boW`僑~x[�� ���[\�u롒�G7z��'�� ^x��6m�~G�n�v]�	"t?�
�J�!kk����~�=Iʶ���Z��(��ͳ)X�b�F�"��:d��2
(
���JHk���
��T9=�X�>0�w�T�G�ۅ'��D���D�(����'����,V�#~FxT�@���a���	��ո���3~�ԎP/Χ���.��v��$��J��f�E�&:�'/k�s|5n��+,V*�Di������m_�у���).d�ro�k�E@��$�-n�����U��_��a�O�ʎ��lY��Y_��Π�!�H;���=�
p��;�5v��&*I�v����<a��
MO<��c��ꗼ+�I8�^�7�(H��E�J�8�ݾs�	��f�Q��V5��M���ȪV������]W1,c�I~�pTkg@��I�~�!Rny��:%�s���
��M{�V�#��������*��,���W w���}�h+�u�����2]�ԗ�m�3¦�?����| �@��	��3���}gH�(�lN�#���87�{T�zn3P�*�H{�(r�EF�Sw*�P�؉�+I�*Tt>�wtI��[�+���9��BtȂ[��	Y��3N&���IJ�ec������<yi�}.!��`z��%�Cy�o5ǚ^G�+�@i$1�?1+7#cqڪ���MW�FqZN�l�����_�2k5A+���������4��	�R@��,�LR�Z�n���]�䧯.�c����4�j��JvE�y�!j���U�����$s��l_�p�A���i���
(dP7	��\�d��� ��K���g@���Ƶ�:(�nX�n2�"1��7��]Qh⚊�ۜc�nW���%r�vO0�h�x27�=YW��;���H؄�]�ހ~|MY4�mmV:B��*2O�~і�6�G	1D�{�V;��t+��3y�ʮ���ef���a�gZDA�1��h���7�z�C����mU��Z�[S������{us���W��z�@�F@��j�a���#i�<���A�'z����C�Y�9�$O�(r��2b����"�3�E.iOZT�>">T.#�+�����.�+L]
:]�������>o��b�k1�������Z`���J�<&e�lK�<K���J����8��Oɘ�=C<�-i��Yl�zi_]~T��+ڣ���P�C���eъN0B�F��Ÿ������o� ��<��O|�:�����Xq,f"f�'a	�:G����[�������7^r�&3���
�aQ�ު���p=o�ի����/)��w�U˱E�9�S�2ԍ~`V�y��'F��K����P��}ڎ�}=z|l�C^���o`0�>%����^p"��&����I��&�yƜ�,H�+ T���S�-�M�$���w&�R��1�m������G<������I3�¶�J	ٶ��(���ȑfz>��o��[y�g
��ؿ�h�Y0,H�3�,�(S���ʩ��D ��J�wȪ����u�Qx'5G�PF��C�Z���i!�X)��.鶊dj#�d�\7(�1��ͧ�;� �J4��\H��qj2��y��z�/�&�/���t&e�W�]4����jt/w���N�@��Y�_�/ɸ�_�%�3�O��úw���������8kZ�2?g��K֔f���N��s=4X+3��Ë�W]K0���2ȝ��½z��`�J�a��[��� �S;�8�ƭ�fI�ވV�ß�o*��h������`�zt��/���]�=�� ��2{T�ݛ)��ΕhŲ��0
"R����O��P�/17*ky�4�4a�ݳ�B��u3P�9L `r�mj�5}��{�$?"��;�۝r����Ԓ�i:��;�-�����	{��k^�[��`)� � ���$QBj�n���'��s"��p1����x��+��#��)��B��wQ�FI �Nј�T��֐noo�$�0��+R��Ϥ�B.�����L^���%�B��r�$(E�%�|G*�Y>K�F�S�e�e�X���v�o�hdPOK%�
�p�?:����t¶��_�����A<z� �I�G7��j0	��^_���;�_�a�N�k!&��+P���A0/�|*�]��������Sr�)��=Pf��'R��@�G��+Il�8E��.��f*Ӆ��Mi�oĘ;�;?�*`��R��>,j��X���-�׵�����2����lb�F�0��$8�0Wth��� ��ה�t�R������fSmS���`�9�n�i;&d�@2-�˦cck��-�Ppld֙�S���b*h�Z��@H��7L�H_�}=fl���]rn���1�v8}@
�א���\�B�k��Vb,�g��XUC��_�I��6��҄2ó�}��Z�S%Z�yʳc��c��]��o�a٨(Gatx��~���U�Y����?����x�>���vT��(B|� �??yM^��̺�͹��D{�K���ɨ��2���X��  $�L�_�R>G��Ee�،o�w��p)LX�k\�~��O�Ş��G¼��vl� ���1Ht����ާ`�h�_htB�衮'#������Ĳ�WZ�&u��[����]�(�5WˢO�E-)j��i;� V���䂙�/��[�����͜���=ɳ���;��8�dx2�><�!
2�۰i�"��'o�m_2##������ĵ�	:����~\���Fѧ6��m�c�����I������?�w�r�e��0�/>�?��6���1�m��0�5��	�~�	W� ��RD��b}5���qi�m��M���5�(��b�����N.4،�<?z�u�YP(��!>��w����᠙v��q��[���q�`�w{3K�@B"�_��h�hh�1 t=R�
�7���y.�Aq���<�Q&	�,F�Z�I�;�du��!n����3����o���i9��C��/r�؁�ee*���>�D�엮�_���:�ЈI��!b;}���j��M��K ������&+�U�$��q���|�QA�k��,b��Q}:[c�;��]����!<|�Q��8��t�;Ϙc�ۄt���C&��\�Ef9j���)k�OI����f= �2��ۭ�b����xz3V@��>�P�S��b��{v�OZy��6Hr��"A]<����F0�cGӆ1QY�o19qU�z,Ώ�(8Zfe�ż�=���j�x<U��'%[�5�6�oa@�y8��7 ���@1�IL��*0e7�itD�����:���Vm�e���&�ZVȆ��T�����!\��8;�.���2�����f�Q�z(\�^���g{��7��£D�|*qc��.l�����Yr�m��Gp�$��4�ց�߀��Q���G�$�\{W�y1X	�f�`���"�G���F�M���-���ŀ�5���a�x_�h��Nw?��m��j&G�����̀^��~����)����T�ۙ�k{m�����x��q�^M�]�M�{ ��Z�*h�Р�R��rՙ߸U�{�#k�#jz��ɫ��m��Z�
�R�sA'��gԼpUCؿ+i1������?״�!i��<�zub� l�J�VZ��sM"���y�Т��qf�1/���KG{�?H�l��Y��[��ea���,^���^��ʰ%)	{^����:7*4׋��!�A=�)�s�(Z�5�3>.�iR��׉�F��W2�T��˵P,~3��n_�Q�E�$��d�k���Z��C�N��򤭆����/!ztv/:GM��x��r���3|]�t��軘�B��S�p��ـ���ֱ]��	?�#e��*u����tPBj$��F��Ck�8t�Xf{?��X!/�o+�/�����7A4~DD!-�G��pH�]$�-��R�&�7)���!�+LR��Fk#��{�m�� �ů3A��D�ȹ.�ΐ��d��nX��]
�m|mqQ��%��VQDq#�؅��)����\,�[(q��t�-Ϗوe129oFo������N�b��f�|g(��,I�i����h6���do~ŝ�zĖ\=�rO�$Q428Mك�{��)�t��S�Z[���b�B8��G�	�
P��aUsi�v��V��u��N�2#��?O]6r�UuC��hb.�u6����~���^�}@�