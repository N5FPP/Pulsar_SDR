��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY����B|Y�9��c1��p:������`z�a�)��;�D$MW�
*�^`!npGUQ�8�wټF�)��`Q�=��t����6�R��w�������R񓹚�μ�qm��M&F���s�rHkHզưI��f��ax�����D�r-��?e��{�NT����ٰ{�E��<$�xCѱ�M�x����e]��$��n��2}g��b^[���B!ѿ��cΤ&˟)7M��I�!�p�F��R�Iy��iҾ+�$���a�����"U��j@�8���Bh|Bgɩ�c+���������|���'��=b��y�Z[%Z[ǈ}��P��%�ws����s�\U�|!�����v��<���7Hs�5�3.$l�сӃ8�T���Z��H��&6b��mX�R�
�ҍ��{����V!��Xݦ
��ɳ0i��M��ǧ�ԏ����dJ��p~����V�9yD^J�P����K�&��1?9���G�J������>xvu1D����c����pm�?02���L�p' $��k��g��B]�6*.�z���\�q˦Ɓi8����:F�8$�X[�	�-?ky�� ��m	��F+Ń��&����Ilj��9J�o"��e￯a+>�f����:ݚ��b
l��L�)4b��w�K�cxH3��j����q^Pm����F���S�pR`���
E��h(�P��7Pp2�4���O���0�v�R��/lW�|�d�X_�l�>jU��I2f�j BL(��k����
��^���AA6���:�()���G����(���;�CJ�S3��p��Q�?�˶��k9�:ԟ�#����H�&����R <ϊR�)噂����L�t��+���b@�l�oʐ1�m{�+Bu�w�l2SIǅDz��8�5��pr�ɬf�ə�-��&/��+2Ca�auig4���LO�S+D���v[�g
C�i��N�&+�bC� B�c'�N���M"����w�\�R�X��4)�\�}\�7��}�3$\�8�=�R�,�f�?��+��ҹ(���#ND�`J���Yd���?-��ͥTݡ�V�� �iR���˒���RyX�3k�� ޔy3 �p����(.L�0�$C�Ɓ������V�A�2+�e'WY�L�λ��_�k����W��5���[7�ؠ��s�7�x�[�y��������W���r��ߛ�2)�v��;��:�K�.j����!��$��hF�z-n� \;���[��Pߦ"/�� )�a�ۊ���A˦��0y�3zT�-��.4lDiT����$|<IwbHԼ���M����WYH��ˬ_��%8��I։s��j��M�ad����0�A�hO�P��wr�e�ZfE@����gt���DOͷK_���7�z�'l�t����L[4���'	��>�F� &����j|�a�0+1�����t�!��|q4i�`A��9���~`��Q"�CEKTM2���n�Q^����|i9s3M?��_��5D�����`FN}b�C/9R��E���^��Gձ��W���$�3�=a�a�R� �#�s�ǞYP�a����=.ʏ>��g�fMX�J>a��*q��=	�7?�ܿ�3(�X�/!�7ٝD���\�F�>�&����\^���ş�"c�QU�b�������29��%^�x'�eI��N��M����w�&Mo������Z�ǔr}�5Hm�7^�R�Z��u!���	�����ܥY˭:�3��[�a� ����,��kg� �&�9�5m���'�Qg�=�T�Dn����Y0�=KIc�����)��7�����aA����/�'��)5)d��NL���:��ɸ@^� �G�����bu�M��%��eo&�M��m�c#�r���::�����ƀ[��'A;�.�s�2�j�6$�Vڵ�\i�FFHR���gdyx��q�X�;����Fwؿ\"��)\�.��74��ًe��X�\i�֧�DK{���y`� �ԛk�ֿ��5�K#�RK.FY��Z����u��j|.���NL�pB`׏a;�i���au����T�5`u~\��
�F�c��u���%|�	[�2���P>�
T�d��L�2�����2�W� z*]Pr��|�qk�T#�]mpK	Η��p�����ZƜ/���glJ̐�!�f�<�n�Rqŕ<Z~gn���F�ŷ�C�d�?��"�p�+�t����O)�M�2�XƝ/9m���:�N
�r�d+��"j�WAw롞�U��g�?ҩVx[ٔIƢ��Xɱf��7�)��ƁSIm�)���G�p�'�+)�dk�3<�^~��������
W<IZ��n-f��נ��}*��ҙ&G��AQ���j����C�z����[ՑG�Zj�t�xr�z��y	Y�5i[�:�':W��3S�[��	a)H<��_FW�`��Ы����%�~.K?�-�eV����{*��w�r�П���^�J�j�� �C���uiY	HMk����Ԧ<+�������$%�#0H�IP{^��JC��Qƒ����=g�x�#���kb�	��IZ��;�Rz���Ƙ�x�P੹��QN%pqh7e$�a��g؉8��)�;K�71�*چ1W���C$zh��dˉHn�bk1bxX��,w�N�籃>b�<�e�W���G� 7q�e�;����X���k/�`h�l�ʌ�O�p�w3	���u�:����5A���R �!vE��5�ߘSZU�ŉ��'�L�ˉHJ�͸n2�8�����ȟ�&�B���t�sY!��%)��$�e���j_�v΁�#�wVb� P�S�?J��
6Ŏ
��|���w��J�˪�I�h�*�ڞT �jd8j^��437��c��^6�ڰ>\��]��B]ss�-���N�_�]��I��R�*ɦ>%��k�0��pD~t�*��ԝ�(��	���(oR�(f�j�q�k�Ο�M�=-������h��T�j�k}�R���G�sZ�*N�������2���]�OÇC�go��3�z?� |��`N��2���zG��z��~�����~	yw����t�Ɗv���)r� �%ӊ=�.�86.�c�3�	Gb=��K��*���9	ܫ����u�ݙ,;��	�G�r����Y	^�Va�����)G%˚��E3�������<��Iwi8�����13+JV:�z"o��*�70^�q�'��vx��e%tw.ֽ�$��&QFNW3�V����(���zm�3xn��[�9
W��<��$HSx�7���ʶ>���_�p�Frsk��㳓|z�t唹
����n�+��c	k���j)V^���(���)�w�|
�$L�Tb�_��u�Z7a�5�4����<p����J�W�uڭm�P.!gʚ����e
��d
�����>U�ʶ�����`��̌Q,���j��Ƴ�H��˛o�r�(�ߟ�Sm>���ȋ��9t�N[��J������Bw�Wn�c�l2ά!�6IUqwy�Rq��A���@����J�/F���)��}D�c��W��o�qAЁ�����ޚu�˘��CÎ^ac�r�Gt{lҏ\]�[���m.D�k��Aٚ���	���p��ƶH��e����ҭ�s*$��f�����b$: ��Ft���h�2��i	�E͊9����[�{@d5ئ]�����g("0�ɝ�?��)�-H�J)����-h�-�⹆L�z�U��
�F6�o��hf�¯+IYNc6f3�j��/D��A��f��-��9k=�7~pJV��c_��=�zr���l8�<�W6ݒ88;�^��*�a� �CI�R�k`(��3WasYo��-!���|C�>�nF��m����~D�C�|C��{�t==�iPu�z"'�.��?�����7PI�����@����%��d-P�`]�em#�<
{Ɨ��씤ݚ�y|�|7\��0���+Ž�/G���Ƚ�f�#�[����42TF�G���tӫS���暶:�s%[�*��Gu��֛��s+z��ꄧ��Cul�hy����蟔�
ΤW]���}f�Ѐ(�.tĘCl_�1���s߆�p�W3�뚡r��.0m^�CQ 5#���9�Q��T��R�oQ�!�]���غ�(�͝��\W�*�>��ʁr#���.��������`\A�w��#�,�
�5�Ґ^�JܥI~��p�����9�0>���Ɛ	��=!d�B�"�'w&SS2�ɾo���%o�Jb-���E��I-��sOe!����O��w�p��Ŏ� Ԭ�!+�2$����NA�M���qDU�
�ed߁�����=����P�Y��)7��8�� ���
̧
�$����բ�n]�Ӌb��d�T��{�B"f\��:Sn�h��/D#|qK^�/S�de?�IZpD9�.hl�S��w����c�5D�E�h�+��^��,�\�À�!|��*���y�6�ȳ.�;u,fշY�^�\���^�Q���J>� �xq8j�����m�WTL�V����a��mV:D�q�"Ei_	њ����5G��K"d,!#��M�x�4_��q���v�i�r~�R9��J'`w�<Mʠ}�x�jV��&-U�۠�Ut�P�R�?�j>ij���7����]LL��(96�a˴�L�{T\9�3�</_�O�i�)9@�ɀ���OC������f�����.De��t�Az�૪��R1|0��9D��nvy"� v�|�,�D��(M0�''7%[��%�1Z˻���DY��{�K�>3᳧	��ȓϊV�1�=���H���
<(&��]��$vq^w�E[�,�|�������q4,OC�g�]�Lڑ�ýA�������6�,C�\A�e�|
R�g�l����6|.�r"��,4W��&��>���w8�J�:�y�ƻ_x�5�w_�6���!��z�U���p�����}b��^F_j~t���%bf�r� ���ZNo����@��Wr`����c�]���S�hA�g�jT�p���1�4��2�������Ì��U�r*��a�~�y�A4�����3`�yzfּAK����J*�-�{������$dK%��SYڤ�A� 2��<Y����])�=�25��&N}���!�QeX	�~(�V{�e�u'e��;�bc�k�eu�iΤ�Q~�~�!����L����6琫Z|s �e�2���+��f��(s3���%$�0�X�Vz"4�K��/�4û��v�Ƨ� ��cˍ��?��zZIi�B(>ƍ�����R��·<uZ�s��BU��Z���ŋ\n�f�+�#�[����X׈V�|��w��3���N\���t�n+���z�c��	�:	�)C��H�`;��^��-6Hk��!$'����QB�]:򺭗[�|}��l�{��#�DI��@�2�S���j��綼w�w%s�g��N�H�n��Fdz�FxMXc���,~11�K�-���sYwT�5�q=?�ES��2G'�5�D�ߘ#�����m��H��=
�'xWyyi�"p�� �~�" �HVy�O�SBVN�~_���=�a����y{��b*��9����}��4X�S�MI�N};�g�A�.\����\���x���HQ6[���NΞ�W��8'���h��`u�>jó�GΤ�߱�®+
9l�8jx&/=�T�5WM]bZ����y��Ұnu��h�l/S#�b�	�-�~��^������o`�}<��Ӗ�,��X��C�;�Q�U��)�M!�hH=R�d敎��'Lp�v7��fA5����i���\ꂋ��=�fg[�k��kW� *����;J��lD�ϛ?�1���LIF1䊛T;���k��A~^�U����^�\��ةlڗt����{��6΀a��ݢ-}̧�Rq���W��� J3� ��Ӌ�⹬&-����/z����(�U�WɀpENӠ��萪J1'��Ko�6MX������J5�5S�t׼b�Tm����{1U�(���x�E!��ik���cq�l��<�Wf��*],�Z(vIA:��Kj $m�,UD��ku�]fs䈃)� ��^F�$|�*埛�2;�1\�Lb�3t�����'��p
���jȒ�X�ΰA6&���8�f�=g�wtU�+�vS��,5�� �~A�R�����Wn�p)���~�7B�� 3>A��_{J�7�����B���S�M�w���$#�H��c�p��q�V@�/~�̪�9��;E�[����aTe�˸��"w��Ú���w�D�M
�df�q@A��>? Q��sf0�yp"`�vJ ���Ξ��/ד����DǤ���i��]ܚ<ķd/a�������
���2���J.+ϵh¡6�U��?�'��X\�H�Ӳ!_i���0�U@�Y>��#n��� �+��4�pz+X���}G!u��_11폥���/��5rh����P *q@]�m���dѐ~V���Q�XbY���N��98!9-����-�ɪ9�E0��z��J#��LL;�O'4t˓�Y���K����8���6Lu��n3�ʑ�:K	ncS��S�=��|������v����NJ D�cgg���B�h�� ����Q:EQK��F�&a�v[��ܜ�sA�T���Z)ᇰ�?M��}sx�X���,E���S7��{�q��Z.�&a%Ձ++��'+��K�("��H�ڱ��ܞhrjԖT��d��%�!��ض�[x:Ù�n8?^~+��[30at7�C�>'�-d�C��� %A�5��猹N;;�0B.1�yI4bam_s�?�+R$Bv�� 4CIZ�^�j��R#��~��M���쓑ȃA �A���-+ {#*y���9Z��F�D�;\�^��5c?�	9���	,�^�c����e���B�*E���"ȏ���qkV�}�ekt������sɱ!�ç�d��5�;�9X%[G��Q&��9��Z� �j���1kk��}����BJOQ>���A.n��1�O( "q���h`����D��|t�V�d3���4�%���c�_$K'm�|�0\(��~�=V��IVJa�������z���FB;\���x߹�B� �x����^5X�N��`�����w"�h�T._��V���.�vH��� �s�r3+��>=?-d�� ]R��7d�^������?�s��&F���װ`5�PѲ�����Lx����v�
�8e\I&�j�[E�Od�����]^����I|Hv�a�Y�'R�$^#'��=�RO�Qe����Y
�p�.�!�.�w Losz%���[S?�B�/�do��_�@������c��O�������$���0	S4����s�RA�Y�\k��맬]����v�:�
ύ��í>��|��#�Q��qa]��(Ϸ�!UG�I�i{vB.a[}�m�+�_
È�V�'�p���^�@c�Ӈ��	b�t�i��������TUa�C��I��H!.�}8�#Ә<��!�z�J��<Zѭ�ݲ;Z��(�^����!p�(T�Ɋ惪~��{w���n�<�����j0%\���.��:y.�](�$����s6���@�կ�⇖�Ex�R(�Y�Cr�8�c����w.�݈GE�]h�`���S�m��jP��P�(%��ԚO�Q��®�Nw�5��rMj�	^�$T�c���7�]�_��Y{��N��^�&L�pT�g��#+�"�����:��<��A$��4����8�*C��MG�q�~Ln �j�r�)tI�Xj��Ƭڦ��a԰�ntIs��$��u����S�9.Y�x�#)yH��iP�7�]���4�>�=��\ۯ��3��y���(�G�;���←cF{ـ4]Y	ROP>��n�����4(��e��D�G�E���P3LJ�a?e3L�5���<�7�fڊOdP�jF0z�I�Լ!7ü�@�0����͇��@��wq��n�_��~�ys���	͐g���&��O�/�f�RA~U���y1�]�0��t3V@G4vĕ��Od�M�'�j�p��7�;s��H�H��G�}Exl�]Ő����Ul>7�RɭӴ� Nʾ��Gj�2�)(�]�I����;�B�`�ABs���w�{2�D��5r�aa�	gw��z�\����M�#�Al�,ME�]Z���I��>�S�����b���_��;?w�����h*�W41�nTR�}f��|;���ެ຀�n�C<7��
h��hy����h��T�! n��A��M�����`��>�������)Y�����wRv*Ƕ
�pż%�n�M7�ė�i�V�0B���
o�r�r.:����E�Q��UbY�\J���m�~�n�����d,h ����J���+��O�,��(8�ҫ�>U�F'@��#9���͏�,��W�mR���C���h+l���<'L�E�U}��RL��I��U�y� B�E��%����zl��+�*~��G����U�L< �5���_���;'֜L:
 `�D���HR�yF-�S8�Y��~�QK�R}����yϴq	*M=Źd/D-0��1��)Bj_�I��$�?t�{��?|�>-!�6�O�O=+���~�k�5]�n�D���ʟ!AO���c�.j����v ,��G�s�}D�Ο���<x7�];��.T����f5z�q�HGMw��\����Nr���2�P�<�tB����.9��h+h��Zr�e]it9�~(�=7K���ZW�D�'��4��x
#�7_Οp����p�N�W>5Vɥc�Mj�hxN8���>�t�vZt������/��"w�ٛkq��ٺp�/=L߸��r�~��2lo�*�tØ5