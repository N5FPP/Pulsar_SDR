��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ;l�Fv1�ϯq׆������s@���'����j����դ�P:�Cb�{�'�t�ɟ�>��(Hw-�u�� !i�^lZ��C�{��И���i�-|�|�I�Dd#����i��	�4�@$,d�������v=�3�A�pO�w�tE���M�ȼ{;��?4P:ٮ�7���F�ڦ� w0=L+=~�&P0q[��^�-\ߛw�T��e�z�"�[S��B=q��È��A7�D��]�!Tl�f�+K������<d��\�毙�����gpȷX[���;ފ@n�%%�WNr5��X�hqҶ�=PY�0��WΈ>��uX�+4 ʿ =�������5�i	��,�Hɴ���d��h�(P�pFtk_���'E.ݷ�T�q����l!�&˃S*��, �FȽ�'(�k���=J�?�>:̃�7�\���9����Px%[�C��a�d�%�}�qyh�!�ۍG��x�58��Θ�|l�zFSg�\j=)霃��f��L�U��!�@C(����U>�RRrT� ���X(�A�G���I?�/�I��"�?�Z��E�T�w>�3p�>����G�FJ`Eޑ^��&z9P4��,�N���*�
;�˰d~4�� ��'�L�͛�e��ث
|%��QLZ��s����9[S��ʝ��:W�7��������gG�^:�6���3=x;-��;
�
��_a���-�V�,+Z���N�69"|����a��tZ>�G�.�/�2�7]�Mg�S@~_m����7�ZҫӁ(�,�	2?���G\�^�����c,Sʴ� ���F�g�\OA6��-+���L�����**l�K��:H�\��B��r�A8��ѵ��1M jp��x���?S��p�k��ʷ8ώsr>!w�2�O���q'y,�g{"�b���ipD�L���#2d��!��K��VFha��_�
]{P���(���*8����N}��^�g����~�I��!��]RҞ��ŉ2�$���S&{=�2�*�tˠ����ě��Z�l2^{�0dR�޹��q��uΥ֕%C�
�~�Y�6<�~���*3f��T�\B&�
���hp��Zr�*�u����TzO���~~��_�9��8�J{ܙ=�j2l��$im��F���?��c��	��L���؁���*6����L�ήR���H�4�����
m�����O��i���0-(��t0;�&��D5r��P�-$�`k�Q���hfk�TnႢ��f���u�[9Ȩ���c�<%��1�S,aUb�B���dړL82��$c]�長�4��iz�Z|˥�H���,�<�Q��"��U��]s>�1�n���oaR���gs�ZT������%&c?�I��9Fϊ8����E��\tw)T�l$���i�%(1qF�(��z6��%���u��?b��a�l��P�=
p��FY��&$���#o,ϣ6��Rl���$��,�*��~�|��͊P#5(�c�Ʀ�%�Grs;��1D$2�`���P ����E��pH�w[�� UҶ��F{���$û�L�@`e
�ڎ}�����k�2-���u�z��Y��V��h�"�G���N��Y�S�2�B"1�Y� eU�t�/<�h٠��r~�$�y���L bB��>�LR�J\ (۬�,��d.�)��A����5%��,�ʓ�]�j�eX�\�[��2(�[k��v�7�ݽ�$�'ѱ*��Pm�]U;ვ����I.�Ao�<��F����ŚW	z���[()ً3�-�F�K�N9�ͱ����6�}�+נ���/��4!�om?2q:�MA�+n�������L�-���:��0H��1�=���o��l�,�KE�;�M�m�Ȓ�3�]ɿ��&۲�f�&�E��W?g.���:h\�����iJ�en��A�9�� ��[��o)�0�.>oHO�� ��Df����j9�O������\��d�����)eg�kBl��z0*C�#�LPN��v���߆թ�uL��7���ck���;"k��5��x@P�;��Ux�aa�D�'lZ��<1� (�]h�ǭ��A��S�u#� ;��=z$����Q&kP�'�l�c�6`��W���@(,s3�.1��n�_�]"ayGo9$��opG�J���^��H[���R�G�f]�E�B!{�#�#��c/��F@AYy���z�K����]%"yG}�ҧ��|��¥�|����\K�9�<c�g�Y����`t^	�	ʲiD?Lm)B���(Ю;�;�yr@�{�^q���(�|X���h5�3&��R@�]9�n�W���#�
5��	H^Y��;���Y	C�V���W�0��}���-9�G)��s�e�p�0_=U]�	�>wV�vW�	p\��?5*�F4(x�²�Ү>6C�Q�W�O�o�hy�nj㿚�:I�Ĥz�6�:veǯ+�W(*���,���C��֢���h���!��`�X���x��ٻeo�\��V�_��t@��n��I{��[��OU�Y�A�z��+��Z���>Qz��	����Z�<?Ddɻ�Cx;�t
�6����ޔ�T;��R�J�Ь��T@���3��aNU�����nt���xb��55�,���@�q��8�r�Ċ������Q��_�M~��#3p��6��1���bF�P�^�>I9Qs�Y4�Q���}�Zl:�!�aӮ}�ƃ$�2k�Y��ˡ	���_\����vߓ��2W���Y�'}7TJ_Na{�N�l�4�׋�<��a&�.]�O���A�sA#ٓ�+��⏫;_���k�����1��1N�o��f�n=�:�����5�3 ������<N����7�VT�yg�?��"�D�T#ޑ��Z���9E�6�uHm�YY�X�2e�|X�q�u�&� )�ۣu�� V�I8|��Gc�!w@�EҪi9���N���Q$cE,��7]s�O�5ş�F�nTY�`����.i(�����F�3��t�c��6�x �6��)����8�����(_M���sOC-A��� B�4it�}Pc�q�Z�-+�2?]S��A8��Y˟���d0����E9􆡆�7�{�!�)/�ivuh7b��p4~'�E2D���z )
a�[d���_(�2g�//&q����3��+K��Ѭ5��͗4j�T2�F�/ֺ�s��\Wv4r^�}T0�L��] ��Q�-Ϳ�S��7�ǉ"ֳ���/��O���q�|9��(�2\�e a ���p�c�I"Fl�	�u�i1_�fBo�x���m��[�/۫8���P�=���`ݱҠ�~<��R)�2E�*	]@nm��JZ���{׹�շ�d~�$\.R�̻����k�Va�;���۰���8MU��ZH��&�o�%i�.d��`�<�c�6��|����a�&��c�A�L���FV�g�-r(ح �r�M�\2���C��XO6��k]* x�d�˰:�/x���������bw�$ �tϮlO���PA_�3�	��I����u�)�9�y�=*���]���#h�S�ζ3��mp���2Y\p,Z哤2�c�1olA��}Ar� �-��(��$ ����$��-��+Ct������H�J-D��c��%��=����c���=��њP���:�O;����eӾ8��~�<�I}��)��c9�	S�pʣ�T��b�-��
,���F<p�>��� �S ��"ǉ���ܚ_/o��.x�T�T����	!.|�ᢍ}�6Ĭ�����c}��@oo��L�x���c	�l�{x��I��g8�)�=��܇F+*Μ2�ؘ�Gw�;���>~d��1����
G𮣴EF'SmX�SKS�ԝsU!@�L�H�"�|�M�[5�{�(@z�y�}đ��-��U<mc�L��}�eJ�J�_
������%�w�@�Ѵ��m��vLR���]p���݈�q�ǈf��Ѧ��qvyy���I�A�Z0�����kTԀ�����,YOɜ���x%�rN# ��E�;���dg��K��	���$�,e��	��O[����Kt���;߽D�K�������;{�.�U�K���\q-���ˤ���reN@2x��쉇�`��R�M�Q�3`3\�}����=���M:Jd6��N�U�|i����\�f�Ȯ�����<�����˲^��7 ���})OK,��Y0`��'����d��1����lB�ϱ�592lձ���T
ݽP����a�[Rt�$�lY@9o�?�Pb��5��w�#zYw��NA�A
�'��b4�BfÏ�-l��7W'z��p��:�*����r>��0�U�iɇ�;� �B�=����?\?��e�νJi��B�ʖDG����֞I���Ȕ"��2�P ���2.7�̧�k���VS�+a$�t%�
Ƀ'o9�q�#�zk�U����L��5�e�Sތ4��xh�0F�cl��4	�/�M"����`�r�,���~}l�60�WK�\]�Rm�ho���-���Գ��P���7�����3��]��״�:2 � ���m%k�󫶥�/3I^�l�����G5��n�I�g1�����*�`����Z���t�TP���*�N.�jv�%U�y,gN��4�f.^EJT�ʚc�h�/]���EYܤ�R��ŚP$���G��ҵ۶W ��R����g{�z��M%08���&b����GI<(c���_t�|%Y���Ib1�VYa
���ȓi�_̀��>���^�L�7�5�;�����t1,3B�|.J���߀)�������w]���/����=����JDT�/�`n�5�۫��c�3;�I<Uaӈ��Ξ>��bE��;�)xe�GR�Ñ���G�4�IC,�������An��W��#��\��uG�DQ1�&�X�H��/a ��[ZTfk��_"�ɹ�~����^������m�8��Y�m[����ZЩGP�QP�e2L��f�=�ђ� �_󡓙�)G��O3�qks��&\�b�"	^�k�By�1��#wSs�A	}�/�ivL����6�gts�iu��u�3]�=�Q0K�	�i�*�4��߷m��o���X�<��,�Iy�+[�٦�hb��P�~�/�gͤe����#��P[�i���Kõ �Ǫ8ra�����Ou5HI\�=:��8ޜz�#�r{6�|-�����A�dm~��E�j�%��b��5E.ގNl��\�ja'	�U����e�<�x-�ɽZu��Zo����RnB�]%��s��e�Y�b\h�?��u�1��O.�@[T�+��3�����II&w].oxy�/���e��_��j&�l�	TИ����l>%S���ì�_ -(��ዒ28r,��/]E�b��'��ܛi�������3h����@Ӓ���y�����
��b�L������ܴ���ԍ���v�����O�5#��7�b/΅����Ѝ�Y��l��c��l���><}�ҕ{�n�u8�>�M��P�0�zi/!��)a���u��!���n�U�d߱��SH�,;�kݿ�>��Kfb�ԥ�d�[��@��2s�hJ��T�#��v�b]�ǏpH=�V��H�8�����>�S��'�baJ�pf1�����=b�q�3�'�˦P6���D��L��������I<�3�����h�ʇ�`*b>�nv��cgʍtح��aVJ9@��mF��@�M�P����y[M�n�l�=˜g˸Wu3X�Ilϖ>4�v�g��n�$��-&lQ�Fi7��|�80�����_h:�Z�s�c���t/��b( �cc�2���&©�D���.�d��e3V�
���mw�p^���R��Ĉ$�N;Z�%�k�D�m�܁؋�eKW��ҾhN��4���'Y�I�b���<J����p���@�
�Ⱦ����w
�V����������C�ˉl/6���g%�!<�:�� 7��x�Q'%���U�0�j�v�nb�yi�1
I�b8��~�y��߽9�=��y��G��%A$s���6��S�o�h������*1䮂{�]m6 ��$�I�pOeV�}�E@
t�������F��p�;�m�H�o�],� ȼJ=C*��Kc��ql�i�|�ia�#���IA*�u�EH�N�2�~s���w����9��dO�W����p�!��dI���l-�R ���]�
6}bB�1-.#ƾ��iTw�ܝ"(�&��*�߄V���&���ꎦ�����2�Ҭ_=��p.�;��yq@��>/-`��s�ڼyn`��*P�C��T�f�������#�!�ِ�8��f�z��K��$���:��py��n�Cy
>�&$=��ƌ��)�jYb>.�:{�鹃 ��J�ç �4sQy3��t���`�����!�R�WI }�j��7,�x�5��Ya! �V2�:��9)&��"am���?��N�ϗ�Jz7n�;�Î{Hd,�>4f��	��+�P2��\D�.�$Tȕ�d!�Oq�n��!W@0ȧ�I���c�-( 'ncd9��Ts%�[
x�@b)w��sH�Y�>��8!�P��%`��C�����O���<��X2%�O/u�ه)�.�`�����dM�
t�#a����@~����4��ĉdz'�4�>B�rC(I�@h`- ��Y�=��i�p�ȩ�RH7o�[)9&b��q\��kD}������H:U\H1��_+�	�{�-R���k5�C�"���F�T@�����Z��{��
�+dH��n̡n�<
ЯT�4Z�F����\8�.�Vn�3���9ULR' P%$!?`�Ai��SL����X
�%EPL������l&<����[���f}=���o|���)�[���~W}3����@I��\���Tp�WA��м�j�C�,w��Wp��}�}�c0���8���������R
M����c�JzB��j*�]Ja��9>����7NrH�@M��U�j�C��*2u�3K���Xc�� *.z@�C��ܳ���p�*�rc�۰��T���omc�V�m��m�d�O4�F�"I��떃�8j
��O(w���'�I-�Y�D��J��JM�5����ò�����P���4���R����t���KY'@�
����`.�d��t�_��V)w�غ��	֝��p���Pc�Y�e}������>k6m�/N�,�^�����2V�Ap9	d(�����];U��9$H%D
����g��;q�>�E����'^�9ϕ�O�M-�_j��x�����zH�QA��ɼۈ�a3����c���U�)shÇ��䡲�'i��T'�k��5�3�z?�:�
G������d��s�6��S���u��)��t��M-����ʹդJ��f������Q�kj�~�����袦-�l=1«�|+�B���v���izĮ֦�+mω��捸A`2t�4�͒�jU�i
.	�I���Jq�	���pV�t&���f� 0�jC���	_��y�hx�"}3�	�I�r
��6T� ��A׽"�<���wc�?��X�:[S2��7�u{A U�#O�\{����<S**na\����2��N�"�/����&!��7���� ��zr�������-������n�%�`�I�hà��{�^K ��S�WBRp|����`�J��U�W³��U�m<\�Ai�tF�>���#�>o�Y@����L��:�'�ŧ-�}ڢ��V��חS��9�D�~�Y�4�{z1���R���I"������_�^��jX���=}��B_��&" �'g$�H����ܿ�X�v(ӡ��$���&�R����3=2�x���ҍv��M[��I�c�Ŝs�}"؃'�ӣ�(�Y�i�1ﭹ�m�a�&�P��QkZ*�7��9:HP�zQ隙��L��@X�)�� �NQ�"U^�ͯ ��Aw8�
�"2!@�<�.M ��7�rN��k�'�n(��)��~�n��v>MQݍ��K4'�P:�-��00���"B���l8>�&F�е���& ûEp<׳�Ioڀ;�._���h�!���:O���՞��J�2յ2�r���P��~Z�?��4����5+�m&���<��=�}�1�!յ�w����o�s� A3=s���+3%K��0�֖��*/r�	Ջ�7�j߫k�J����`��"i#u`��BM���Z7i����)G Ⱥ��X�/G� !yB@h �
����A1-�ĠFwq�[ �>$���݂���5�j���HB�U�'����d
9x6?�b(�ìs��+�~�~؄+uQbU��w�a���Ph���L�\E^���#�d�_�gm������:���ƣ׏.������z'x3���io��O�.���ZTП�i.��ڇK��j�Ff
x��O�����������{,c�Ѣ:�k��a$�%#^�~��_�JŹ�����ϟ dDa�9��JC�$���"�іõR� �H�00�DU��I|�4h�Gfُ�q>$���9�#1*�F��"�>#.	��b��1�"/F����k]F՝�A���xR["U ?|��	sB��F�����+{ğ8B8�o�����i��T8�v���o���<�D����X�K�x3��T�J5_�|��	3�y�#��'��?�R��G��2����Ze�q���L������-W�$tE��k���mn���T��k���!�T<;r�r^h) �B�l{X|ى:e���X�h�O�j��K��,��~x2�2����7ϣg���Ш�1'ڍ�����*�c#8Xɮ���u���N]g�4�s��e�q�Dy@�n�gIC�Α.Ɩr�͘�5� 锻��0��/�W�i���p�W�P1<�Ln�K	n��6��9�b@��Kܰ�D��ȓ���D��{�+�O����b6���$��c�]�Y��B XwT銏zVЬXP6�� ����Y�=Y!�,��[k$h�E:a�Rj��t���(�[~���hV�L�?����*�����_x��6�8j������>6_����b�7��W|���m�z�eݞǊ���U����W#�؜g|��s(f�Â<�� Rx��a��3[d�#�$�l�)��ha>���'N�k4 �����'�	:$Eȣ��n}���ZУ݋
år�/R=	W�7�hiz`H.��4;>^��<���B��h�H�y;e�b����w�0��v1a�D����Ǿ��[%��0�_F�0��A(w.���x�F��#=籦Ub������
t�.������^jk=�����T�߭+Y:O��N���N̶	���њB�F/����)d�� �7�򀶟�R�C�,A~�'x=�!/�^�e�4���kudr���'dp��r����°�I�F"U3>���"b�b���c�ɩY�����"��`��^\.��R����]+��B_��!��uM���ҿ1��eG�r�i�@���K8�0m�P��5��B3����;��&6#9i�ܼm(����]S�w6�
�| 3��D:~��	
���|[���⇮��f4�*�p��Q��<�
0�z*~�TC�z
k��!��:W�����"������D�t�)j��]��]֊X����-��@��D�2&�N��&\�%�`.}jc��S�t�Y^
�`���5���|�%s2�u"2��=��7�~�X}K���;t)�ܕ�tjY��?Rm-ŀ[J<�ɐ�B~���oͺ�<;ū���IqN��7�G�j�������4ɯ�gǩQg���-�l�-A���D�V�}Dy��Ũ�q���
��Xy0�_U�ʎO�C�Q /�&�@���Nq�{�Zv���@�U�k���t��س�w	{@L
~U<�&�$V#C�ɂ�����S E@�����po,��s���ķ���o^ܧ��]��/�=�PW)6����C�W-����(I#Z�Rm��'0=?<�A����B�c!���&M{���!.븭	3�@���4C�x��[��lݴ%��+4��o�@|��#�2Y���u���!Qy���]�}����d��+����#�����L�(Im��"�"���ࣅH�>j_��;�ә�B�~�3�1z��Wj�N Ɇ��p0'x�}��Ra�F�u��Y����߯��`�o=A$M�3B�+��+���'�g�{z�Q���2�4y�}>v���48-VG������m�/J��0��U��xa