��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|n�\&�����[hc�>Z3�S4���"KP�$��h�I���@�O��m�SP��Y`Sڲ�G�����'}�f�n��Jf{�k/I_8�~5b�(����q�OyC]���w&���{���t�Tג��wr��[٠_Z�m�Q�p*K��-�VQ�)
�
tv�ʊIF��(��D��,s��g":jn0ȃ.:0"E�p����<""=OA8�vWp��l������0�8�����b_��p�r�g��h�}��=�d����U3�֛��;yO�QA�����m|U��T%�s�I�hb�#�ق|���uu�sD�Rz�Lc�fI��n��s��(^9���Dp���a�
0�2��WS�/���l�*��L"�����L��EE�b��ł��w��H����V;bﾕl�����h�bsʕbH ����?��F9.��V8����-�*{�@��s8t]l�X��7\=������$��r���k��`��ل����Q��{�ءp�u"א�s|e�RtY�%Z�zc�k�� H��c���U	s]���-T�F����w�������<�?�h����tWJ�b+N!7a�6��L��ﾰ��C�3;��4��K����oKN���FZe|��xkͨw���Ψ�v�h_sM���C�f�ő�Xv[�G�cSl^->f�k���@ܢF���ʧpS!w�~<�`�=JZ���w1�@]lvk�� �'X���N�|4�-B�$����<��c�VB�|/�\�Zzl�sJ�%��&~Ŵ�E�e�Z�e�y׾hY����#6ݩvoy��|EwW	�Ű��ƺT�S8aOC9�'�������t7n��0�o�,���2+�T��˸UX�#8�E�eX���0��"��L���6�g���T�ѽ��� b�(��m�tp�(
}wԐI�S���UTV�-�V_�=X��O؟hs;� �
�>�3H��ٻuv��˷�����$ �_�:�dZu��e�m��l�/��nԆML�v�'!� V��b��:܃/!��,3U�+��#������Ȯ!!)�u���4m�������A �Ԥ��0�!�p�4���NF���"��q����L.=p )+>��������a^~��Po�-��m�m���O�
Dx��ok�C���{�y]|��Y ��E��u^��w~���p���Ty`�wE��}%�, ���pE��őS���c�6P�0�d{6�~�Jkz@T���j�gi����5#���¾���o����a6��	�~��b���#���u6����zH�+�Ҫ�-Pk#u��7B��T{*6�#��9��ɦ3RPI�Ƶv	)��{��yc*/� ��Y_�Z�v0��+��h3��#�rrV��J���O����F[r��FH9�l�+;:C5��lqf�k	��bJ� ��[jG9;�伲L@l���]/��O{�����*�w�5��=���['v�3#>�c
o�ǘT�� ����s	���BQ��l�:?BYt�ӗ��7I�3ѯj���m�m���YB���
�R-���DߺR���7	N�с��!,kuy�u�y|bƷY?j�������O@�@i���O���GM&����2�K�@]6��X{���h�9f��M�{���1pN�NVi�?��������G�fK���3)H�nIy��p��$�C*���$o\d$�~E��j!F	�ɐ�z����v%ѓ��,�;~Π���_Qi�J��9��f��eܭ+xe�Է%�Tw�%�.j��b������Gd"lf7�#T�����P]AP���J�?o�AȖ�>��M7B �
0��Y�W��g�q�b-�^���X���m����9�5t7�,��e�T;�.���:�ER�yp��{p_�"yF������½	m��"��O��W�\e���̻L�1�pɻ�����F�׵%8��6,Eݢ�U�g<�.u�Ǡ�$cGٵf�R�@����j1���?�(���Mh?eQl�s�ړW��2�C�9�.���f���HJP���P�`_K[*a̢D�����S��0`�I�N�D1��k�a'�t�9ݢ^g�I=H'*��4�r�"sՃ����L�I���w�/{�904�=R��C�!�/�����B�~���p@�nlEÓ�+��5R0s�U߯M��$�h@�l��u�I=���FR�x��+�9�<8��]-�a�I!m����%�Iz���b /
��Q �V����=�T4��,Gppi�݅Ͷb�	�bՈ��9�-���5cN��K滶�
g�A�U�^����=�Q�ޗ��!Y��v	W�O�5�[L�Q��ˊ�I�g����q%<��cЍtwՙm�ww����܂=���#����>s]��cя� -���ʙ�
�I�7Iŷg�������ҡ�Ԉ��Aɩ�����]�Z/G�Z��1�^�i�C�UX��U�\=����q<(���(B�H}�Uh�#�������o���HQ#�!�(��8(w�>�q}^���ȇ��4�(5�f4|Zq<��S�m��f@�SJ9����"d!�u3?�iE�uk�`<�h�`�e�cC&G��uUJ<��l�@Q�/b+Up��Y�ԛ�YX����e�ҀQ�ɝ8� WZ��Loߩ���L~I»�Ȣ���~�IZu������tq��ctbM9��?E�ܢ�&��GU�+��C-Ό\���������w�i��X���x��I��pIC�qݗG�H~4�#4"�R�&�z4?J��Ǯ"9�ݩ
���o�cb���>�7?��rXP!�u';m�˓lLZY�����7D�|VR)���_��D>J�����Jp�������m싼�RC��P��,����uS���I�q��]���IڏsQ-�Z���q]�\�K�c��·� ��o����=o�+e4�G0�ӭᴈ�<��[��w�Z���*4`j�bEZ�I�����M�N�,�8��'��u��QM�(�~�m�A閂5��l��j���8�V.K��uDk'����c;G��| ^cupZ7���_.�5�)nڀ׺-�8�e�qQ��ծ����#�(����9)Kz(��D!��B�~�$��=sf6���Ev�J��曯�v�5��o��rµ�z`P��F�"�K�Ηr�R�-�&�4��P$����c�l����{S^�<D�%��+A4�[5Qm[Πӯ)�.�A�'��df�nn���u+#W�i7���g�X#��]|�����T6%��*V����:Ƙ"�v��}���y�\���%a ��XޫS�M�S%��_1��!פZ�E)����u�u�ū�of((���?=�+:�f�����A,���'%sQ�����z�D$j��;m���7A�AN��'L�EB���,����g�ǌ���x��V����c+d�YS�v�*�����c�%���DF<�f�Qr��hN|(��_��� ɛ�%?^�:��W���:Sv<�b%:i�P�(pN`D<0'����#���s1L�ђb��^(o��qi�~)i2����?�<h�4��f;�WQ��,���7���������6�P/����Ճ���0�4_qԕq������ub�m�	���x϶�|���՝���'EzH�)��3!�:e���O��mJ[�8�ԅ~ɭ�_�c�G����8� �
��Qn�hy6��cδ����.s��Xb��Q�������)��$����n���-	P{.(��,�xV��FMjn��Y�۠�wZ]��
�xW�ַ�0^h.� �kr��R<�Ada�J;
V�uD1 R^U��%�}d�S����A7�x]s������a�1_G��U��2�Ǵ���,��~#���ƥ�9ᑩp��
�Cll�NK3�*o7*;����)�e�߁ifB��Q'��|�[�n���=�q�5�i���~ؓ�n�E��\8��3�������o.⸆Ԁ�z�^1�|b�����Fki$�9�&����h���y��~eCGr��Ÿw
E��
v5��'r_���#U�	�Š�І��Cz�)�	}QE��x���h�����N[�#�=�z�U|_͢�m���(	T�ȏ$�����k��2�-.�;ڄS/һnN���f]��$�%��j����q�i[�QH�w/�ֻ�|��ܤ�}�r[ɇ0N��3&�a4���;:�Q�z��MEݩݮ�nq���%Z���F�����7��B�AdrS+OtՉH���:��!�j�-�oD����=�C~��A����{>�*G���&>.��%�QP�(Q!��f���",u���K��
x���-�Y�eG��v}5��V�����W�)���O-��Ѭ�K��B\�g��|����S��
'��H	�K�ڹ��d2����F���LJ���v���|�/��(��O��oCO�1���%�+�^�>�m����V�MQH��^U���%D�3��C~�Yx�vh�V6�+ԩ�1�Lo�0+�r�3:��iٹc�oz��k��P�p�L@;���t���i�%�ɐ��IWқ��Z��"��S]�f�2�oK4 ŧ�� *��܃�ر5Od�!���D�����e%W~rN�[�9��DF�ﷷ$1�S��MJ�g�1�Hm?����M���Rc�\�~\��ty��� k^�Z�ͩ�N�S��iC�M�}/�\�[�_o��d��C�S��6	��O�H��!��J� �yl}�y��0�l����?F�d�D(&']7J)c<O|�2$s�>u�hA����r��a���E{���4��J��LґLz���I/Q�B~�3/(�ֆ�[S�y�IB�A�gz�vu�yR��xX�u� �Ez*�<ףYSBz�A��pO�G���8���MzB���h��<�� �>W�+Z[�o��ĸ�n��g��Zz��s�,��	���'ة�($ʊ7��K�|�o��
{]�˘W���s��# ��l��[]�l��70S��
r6�x�2�Rb�V��2����kJWP�=l&�n�I/>�x�6i�!T�O��9�`�i�  @�G��«�jM�ي>�B�Nc8)+�S������Sw\K� �
hy0���؁蕙���x�%o�3�U83���l3�vQ�Xb��q|�<��;��l'�ՙ��B@���ܯ�H��ׅ�\�bΤ&�b��o���e?^�(�T5�e%K�?Hu���{9���8g'�=4�W��O������#���U���m?�CLpt?6�St;mC^�?�b������0^�CQ�*q��B���|3v������o��-D�]�� �:�B��9�����mF���1㑀q��i?�`�>�4b�I3E�
k�������4o�E�|�e������1r ��<|��1�R0�P��B�4�A���G����f]QF���?	�Ƿ�>,�#�u�ʏ�\�d�^��:��W#����}=�q=���T}�JP�3u=��FCI ^�X:V�l��P�y�jl�n�b�<7�̺<��FV��C��@�~8�0����r��6Q����y�`j`��n�]�p]�G��eX���B�>?�9���s�!���d��E(���L@((ɐM��'�q*����kBf�e�G_���:�oDy{��J��b����~3�8�p^3��ܭY�>E�df�Tt�v�4�ai;��os��q.1{U�S���v&�M,���.�J���N�Z(D�I-m,��!�Sk������Ob����U�>%1��BE%i4��_���9X�}���	^6i�t�����ŞC5�h�x��~My*x�r#����E:"d��M�iu�@�]�ΫW��\��;��cZ�d��i�����S`��D��m�u��V�ld����N�kn�5��<2Z�Frk�$aŰ��۲#�q�+�Y�S��}�k�=�;ը|�ę	�;ۄ��m���%ȇm�#�WJ/�7 ���x&(���,������jlҦOp�f�]��W<,��%�+���к�&�X�7��~:�NYhԸޘ1u����:\�YA�xb�������8�U�o��(�\j�!UY;c����:�NmQT�K'�	}\.
��p��&/t��4<?�������e��"*�������\���x�ʢ�H}iA�%%���\�����,/X
"��J��c����|on����۪�.�6M�Tp�D\�0<�1W�~k� �)��%�X���3�b�Į�D�2�C�c�n����u8_�sV��E����V��Hl	r��I��R�H+��I�j-u���F+��"E@�c�����:�6x��)E�_1�C�K��;y2E�M��x �̷�8�y�è��g��M�j0��}S�D��%���$��7*�%8a_o�BQ�#s�Z
�(�����i&�b/`�'�cg��N�N5N̂M9��_�Ě�_��a�a�v���&*�D�eqrfV��eKJr���4{�C}6Ә���l��%Jχ!�䓾�ډ��94�'X3	V���|���_��F�� �����xÍVo�#0���O>2b@ѷ8S�>������0Z�ӈT1�Q�Ь�"�m<�7����L*2�^�"s��ݵ�3�ӽ�F���(�	��k��P���M�m��� 9}C0�S�t������B�۞�U2�N�[�������b<��P qO!ܲ�4B;@<K��|�=hB�$��l�$�G]���jo36����r�<�S��Efq�1�ǚɣ����d�fj�`��<i1e�Ė&�2�-�F,b	.�{)�ֳBMl����7�E�!�C���;Nh䚒�o=���X,��zmf���y.�X/}��.+����[��I
1q�~Um6��Xt�Ld���ARu�W�خ��/�m "��5�R��V�q̢̹�h���/6�x�AS�D�[�Z�UQ����)�EM���U���5�O�������,�7�-�J�|v�T�tp�������I���4����R�!�T�!��{aA��JW s�6!֔C]��I,����~�c=���6.}��J,�s�*��Y"�O��:� ��G�f��B��:�	{�HTv�=�C�
�v�8�9�][�;A��7%x�YSM�R+
[��2��b��u�s���OQ?�(ݸJj�}��3'�B���g54mR�Ӵ���8* ����Hhw�C ���d��F�������A���������=�4}�H��#�����]G	�g'�q�{�T�>��>5ǃ]�DE 5gb2j5��u��FKl��(*�$����[�Ao|}@A`��,-�"9� uvv�������\D?�t�����+�m(�t�����5Ebe��V-�5_�)J���`�(:�h$X
a)a��u�a$��U@0��7~c;�%'�Q�`]Vv9N����"D��`̳���f��<=[���j���^�x-6h��c�:�q��2��S����F�
�7�A�U}�2��U�Bҵ��NL}X�U�����8�>��"�ՐqX��;�mÂS��L�B^;�9�Ii������n�q_��t[�a�����;��*H�O�x��r�	��.�dee@��������B$�M�-h)>�.�;kB��	�y��љ�oF�M)B�5�Kr��2I>�e(�����dՙy>t���U�g��� Lon����	�y2e�n�����>@z�I�J��>=:��C8���(뷭:��<���kB)O�Rؙ��j�m��T�u^���ԑ���>,붋���t
겧 d
�}���@��v�����Y�C���'�q}���q�>A�������z�r���H��`�P�k�����X��8<�@��!��ŰK����{��iƷKC-��u)��3<�,�lK�"�"lkh�����G�?5�{�:+?o�ُ��هU	{���_^���jT�t�G�z�u�a��RBM+���	g����N�e�F#5_(�Su�Dc� ����0㜴�^=r���2<���)g�.�sF�7��+@8��< �$��
&f��b�Zب㊗E爛Fh�TJ07菈��j��G''���]����a������ �抐7�A�c$$SG�
o\�cM�o���E�N.���;2
y���mq��Jl(�tj%�\�j���)��������Վ% DP�`ݧ��@H�Q��QC�)TG:���1s�!&��?'P�q���ě����8��j*�1I��n���RϏ�b�U�����?$r-�^X�T��O��K�	gv�(��Ұy�w��EW���tڙx���3b����7%�i��Rd7�:�+��6JNѡ푍jш=�t���X]*�h-T�U�y��SW�c?&����@x�3/&J"#�N�6�k,�7O.��ၷ%�vJ
�߾����~d���b%px��T?9|����#�bk1�l�36����T�Qt�N��S�)?��YvG0�4�"��f6G�&Vx���،�a����v��E�W�{�y"�oc��mr��L�L��z�!Y��u�t�e������j�e��\fST}��4����&��߳V�u@oB��pP�L�`�C�U�)��kX4�U���RdMER�b+��%���l��^���9j��1��U���h�gL2���!V
{����HL���<V��&\E�bu��2���^!����AL� �tg����U�%w+��ȳC�{#]��7
d8JY�{����mʋ@N)��o���gS����\k"��*0�Z��\ƺ�Ø6Ps�n�ׇ^ebu#��n�j����EQ�z��RQ2�eW�~>a���Ƚ�9�\� ^^�N��	���cg/���Pg%�5_��Q&r���*"]����`�Mi�<fx 2�D��:	�|LǋA��<9Lۑ`&|�>�1̺_������<Tv��hӓ��ɟDc���tfDXk]��M��'2���."���D� ��$'T{�Ll��7D,�>h���Oo'D��*c�J�����N-u��G+QD������x]3�� �|pf�O0�
q'�<Yy<����;����Jf����%��a�D��B?����}ۂ@*+|��㾈/o�K��K��
�'��>hj���'�٥�8%�.��(��%3oЪ�ۿ�)L|x�|�Z�WN�D�Á�S�#)1�-����`����c"�Q�Eb|-?8��V��۟}����0r��B��āy�DU&�1��Z������F��t��_Q���+���a��}_0�Z΀��(��v���0��gJa�;�K��<�R�������k�(�������x|���j d��;x0((�dA��m,����(����{�1䰙�F�_���a�A��y�N{T��iY�FQ�a��]=e�D��I�2�_�КDv�wX��MC�^p&L��6P��g�[�HD�d�����Ģ�O?T�^�g��I֑�FѶ�4�������@�8��ƻ��� ӓL�b�U�����%�vQ�EG���WXE@�R��FE8�b���G�[|��|�-@˴rs���^+L����d�o��}��+S
/�j����ͼz�<�6��"��Әɗ7gy���Q#��ov%�ӧ��W;p�4����7\�y+D�2~=�UY��4�]�����o�i�}k��G��S�	N�w*K�K����f|
��Q#�`��h�O�?3�����K����a+?B����톎��3�����'.�<�?��nH%YV/7�(�P�%'
�2 �F^Ntl�|���h�@Tn�,~����������L�f�6s�b/�M�p%x�''@��wm�=���nr��q�KW���N^��^s�j��esQ���±�G�ڜ"�G��{���v��G�8:/��x��[m����DλDʡ������Z9Q�톜k�iڧ�Rz򘢗=�s�%Q�ɑ祉�	#��DBp�?f�4�ۼ��&���^E�n/�ʟ��
]��S0B�J�唽�b	� �c���AD�ۙ�#l���vM"<c0�>��T��"�(�9��$HW�!�C�l2m��7���Gd"g��F�Ꞗd�#��,�z���v�ɥC�EnM�C��x�8&�Gt|����q�l�tA'����Pg��V�J(Ѷ/� '��%���hH���O�y�����%)�a����<R�Ζ�RT���Lyg���k����! ����־b.0>.�ܱфr]�,���O1��Ս��{��7S�%���4��<������>5t25Vp��z��郉ԋF
k�m�:�ω,ƈ�%ϐ2�j'G��D����a��đ�4f)�d��x�2�'��"Gg�����Wl,���%SN����-E6�?��fs0���K_��L����I�3}��Qp1g\>o	���Y���=�%8`�ψ2��Fĵ�^lyJA�*���jp2�5��.���&H$�3Щ��I��5�x���~�}��|�� i��ɘ��u�M�7rR�6��k����MO�iI��nK2
.>��	O�_���,�-YX-��B;z~X�[�Ʉ[���=,|��A8ɯKmƣ��EZ��o��\`��`��Ͷ���Z�O=�k�~#�:�E�M��pgV/�/c�qFA�4�I�@t�r�O�'~���`r����px�\�i��^�[���G�C\�G�r��ɢ���nIveв����Z5���m��e#�%���-��ދ��bpN�>9	��Jc7�\��s����0�&�F����_�~�6�؝X��v�0I�F�����ک�I,R9s���Ip��n��������LrU����eQGf[������gd!�c�/�ϯ,�J�6�}��1ݘ����-^A��}e�eW@8VqWίL�O�ՠ��~���	�on�s`�4q35ޱ���	��8�7P�A�I(��F��\&C�[��w�����\l������T�_�)�W�S�~���8F��;���{Ьp`��-".i���<;�.y�P�Ƿn1u�u��ѯ��PD=7�>2���46�&����-[�-�9T,}���>�RE�<J��r�r�f�\��Iyg���F�pN�w�Wz�|B?�Y��=�Ȭ��<��<�W����.k�\��z��f�1�:��l�k��?�>����K�.��Z��K_��z�t��&D�-Q��C��A�tq/��!
A���#��RxV�A�<9Z��H�?��DL��^(ZS�g�nۆ�9�J�%�ʘ�ij_���kR,��IR�*���R��R6%cw*W�}!o�j's_˟�i���p�{Lwq	
|J���[Q&�Z$��ظGC-fV z$�nƆ]ᔣ,l�F=}���c�듌�F��}E�mpnmӀ]�NĐ�H��CJ_!���Z�"��<q��[�YZ}��E#��"��]���t����X	+<:j�A �2�@��x���M4|�
���o��![z^�(��U��ى�+�1�cy-%�;�b�����:#���(D)
�h�a�Cj9���(�Zt�Z��ǘ�p>��$�^p�����A���Z*�\u״b.Q�I^� ��Lɠ���OO�p.Ghtc�f;����]S����e,��L<�Z�<YpD��*_�C�@&�!��R{�?���%�j���X4�;�bU'z6ba!���w���P��oiC���v.�5��~��Ϫq'�x�����B���Wm�>{G�-��@)RB�a��y��&�*����*�E�m#�O�Ǫ��O�_?#���1Q� 1g��ݔ�mn�KE �q9��lO���*$�h��=�$�u1~�N�梊O��VI켆�k%�,Y=I��v���z��B�
+[�`�ӓs�ثVu%�*y����i�ۚ�|���{��7�4h��	#��x���/]H�	A���IA(��y�e��߱��ڳ]:�|�9���lԻ�$m�)�S;���I�%��u!����Zxm�<�Y8�$w3!+�k\ۓ��I��c���e}��^s'�D.���=�a�[��g ���uKlWv�O�態˳�"%��=Y͆b�nKX�>�~5�EH�Ƚ�@���7$��6���T۫��Z� �k9�}�C�P?���xp���(O�F��-�ហ��,f"�_8F�<��!�1	a��s�J:o��+P�����!N���/\Y0ξ?��@P�� �f����U�ן��.\��e��
��=�l�GO�m�'~��㿐��*I8~3o+8�&��O���O�P��~4k�c� ��]e����a^}��a���Du�������"�#��DJ⛰lD$��P�"��s8�Zk��h=�4���k��~� \mnjO#��\�/�D�
���I����.�%|`L��k��R����3Xht^�el�x*����B�FA�SjLб�?�=o��ۉ�6e5���j���̫m�r�掣�b���څ}Fi9[! Z�>�dQ�i���X��y?Z&�|���Y�	�1�(��I��t�����+}�/��=��ڑ�8� ����fY8 	Q��8��ѧ�3��Tԡ��?V {b.� ��R7��|��Xh�o�w����'�⾽7q`@'�
���'0&0ڼ.���m �E��CW���ݎeg����Q��)ORvC�߂<�=���かI�삸�v�=�(��ulKN��e4��=�C��_�=D��6#@)��vHz�]����񲽤5X��η�gE��QZ��Y���ԇ �0a��ށ�{M_�:����>�$��0��B���߄�4�8 l��|lV�$��@<Ц��/���%׾��ء�6n-��r����[R�g�ኀ�g,D=�w������#��+S��	���K\U0�Uà�]:�:�/a�T�����gw1S�i ��R9�zr0_�|�A�wȚ�%��g�7[�|��H���3?*��H\UN/���"&es�]��.���ж�@�����t�xh���-�U��blE_���t�����s)Q��v�U1대�:���E9�F3�Z���lVoMޓi�)Jk7#;}�?�[8�������	���#gC�v���Ԑ�a���F�\~�-�k�����sQ���פ{*q`����{�J���2uĒ�2�zf������ NQ�y�(`����u[t�;�Z���Q,�4���KuC�n�ڑv_��c�.�v.mt���FX�K� �fg�s�1�㗖����ȼ���#I��׭��������V$g�ʂ`cvz>�H��.�1~�-c��4��F~�p�~KK��� Ec�-U"�J�Ԙ=�$��a��\�����{���t�#~CԴ���@�{L����(D����*�	��b�[ZO\Qz8X��Cv��w�7�bI�p_w����Q`��lƴ�p�d!T��$A�	�/�����F>3$�Be��VY�U�:��(+x�Α��7S�i�z9~>J����!��L�j�}�,���8��/���1����	��,�t���L0ucXdJ�+�~mt���&p�Yk��𶪳j푒�H��-j|q�pJ�c~]��}&DtN)��OѷEQ#Ei/��KG���^?.�t�xm��9D�`C�3{Q��+?#R��W���'f��,���	�Ό�
lX�ޘ��Xv��1#�[�n\�4*:?���
+3�s�o������a�3P�NЍ�����S�p�)�M۷��q �<���p��$j�������Zq!�
>�	4�3�0؅���:	��B�i�K��ϻ�Z`Tj�CY�P���v5��e��B����M��J�9
'�9h���0�3��K|��r6�uvu�!�¥��;����lL_��K4z���4���1Ζ�@[-��[��/��{�_2�'���m?�?���1m���B"�c�\$�uD�^_�aoeC��C������[K�I�r��s�]��uO�( '��CV;�I���>ރ�,$��dY��j���-
'ѣZ�?S�ɢ�#)����dϬ������:M����g@ʸ+��4UZ�CrV�Ԉ���p�����M��H�zȉ;����:���<�w���䫲ٜ���ɕ�j
��9`��	���kKF���q�8��.�����|b��@hI'�E2�X�T�_ÿ�����T2�{�p��_!��񀲂)K�0���l!-o "�p�np��!)�%~�u_�w�=v͹ڞD�����Pf@'m�.g�} h�n���QX�P@$H�8v7I��ݝ&��']�Ht8.U���eĺ�ҟ~�,f'����-Ж���*� ;���ml=�����w���L�(؞�T����ѯ���a�"lL{I�a�ؼ�U��EQ9r�3���� ��
��7�
�^��@�&*�m�2�Ћ�9�X+s
<�h��3�L٭EI�Q�/�?!ڢK��t.�̻��k�9�u�`�t��JTA0�/�z'G0�7�0�EL�Y�˘m�b��/Ïp��5-J���$�X<���4fIL�F��Rw������<�T��V�f"iأ �!�}��M ��Eľ�ɝO�8��Z�F�r<p�4��%�0Q-[�-��<��O�v&-Y>}�A����V� ��f?���[��{6y�b�vL(3Tx)��Xbb:��4��z凮�`Lpȋ��5mt�^+���6\&�3Qt���\��.~?��s�C�X�%�L�I?�2����!4���&&O�o@�(�~��z���K_J\�&��$q=��J���%hu�u ���{�I'��������ӧ���|��9j�qc����ū%Ym(�WV�}uiSB �6z����mB�2���Il'C����~<����_�b�#�	RF�gv��<ƹ�ʑ�n� q]Cأ��"��+�b��/���b������S�l���-6gU �o��1m��oU������3?3kerxB{f�`
Y~���