��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��V�^�Z�4���%�ڢ�kU�j2��.��n�{VoR�.���g��ɡ��80EFj��ƕѻ���vBͿA���CeŢH�y��?Gɻ�+��aFqB��X�ذX����D6�y6�� ���Ȼ�o�+ܚ �'�J���ڜK�]?��p�
��Q��s�������K�/����MB?O^T����	�/lRf��L}�^��n��O��� ��UQ�%�e�r/��^u�gd(>���z�4��%�"�V��X��+�Q�RM��;��y��u�}�њ*����ʾY����ޫ�)@ ���Fÿg�Ee����#<ƥ�ui����K6�b�C�R8�f���N�����g����N7�ƚd��0�f~��M��ȿe��@6�_�4��� �#�I�1w;�f�Q�_�m<8�j�,�'�g�gX��v}���e���X��������=m�V_4�!�avKxApaj�Z�~�9���af�9��1��Q⍪�ih����G ��n��21�p��Htma� �򓋆P=fl�`�z��Ap�J�
��Y6!�B�����3�GF��~�͖�Π8:��S��K�U�����G��Z�+:�dc�]07�������`-pwF�l�:v=�}��̿CZ�Q��;���U���o:?O�<�*�����`��D�=�R��o�ZbRm�����.\Κ-=�+
�[
c��+f�/,�G��װNgEx�~�������J���é��Weڊ��^�<�`�����aI��{�h4v�]Uܺ��+�O��`�\0:�$���E]�'�����Wi�q����c�Z�N;�8��wd0*HB��糾�H&�/���~��Cp7*/�z��P>����U�\5.�b���6�ƽ��K񘇽o�w�V�+�cE�D�1���_�d/���I�u���{> ����H;���62�Eo��N��;��$�����~0�t�Y��ݮ��я����`	<6�u�e�qR��^�����-��Ѿ;>�4����7�~���o!�=�̓c�/DH$�z_<����}�@	�t.<3|NQ����X�\�W���o�~/���M@zu�m���%�n�ߩ^���A8��s:�B��k[s����,���j��A�e��d9��셆��؇��+�{�-��5���G} �B<�p�,~2�ޡ�س|����{����&3lp���������L�{@j�`����b%lO$ ��R�hG��Q���J|�*-�m��kd?z,�nwV BF���DT�oK����HT�tlބ�*ua��d)!�ƟV[gƧ�hMܕp��E�%l�q�7<S�-�"0u�3X�)�&џ�dq�o:��� S�P�0�bR6�%�l�ԭ�@J�nk�=Vo�P��v���`q�
E��NR�>�p�-��F�e�`����<��0QM(�<����(��h�W�Ԡ
��i ��=�Q���+M<#G ���}��C��]�ɈH�+�Z>��ړS�'��?7?"�2V��N�vk��-iO�n���DPo-B�C�S�ߏ�o�������Nk���M�Ӎ��	�AHp����]��9�< yaR�d`���r�k �n����l�9�ڥ-�o������H��X�Z�+�^��pt�
/��+�W*+�1dulP�!��bY���_�F�}���c�	�sp��.��u��x���H�M��:��?�]C���ɟ�^�P��k<��-'�ʥ�u���0V_͌��;P�n��.ӷ�ְ0>�^=�7F���f���������N��c�3}t�ғh�6a���g�����q�Y�l �H���-@�h�����?N%�Md��ܱ�A���6���J�t����?|"�qö��[n��N��-�$:L����4C�e�[�,d�y���	�G�3_��"&f$�6g���ڰKh'�Q�?n3)�	�}�H-��h˕kuE��|��R�͛��PXK���r�[ˇ�j�S���ܶ�lT>G�����`
��9U�(�lÓ'x殟B��L�!����x)�Qn23O���R�z��î��|�����YtM��ڑ8��fҲﾁ�� h��k�p�D	Z�w��8;�mђbG�m2��v�i��q�5�f�#c��#��Nq�̠�_��kO6��̐p����x��)Ě���.��YȈ6�Ú,��"Y�8�S;���QH��Q<L�qQ9`~_�$���[�[s6
	PB��&�l��N�bgw����
�ٕ�t�<y���@��m�WF
�.�?�#�0�F❣�ΑZ�˄�Y��}��:,�*�&tKJ��{kol��yNN'G�E�YD|5��Aa�W^��L��m%���"����֚U��wG�1tK�4h�h��C
��8��	tk��$4��Ä���h�Ly�@.��6�W���c`^9_
�w����P4N��wې��s��v/�8D���ͪ�'�g垚�"1��5��$��~��~���S�UI�p������4��~�y����=�b��l=���>~9^�mG�CZ6�|���̨`#�q���>������ٗmI$�؃����)��q}#�8#�C�s�P$z��jbK���9wi���1�Nu
����C� H���" �5���_���:ʽpv�s�|(J�s8/�����v �2z�<���W�Jz�II5�V&�4���VU�%�%7��/I��}l� �%q���s)\?٬���#�^t��؍X0���s���];�3��u�̩^��7�^����i8s�)C-���T|y��(�[�Υt>�I����Em��J(iK��Sb�i�Q��|��!���CPl]G��Ɇ���R��K�N�쩮*�a�+�垣~�h�1F��=�Py���uY6��Y2�Œ����D�:߿���y�}3�5�DT�-D�D&LW%ܗ%0f阊�\�}��1�>���,�IP�e$-���x�dŀ7�x�
[�ɂ�`�8���w��HKT�m��D4�%#����=��%��隌o�Nc��=��%d�Jȃ������z}@�?��gw�9H��L��=��h�v���/[�u���A ߑآ1��S;'p�Ve��H���(�^��P��x.Q�B�{)���^�Ԁ�������Zm.ɫr܋<��n�]�o�d9��g���ۚ*fى�V��N�8�H��|����Z��~w�����x#���`���� o>�22!�$�)V� ��x��jzŷ��g/�����7�xZH�o��%]S��U�� �kkk/l��q4 |�EvbJEW@��R����\?-����Z��R�hZ�UBMg<�rtilD,ۖ?��2B̖�<A58 �P���=��!����e�3���g�fG�3��&��R{�Ϗ�0ߊό,�*G?�E�����?�b�4ƁDȵ��rʒ|�E�L-��:�Ƶ`����n�����a b��d]y�����J��Der�MV۳
��A-f. |߬�y%�]��|�
$hL���<ξ If�C �$�{����ևK���Z���r�V ~p��|�W�W��6ֵ�)ڸž�9�c�AGƆ���y��N��i;�[R��(!c��h�(����0��]H��p=��İ'o�#�Ԟ�7_ݦ.�l1�Ǒ��8`a�e�m�{�u��o�G�%�\�E�MNq�/P�4�6��� ���D#S���:�q"�z����68VIJ� �z�;W�!j��	�u���FkEɓݣq�Z��[۲�ߞ%�u$�@!E)���g�N�x~�lGo/��[_S��U�����}����0��|G{�������I��K��&99��Q��Уo�<&Y��ˆSC#Z�/��xy���Z��fі'�F�R]=v��������:|#5�%�#�;8D3�Y)�/[ g�1� 0�j�ӈ,���_��'�������'�&Rb�kH7~��G1���A&��U@4��A����˙d�=g��m��/��&���9��N*/�$�m�X��m������B�X罍��zs�xpը�^|؀<��;��R�c|<'��.*�y�T=y��M<ՠK]��g:���k�g%o	����9�vF���߯15����8됦�0���I)�� ^~���q[_Rx��[�c��kOD;K�g4ڶ�#t�%�GZ�����H�h�;`�zf���l�Io?�N
B���ٷ��
}~9���)�=����}����o�5�g���j3�����ᶆ���Y3�&ux���x<��*H�1�����K��|#Uҥ%��xO��.%�|����G�h��V�vKX�n���eR)EC�G?�q0�&Z��禅���K!i��LK���i�5\��0�%!W!8�ڞh�	��Ytm�Aka�!�Y�����8af�TOO��

�����g=��
���"~��[�����і���Y�9�!�xNI�R�spo�/�hƏQz���,锦�~bEa�-`�$�g1c�%�ŭP�� \A�@OEe�5F���wB0`f?ў���Y
ZO�\�N�,u��h��n4�	������0�
��0k�3\4"���pꖞ�І��k�8L*�S�Z>*wwv�=�Y++�&�t	Sු/4��������%�@��~��2�e��lY�t�?�F'��7��I�]1o�_�������D$����w;��p�V��V0ZB(օ.�PG7���7Q �����6����8mhd�
;���GL+�bK��>��]��r-#�ӌS�E�*ab���WC���̴#�cqEE�#	�*#����e7���,7<6Af�fZI}`����9E�{<��?O�V�X���'X�y]���Dl^�<Bc��b�'�\�ŉ=6Ef��=�>� RU�h%kk|�Yج_v����?�I�����H`cKrD~p�?ޔ�(Kpj+��V��^�؅~�W�ko ��5L�Q��_]L��{q�n�6�_�&�"���S!0�� HTL7�A�^NTG�l l��F-�j���Q ���3�'�8�P��yu�2t�l���<�bK��o��&:��p��B�ە���_\AUe[�a1EB��|4�O���7��`�:�����0w'�Ҳo�5�	N���`�դ(*�w�H�$>/�`�A�E/��C�/��]�5tǷ���� "{��3RC:m4�{�^J�c���ka���
���5G�7[��j�K	ז7�j�%V��-~7}f���x�s] ݻxR�}G*婤V?1�J ���j��'i`4��zsY���:rr��϶�fA:�q���]n3�&:�>l��-��$�=?5͸�������� �S�zH��Zwƣp�Z�u$L@��59����:���W\�oc,��ܔ���|s8^�RVLOh�¼�*U��z�{D\0�u[PJ��������fn���U�8jh�ˣf]�uܠ��/#w��s�£*���g�-��*x����lL�"l�e���7���_G;1�a�� ��ӵ�^�'�;Rč)�=[n���*\+T>�B��?Ǌ%�>YI�J�����ۊ�o�'���+"P&�N�s��U�B��M��{B�A�X��h�BTͺ�E-u����I�~ ����鸏Sq��u��4 ��Y4ٳ�	K��_�nE��n���%��4��|-�����OC��Y���T��)�-ϗy�TRϛ�C��_!���}�XPЗ}�&L�L�B�a
�y�����<|���o���gV�q^�O�»�R�h���5�J!��Ӈ����}���ZT��E����N����*~�k3O������3v�x����<<�3�~|K��z���D깇:�!g\��wy$c�Z��7��hs��~�h�$
Z4��5�*���S��;}!wZ�S�}�w=�ƧK�noZ��	!�]��w��տ2�ǽ� ��˸�U�&+~^����3mq?�f�+ٟh�łP6������9�<�X��.�D�8�+P�,�/�����]��j����\�}�El�$+]��@K�Я��U�	R��r�_�U~W��=�g���Q���7�xkC� yĴ�?çxq�����!(M�=pPT���b����R;����P��1��cE��ڞt{$�x4J?�]�kt �<1���a�$P�ު�/'�v�]�c�>��ܹ�K���D�P��XS�p���2:�"��Hr��U�j�[��߯m��R8�X:�&����\�D��]�bW���14���?!s��p�9��`��vԬ����&��}0Pj�z��]w���O�N"�|b�'��_ӥF5=�"�u���d��Qښ�.$u���4\�:u���)�i�+���0Z�
���3T �u8�󽅽*f~[
������[r"|�ꍠ�L�f+Jm�vfU~��v��6<��9NZ��G6�H>��-AV�0�����-�f=��s\�.�&Ue�ZM����>��"�Oj7'�lkC��S��T4�B�U��Bb�ȗ���f��}a�q�}�2��9���X��c��R�
#��߷�V̭��50�w��8��ǜ�y��D�ɑ������֯~+�V�d$��sԤ� uĹ�~:�(�v�'�;��3��(!U���M���ZIذF�׭�K�6���w6l�ݰ(�IW���B����L(]�"�9hі7u��ͥ�dE9����u�c�c<��e�zf�y��S��:�zs��N�W;�ǻ���~@�ŵsI��Twk��2Yk@p5�ώWU��Q柰��̡g�q�
��8!�)ʪ,�Y����^��Z�)f;��f��l�B�Q�`�z�>v�V���Iq�«�GQ��q�"#pߖ%^p�2�.\�F#�[�Y/�y#˔I[��XR���[:ƨ���i��E+ (�t�^��$�U��K���#u1� %��H����Z�{[�ʘR� 3�_s�!��^�ĞC���U��%K9�,��].�Ɇݝ���v�2iO%]]z0�E���W� #�n�*�v� �RE�&�)x�M�.]~���Y��w�Y�o΢AݵF�e [�v�Y˹ש�$�Y-��o��+T{�%IF01��J?{��������O����&�c��W�>U����Z8z$Voǽ��xW<����Db�=Օ5+�?7V�y:ٌ�h�b}��9H&I�ӕ���R�� �B�<G��o+J���H��a6,r��p`T��S�r@�i��A���Y��Q���� �e�u D�$!o������yP)���4>gL�mP�:����I��#/MHa��+���������c(%V`2T[�0��^��Z���p��vBH��)�7^q�@��T�	KM����M�p!�L�?f�w�ى��Fv�pY]fU�ӷM�f���9�I+�]W�^����q��%�H[��o�[�ʐD���~�"�[��G�����l�Q$:ё5�:����m���@j���#��}%�+���¡l%���c�#�y
vB#e�r�(Fm)&�^;�`�>X?����q���Q�����̨�:%oΔ7d1	�b�!�2=6\�3ɻ��W�Q�%��F��ɻ�gAf�\n��:�_����k�ȅ���k���chN"�V��漭~�ܯ|��R�M���[������@

��	H��������wU�=�Ė�uA
Λ}	�d����K;���f��n�4#�ԏ}בx�����]{ H,