��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�&���ڴzk^�2�t�tC��)�/���KL:�kD3���1Y,�d1	��Rv���)�g#��5�fŽâA�|Z^���,~t
��/�1����,�ơ��:y��q��u��f���c� Q��:oe��ɬH�3UH�vF���=f�r�:��dї�+��{#q,WƐ���H� �ٞ4S�'.��S��d�#�qx[]<n�/�ݦo\�i��qN�ѱ}'��)%ʶ�6bY��+¢ޡ땲�0���f>A&��!Ⱀ�l_�K��&.��ûI�+���t�����.�D���|e)�x���[�xަ����Bɥ��dr�M^tgw�\��WC5��X�7w<'b��K�*���'�I���f%\.4���G�1N�p+�W�	Ѣ6��Z:�0(-����#��W�4fð�0<�D~����̄�fI�S�H���BU�����	���/D]e1��gJ��*�3��WW�3K���Ue<;�iv,o�Wv��I�����K��=��n� �܁t��b���� 0}����/��tu���@�I�BSXt�9�Ƈܑ0�r.��]f	��z��ۅ�͓mS��upX�Z	��T{yc�Vw�(��#c�}/
�#��Ї垻M�[���V���D�!߰�K�Ӻ�"HG��n�B&6��G�ԁ�xh��k��p6��s��"�I�>/�}�����{� d�#.��y�W޵�J�5~���m�	��*�z�Em*J�O����?� ��9��*��Dyz ��C������>�+�;�6>W`�_���6ӵE�]9�����D�c�_�˫M�a?LC#q��CV6ceHG�d*���[���S�a��}��lmuCc������y2o�������.�aU�`-9�`^ѥ�
6���'f�|j-�zaJXos�j�=��L]�vrsUR�x�߈ ��b�,%��
+���>Z��W�#�����,s˜�G�K�T�h� G���LG��R��<���Msp�Cc^�D<b>�4�Pؽ޸;*|���Ϲ�C� 4��}�}���垲;�L,tҧY�����f^Z����2Ђ���`��<�&�f��w�.�#og<����]�G&#����!����(��#�)�H��mX�&���tc�/�0~�Qv��jnMs�d傦�U����h6z:f�Q��d�#k��ӝ&?n�& sr'}�~�<��~���A�"+a�$R��:x��\�N'/�i��i���)�ѐ ��o�O�@!��,��ȹ��	,����{�	6�@bw�X����m<�Bޚ���-/ִ^:��}R��L	�/p��.B8~���'+v���X�E�QS�4�\ȉO�aX��/�v��V�Z���՚�Ҝ���
a�F�S�3��OZ�ZgEMBk���{L�0ٻ���Z��T~*n��Ux�W�uŃ�~a|ہ��ьlF�
�{5������~�u#�!�m&<�a�)/� k�e.m>xj*�WW��Q��gY��gw�N�/Ғ��� �ˬ��m��v��%,f�S�U)_�3��1e�#ݫkl2N<���t���*XZt����J`�Ga��s1��5�}��f���H=���F8?���u��.|��K/�E��GX�nȗ|�M'�ܹ���	�[�0���ǥA�V��n����Z{�fǙ8B�oir͕-�����"s�O[N��6�J�@{t�2��ࡈ�HM4�0�����'z��Q7:a��Tf_���`�
Z�<���>��H���4�b.L�d#���P��/�ȍq�	���i����!�	/T�������EMaC��Z�{�y�	��/u+ؔ$��{M&>���͆�[�����C�g�<����v�& ���5�ݪ7�wsו�J뙋En��0�6���]̈́��i����0!i%�6��I�o�+	��*��`���{4e/f���w�����"��D}��7ߪ�2�����1 }n�:��ڞSu�:��4��Xu�Ĵ�[��ٷJY�p(�
@O��"2�%XzL2<]3_��_���nc��T�����"�i�%JmS�_�KF��b(}�WM��ux{�]Ue��| ����Ui���1�f��	�B1ˡ��+v�r�`�d���;f;��w�Wt��*\b���U�H���_#��ٹ�WS�H���RYg%�/|C�^ϓZw���]�6����dTt��7#b�X��.��g��k��Y�0,�D�_w�r:�>�M�}���̻~zc\g�_�T~$x	C2�/�2j@��d�>%�XQ����]]���-�{�cD$�B�g�B��i]���E|N��>1j5 Ih*��m*d�#�76�"���g���9�u�_!#'4�S�{̢���q�! #����a��E���R���W�Nņ�l�d�E�S�cǨ��m(]��T��B��1��P�?<S�Ν���į��P7U6��$DT����WY���P�М�5�$�%H�,�-�S`��cS�9�w��X�z�3W�`qr��j5@e�]_Ǥk�(�楁�;g�1�{��2qS#�n��`^M��Y��B^喈����}��~�g���w>�������u�Eq:}�z���D�L/�z���A�����8u��Z��{�C�F�Y@�6�g��+l}R��� 3@}1':�o���K���Z ��W����7�M]ń��z, !���5��c��w-p9?��j)��!�䕭֔����󎅌qZ`�������w+�@1iG�w����|7J�1y?�E�LY�Q�Y[6ɴ
�p�F:(t��C�G0׀l�)�d��|����U�0�2�>-Y���70���Qjr��h�;����0�:��>��zl�,P�.Z�3����TT��)l�F���Ԓ�Ļn�Q�%���[�&w$����]\�󀁇�y��`I�I���ʢ����G3��5)*|I�Q
��~F؛2ٌIY=��J(ݬ���lN/�ɭ���`�T��U����!#F�}q)5	�Xç�n�����t�*�6��H����Q�'��f�ͻ/�x�{�
�0��s��ҧ05�sQ�~�W�P�$�Y����x=-+���e�wS�$ӻ�NOUV�_KN=�Ɠ�_��T�UA-t��M�DX�<ױ����	���Y]�h�E���O,1�8E��V�˪�@�^���-R�P��˻�b�K�]���#P�ʩ�3�!�aA4Fzg����NfSr鸌�z���Ю0��*�?�5j��a���X[V>�G�ڔ^��)���E�ʊ0�߾1��l���?㹡���9�Ǩz#�b�Z'��8�� �y�M��{*� �g���Wv�q����xo�<��N�v&�X�f/>~��xP4���u�6�N�%�i��$�i4es��w
5��`Ͼ�����DËg$ �Љ�Z.��Wj����Zhz��V��N�H-�|�;�"RV�9��#E�B�_��5��ݼ�7���`��'0>g��*e�����s�����5�v<�*�M��$M�L���#�1?՝��)�<��=3������k�~Ll�+��\�ޓ ��x�s\��-���^'��vm����~�K�)5�V���,���$L>?"�#4�5#����-KeYVq��*�λ�h�]I5 ����A뷹�Dsd˓>���T�{�;~�������V����Ćf�L�Gr��#\���0�A���v�
��\��)�5������1�[$Gi։Ah�)��I��1�Y�-�"��)baה���`n�ډ7Vpq�sX��iG��/���;����w{NI���I���;�}ϸ�l��!g�&j��Ǉ�1`�sa��oC��7p��Q�����,�
/(��g��<@V���xc��9�u\y���l�	��_`Z�O�����[���]�gYۓC?���ͼ�Kܴ��xs��K}�!���Uu{��:��C�Wr3��E�be�ݍB��7m�CY��Z($�(C�/D#	��	�k1���|���Yv�����M{��`�F���2����QM�ܔP-���+^O�&�h��������n�c�F�'[��^C��N��jޟ*�J��_� oez����)oj#)j8ɧ�/z^��-r�S���U:&x�CD��,ď��J���g<��Ձ�HǓ��g'�؀���jE' ���;�H}�˃t\��w�����g�����]�ْ�;W�S+Z������5�`Nx�3�����rFv��r�9� ͚�>G)�6�T��(b⏠c���J,��.=(j��wv@����(�X<�`H8q">XيI�aL�A�&�m�p�Vp~��#�8 �9�^�H삧rCE[�?;��Ky���ٸ�X�����	Wkr?�o���}�N	��!��ej��i2M?���,��v)cY^��W��l#���ĆD]�QC1�Z-��WV6M"Ok�9�oӢ���Xi��]ĸ̂�k���\8�\�<%�����G�U��b�	ɂ�;��/�7ځl��r�7��IAx�Gz��>n���~��f'��0l-i;���U�q�c��X����3�S�@U
]�%���a�8z��J�B�r��M�(�9s!VR2I�u_��5�+zc�v�5w?�P��гôZ ��,�����PK3��������@�1������ML�����Y�=�T�Ub���L��dV���]��[o5�N"�h>ss�B�s����b�;�k�A��G���1��$��x�m*�F���b2�(څN_s7~�}q�iV�dH�yb��;oP"�������T�qYEߞ?ſ(<�-1y����=�kE�X��7�MU�k��s��`&�!z���RtP�����;�ٔ$�iI«��ҫd�!uNHw0�Ë��";:��X"�����ƃ+R�A���J���o0���3=v�K/(L�����h�>X���v���k�|?���SŁ[C��i�-��AC�����o���k��C�=�,Q!��=
�������d���w;}K'�1`�Y�F�ܛ���VU;��s �0E�c<!pp(�W���G�[}[/�~*#1�jn��ĵ����K�f��A��Ga�n���gLX�T�>��*z1�aVJE���
��ifg�R�D�o���H7��mj��w��t,�Y�c�q6��) 4$�}Eh#/f�V�ۙ^*W�=�?�WL,���{9x{#�@�4@���Z��� ��~5�'�bZ�_�ɪEy|��
���׫}��W��Q�G���t�!ʽo���/��c~��A|�'/F����P�r7A�̖�'vG�c#�3�1�6����]������8���#�+�����Lc�0�G��T��<�-�M�M��, ��ăou+A�V���G7i����w��5l|ހkz�n�;�9}f��J ?^�,����q�
9��P�n${�J�tf9Y{����}s�m9�/���B�wV��h0ƈ�o���TN����-'�+O2����r鹬0�w�!�{U�N�D�N�8�B+]YE	ļ���R�LH\l@Ff<>:����XZ/X��&�n�������vX��tuўS�P3XZ�����M��^�Q��[�^��0��i����:��+L�?�1�o-n�h*�k�r��,�4�����%!�;~�D�7G��8�Fl���V�Db��b��ߧu�py�t�fCYJ1
[�K�*�@Չ���q��ݜ��آ~��C���ά�5�QP"υ_N6���Yz����óC{��6��}��F�g��J��,C�PQc	��4njI'����{�K��Zԫ�~V)��f��Ty5`�����~l���3.�F���N �!Ki`N����vF����\C�IF��H�q+Y��o.w�t�y:�"85Cj�r�m��4;H��8Kl��y��}"��1��i#6��s��.d��?y��*��1�Ǝ��1�3À�u:��E�x�w��`�P���8���b=o�('S�z��,�蓈qj�.����o�;�
U�4��/::I#@�t�^{76 ��G��wSI|TĂȉ*bJibJ� +����H�#�{��A�P���t��7�a�R���*����S��\U�!rM�;LT�W��ibu�>bgeC�PT���a��4�a��X�U��8��0�A�?�d~�aXӟsw���!jF�|��/�zjq�?W�Bkb� ;��I�^0K��eU�\42���f;�@�L^m���PD�~����Luq�����$�PN�