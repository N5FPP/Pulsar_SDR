��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�۫k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A&Q>�Mx�E��K֎�>v"wTD)3�2C�
!h׮X�L��,�*�� �L��>"赇�b���6��72-�t��x�"p�0%N�+��<0~#�Ѣv�7���&�0��<��;��_6@;E��75�":,h��O�GD��ce�7G{��Llr	tS�����F��#	/GUv�}�=7*vBx���Q 8r���~Y2r𘏸�${o��qaX5��P��2/�|��f��,}Y�(\͹����4o��p��v�*B����C����~@iK)A@���Bg�n
Z�.�:���L�n2V��ɬ�z���};n����-�U2�P|� �ا��#��i3���U=5�
(q�p0���bM�/\J�>M����S��#l�.�������K������u-����7�7j���GBJ1�a8�o�x2��<�#-���L�����sGq#���0V����ul+�I��;�YA���g��\��=�U�-���[y�/��x+уs���Ԛ�VF���/��T�3j�L��(1�bV�Iq�Vɍ���E�ʱ������6,�O�f����B#�<�ED��5�!��
5���7�?�y��~��_��?�Z�0O,qk��ݍ�k������j��7dŇ��$���/��i���'A8[
0Ю�l�-o���n�w�#�/��:_��;vZ�D����I
w7�#�[���R4*�遳�xaX��X�����@}M��Q �Q�/�?rg&ŵ��6���=(��L[�<Q��@�����rzb���/���=2�������D$�����&�9�s?�����\�m+$Ȣ��|F�Θ����S�)�)�`H��3�A��ċ�$��e�����`����I~��TE��\�7JQ�a�#�QU�\�H.2�g�^���h�E顱���iSe	pu�H�nv����^RF7��Eg�/*�]�}�J4�w.{�OI�1:��x�`��� ��l�=�)��g �Z��Bz[+���	}�"���'��H`�4�M�sz� ��GG!vaV���s�Ue��h~X=SBD(�6aE�96	fv4w���v����^@_�w��y�$��ob��桨X��v���
�x�c!�wW@�e��떘��:�Q��7�TcH��r=_�譢ÇO����}q�f��Щ�B\HV��Q_K
ck&�/u��ifA����R�a�%��ɘ�Pr���n�7D������v�x&$~�� ���E��\�@^�K�������)dU�SҺ��4��=�i��2��c#����=�4J�l��y��R/�6���0b5�dz����Zr}P4	;]<��;�a8��Kf-��I�:=]�:4I��� �5oq��IJ�vT�}MB�?�U���IX�A�U�0ԫڜ3{��ҝo��Iu���Ｑo	���6��E���d�=�p,j��c�\{�&�:�^��q��$��'9�t���'�]M-F�uJ%b2\s�L�Q�N�����ǩ���ߞ.MY�Zs>�