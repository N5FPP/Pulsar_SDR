��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|>�qT��>�z��
�����|�L愫�H��ɺ�a��w��$�YF���bںM_���,�0>��z���H���P�0��C���[�;vJ׭Rj.�
�1�?��a�IX��U�ܰꨮ�\��;(�Ee�-V���%��S�I)?i�^ׯ��'@��Vg��?��w��(~���R0�u;S�}�~�����b�'��}
{k��w.��Ⱥ�q��g5;�y�˿
�#N4l���IN�d��� -�� �^A8G4���$<�^5fa�� m�o�4��bml		��2���`pb�c�{�
J�F#�K��2�9������(��L�T��6���UV��M������S���o���-dq���zaT��'�{n< ���
(I�B��x%�ǡm��қ� x��(;�b	�Z��W�K���O������R�c���?ǲdb6/x/���\�ԥr�n��b��^�\����N������~��}��=~չ����*����=��HL�e.�n�t����L&-��P����l��4�nw��ؙ�瀕�F�dp�#�{N�2 ����	�|R����<�1z~�P��A���"�)�U�,�T#�L4��~��Dg������XEx����i`��"�y�|��Q"U�S����vv��,���73�7j��D����p���ת8H>��[0n�ky�˦'H�B�n��_Γ̒4��0��#��~A�8���A]U8e5�Y�S%�&H?�Ү	M6�\3@l�@G�����*.����3j�Q³(W?�����K�f�a,�q���j���G�;L������W�'�;���C��ヌH>SN��ۥ0g��֒?冠����8�T��Zq���y�3���]��lO�C0hI�zW��Fʰ�Q�jR��7�c��϶���R��f&�l�IM�+�Q����/�����֕� ���m��ؙ�z��{h�=��^�
q��T�L��F:m��P��j���rb,5�-K Z���b'�ۋ}EW��N�Jr���$��ӷ����{E���=U�X�~f���&JF&�ĵ|I��r��'k#k�J�c�N��}ጧ���`���қZ��^��_r+oV����|�W�*���|R�4������z��#r�#�a�����uq�Y^p��&�?�$��5���z�\���NA�U%��nkZ��d)��fV���:
*�)�ƿ������!�~�[�?Q�J��^���%�uhk&YI`�1��>2�����R�RA�Ɓ���͂�c��t]@���3k;N{�#u��g�Ƹ��̛b,}�7}q��]J�M0--�ť,h]'�υw�P�w�p^w��!��Q��8�Q�����!	*�t i������j�O
<[ c��c������,ª(J+�\��Zl�E�a5�[���
����ֈo��h�z��qKnh�iC͇:nT�Ԁ�6�����8�r��8" {���_	hd�31������O��H�xyi���+:[�|�R���Fd1���ޱ�AbWIav��ˊ&D�}*�H�R�2
��0��TY��U�����ʆ#��n�֥�?�����2g����� �d:��9�\i:Ww0�6NNi5 �Ī�������ukj�:B��#��&���>�Y���J��h��lX]���'�UL-g�^٩_|{V$�je?���^d��xZ��)��-X���ka�;U~-�U5�T��w�*��]M���LK�"k̄���.C,��tC���k�l#}�fܪ�u�Y�-����5:I�%Q�X7����;_R��lO��	�e�ɯ� <YZ�Ep�l���(Ƴ'n}SKЩ��s� ��|���9�5Y��AW���Pfm�����b3���O�S����W�L�����#��QH}�:��3+�^��Jo�п���d�N�%)��՘�NśvDz�",qYr��
���n6�y�7G�b�хw+j�H��3@�|�8`���!eC�g^�E��� xwͺ9����x� L���*��덏��b&������ڮQ��K���JO�P�v��������k8(�������A^�r6�?�C>��=����iJ_3�9v)35/���ݜ��/ t]/�`�9��s`�é��1r[[Mp���r,K�>�,@Ut���5��e �}�RKm�m�T/��<�Ͽ��6��+:����=�-e3��4�u��1o8��sv��o_�����p�{)��o4�<�� * ̇�;������G�K� ���q��9�� )�����e���I�y���Xb?��m����U�<d�3j�e5�q�i���҂A���C������Rۚb�\q&l�������;&��tn��"~ݳ��A���9�]/D��W0-Ĺ��U�C�7/E���뮔�?�V�[�""=R��$�$�Q��C�k�E�l�U�]}��L�v�=�ԇ3�_t`]9��ߪ���H���	�O]�kf_�$�g��eP�UQڪ��P��z��`� t����n�m��g����]���qt�o�j���޲u���[�M�5g�ktק�}¨�E���D?m�N�����x,EF։��A�C��[U�R#����'���>q{��8Uzz�Ϙ/����`�3�Ō�![8��^ �Ի=I�;|0(�=S��=���T�d�@[[YA�e��r�y`��͙��o����r��s���:����O6�g�mec��L�}���abz�&�h�WD��5s3%ݱR>�b}��Oj,�O#E%��u&�����D��g5"��*Q�x_Zhnn�G =�~O�WFߩ˧��7�8OL�*�T�q��M���|p�׌Bp"`��i�&��R��y�G�͙��+�Io�Y-f1��h������\[�
��m.��T)�҇G�7����U�l���E]'C�t����Y��r���U�y��a��r��+F�t����	9�>d�Ǫ��q�=�$�Y5��¡�>(5���zA���Z�s�s�y�:>�Ϲ0�9�I_��1q���S`ϯ�ؠ�:��W�̒z���s+8c�s�*K�1����o��(����^�(hQ���dY�az���A�Ǿ�8(p����L�R�c)��K)��?cҿ!`�0_�bJ{Q�G�u��@2�(��� �Wl\(��(�k��r������H�o!�nz����L�����L�/KX2|�HWެ�^ak��|���Cg(c��վ���V�B)���HN*��ˠgaSx�ӂ��h`����B+%��Gj��y��X��χ�rU^�>a� e�rȃ���h��cg�ϴ�8I �
�yÿ%n�kH�~E�1��:<zGqqv@�~��⇝|PR�U���(/�N����AW&G���\��cJ�0��i��i[��̕1Cf^��%x,����c�R���8�����n�x��j}UwXK&\n%R�?}`\��>}(�V�W�5��U�60��{j��u9�����+�R�u�����ȴ2c�V?���I�B�MyΆ1�VU��� a��/m�!��'F�/�{ҷ�r���Rsu7]�q�N�tg�(D���+V�da<N#ٴ��Z��=KI�ZY��d_&;�_�р��R�&7'��N�e,�,�]*5IfciJ-g�<(��"�-R��Y,����x�j��E�pE��Eg�m�,`D>1g8r܄^%f�����{]���Ĝ~�F�"1g]-	����({&�h��S8�v5������
��gBTD5ʲ�X�S�тm���R���	�M��͹�Ė��S�<�c���h�y��?�d"�T{�Y%�N[�	z