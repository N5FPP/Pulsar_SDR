��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��e�ik3�������w$����g|��J^]� �恼S哂�O+z��p�˺���pd B�O�v�q�5SK4,]zO�=���pۥ����ʾѶL�ܕ���rtXi�5�a�K�~�Q��mծ��9+�LGx��?�[0ϭ\��mL�Cq�I!mhр�ҧ9�1��s�ԣ1�U��;s*?�~�.���D����S�e�%4�RqM�&I��W�_�b�n��r���~6S���Cc�� ��e�V}����p���d�!�'��t����G�^�'!u�;Lܶc(U\i���ؚ.�	��\�C�0F@ &&2q7��d�4���MxC���I'��'��&�}QXRE�g����ob�q:���W��5�d�I\��~_�ŝ�b��M�[}	A6(�K�;C2��;���VA���5���bl`��{n����^� mc��R�ZpS^�N���?[ZI����ڞ��ee\����LTn��g�)�ک�6��5�_c����N�JyO��}ڒL"�����ܰ>�D��=H90�՚�X���ʅDY�J*��PܲC�:V��ϿEa�t�7�$R�]Q�
�ep�I+~?�B<]O��
��'������J){QGڈS7H���k��ګ�<px@�;14=���AQI@����� 墴IQDI���j���XOx�&�l�.����}[�a7-p�/Gtq���?�A�E���y��m�VK�y�o�|�����(8�AJΉ��6�V��v�SJ���c/Y�;�Ԓ�N�&M!͜i�*�E�nhO0E�h����j���	�1�~j��8�6�1�UDg�n�nuް6��(m����:��~�D �1���>����3	3��l��kp�5������n��l<f�Y�=�}O*/���w����bib�[}UfԤ)�wo�}4�Mz�q��mb�%��/�
���|0qi<-qn��w�0c;���O�O�f��|���p+�|.�l�&�Z����}#r�(E�KEg0nƬp(��X:�X���c�ʃW���Ãړ8��(��1�F�r�ܥ����Ca�):YM��X�	3�!u�����<�C����*���ύߝG��k���<�:���t�Dqi�������^��NX�r�
���1]���].���ee�@�{���e;�f%�i��:��
GD1��5¼���Ԛ����6�*�Ǔ@��m���y`�h��ɑu��p:V0��W�#�]�ڳ�y���lNG�@���z�����x����<Rl*�H�cVL�q�{����S�7��u�g�GU6ׅ(��/��[��0�eX�3�sK�*�hK���w�	����(b0}۾��`����4O38�0�#`��Q����?ː����b�wF�t���v9�;yI�|E�)�E���π�E	A�B����؏s
b0��t�  ���n����6D��]�	�� ����.[`nѲ���je�K�Ց?˚�P�����	�%P��8�4Q���?���L�췷�Y�rL;�����;�S}��>��w��G�����R0���uq��T�^=}GB��5D���ne6�<��������`����M��3��s�z���-ן� 5'�py�G:Ψ���n��ώ��T�L���>_��[|��r4gc^B�%~e��z���OG�}��~����Ӧe�2c��c��I�x��s	ꋌA|9͇t^os�V$�)ɘ��^P����v���*�6-	�x�b���l�C?�`@n�7c���x��:4�ڻa��������M.�]"�����g�y��R8ѐ�b�[��;�z�&X����_};��}^P*��q��L�A�_��3�<ͮp��Ry��CJuKTנ���-����_�lmޓ�p�;��^�Y�*//��T0?u�$,`6_e�r-J����y�LJm�,i	l]uW]<"����7�e����aq$F�+}�W�(��j�sU� }���(x��vz����%�it02lʓ�V/���&M�?�M�&wl�s�t�����MǡM�I'��Q-��7�e����=�`ݜ�HSq��{�i��%T�2�#��"�v�;��v�����9=��{s�s�ȩ_�0"a�)�F]'�˧w�{�e��ƹ��2��`K���8}[r����m�|-�D>�vM@~�Vf�~�Y�@��5�̏���a�'��]5m��l�')(b&A�0�<�>��ꄈ���8^���Xkhk^N�g��q���OCQ����)}�,��j�y����ᣌ(���2N���6,(��>��V���*.�iĵ�	���A�W�&c�/ǴHӕgd�]�4MZeKm��;ҧe#����;���7��a~w�O]-�L����+π"��"~8 �d�~�~�t�$d��zeG��oj�Ϸ��B�C�bDD���r�����=�#$�����,���
�Υ��,���/�E��_/�t�ڢ-}�Ԇ*�F]�� n�w���	OKX��:⛾�n�Yn��F</St_�U�_y��Z���A��HӋ��&R[5�M�%CBk�.BU84�5�g�t�HE�מ�\�r�5�P�[��>f.x�`�N�\��傶����i�~�־��y|�����T�(E*	R���.
U^��w�q���E�Sy۳:L����@}|���s�b�"�-
 Z���,{��}�W�Oy^�@�iI�@P�p�e��+�k��<Q��B$�<U
B5��6�KT\&\��f/g��P�� ��x���Tr(�q����c�&�H49 �;(��!إ	�rk{��K�VpѫS]�,EV
TEN��lk-9� `���AT�6�wp��߈�����Ѓ	c~h󒬌Ѻ�d��*��N�l�,s�����S_=�ٴ朥ƃ��@!���4�d?���AL����{�e!�nSd��
��ow���X���О�	ܭ�T)� )�_R;�#8[�A�]�ӱ�>F��\��
�ڳ	Ov�JNڃ�����^�CF�R?5_5 L�y�%�$rPO����x���l�� P��������e�UBu���6쑺;-W�������P����;]�·����jn��� ��ƣkyZ.��A�]h��I
K�XS�}�.Ilv�����y�@7'p��;��ȍ�@s]p#'����R}'��BXn�-�n�ړe6&8l��x�z��+�VǍ��5ـ��b�O�	��=8S���1���J|K���#�w�1���ƒ:U���6>��H9��Ș���2?O��[9 
�g����7�n�����S���)�?��f�b�����x���eXa=�9�5��a|E���)r,�gnA�"(�/�<;ni!�ȋ���n~p�lV�R�A>fųr ���t\2�+/�~�5�"l,�
HJ��C�H��ɤ�ױ~����!��rwZS P����w�\�$/2�k�<l�*v�7����s��D-���V�;��yA�����?�,��f+,�m���د 1�<�8.DJ���D*�\�L[�^�}r��.�d�M4���y0UF����6�s����KAޠ�r�]�����|��!^YlI��X�S^l�[���9�LF2)��#y�G��NT�:1o���dh����Ba
��I�����qBR��o���B���P]��<9.Ŕxuj�`Z������9��|aX��I�R�u�1)i�����:�CE5,��7?*��^a��oa#C�潦(�����T\��-,iX���J��/�!&�Ѵ�Ȱ.!���s#RMm\��	�������_�g�ٴ|��Џ��	1��Ս�� O�l�+Ԉ.�"��y�wKg� cL�ݫr����{�W�i�w�֪>����
�5� ���_!�&i�'�8�O�0��:��$.�o�8��P{XL�!۔eS�,ʥ;���{�f�Z�:0��޷�MC"��YF���A]�����;t�����C���`R��	��8%l�᜗55=S#�G�Vm�-��U��n�'�H�D��R������!�G{o���ξ����<~q��ˎ�bL*T}���p���۵$�{|�_*�0;5>�V�뒋��u�7!�f6]�)}x�T�����}�"ú�������[��>�*!k�T"�������s�e:q�"�����)Q��-�����`��l��
_Q0%�|��.�tk��J��\����E��+F
g�@�[�^��-������ u��s�O���쥸�Q!I?�kd��g�n%�o
�����vN�y�0Ѕ�)������c���A�<<�F]���E9Ԇ�7�T����.��8����� �Ә���
X2�%����o��J���'��#C,��[��He(c�э��`b�$�E��m
�$4N�\��sO� �gPiӦ-c5�*��J��}$љRRI�8��ǵ�R�=��YHF���Q�j�a��7ڛ�
�%��������G���l��$2iڍ\�pl2zChua( ���).;+}e(S��P��Lԩ����ҋGsΑ[�Q�L�GژA�Y
��7�R���&
7����`����a�'
K��D�Ǩ�O��~����������Au7���ߍ3<Q1B����v�7���G���3���Vl���Tsi�����Y�����]���f�{�qO~�~�=��7������X�c��d_���G��vm�|QE?�6~ Oɋ¦���}T`���� �2��t�(�??8�x�:z؝�NI��#��G�9
e��ؑ��a�n�)k.��ҽ��Y��:�u���є�z>����m�����nAf��Ouf	�����iqoH����m8E����G:��U*���)�A.�ɒ�sPr���Y�ݾ��@�Y5"QSoO��C{J¼ۜ�e��@6�p��v?kÒ0Oe�P'�u���?������� ��^N<$�к�;J�]e5N�Ӱ&i�1����� 8�!�-7�����s7��	�v�%l4Ac�ׇv��DR)��).U��kK�6�G}!�>�̩+3b�RcA����q'ax�X�`$�W�qpձG�-�$4X����$Cg��Xq.�7B�*d���?���)���nR��Q~Un�ȨfkA3�&I�EK�ն����z7�j�q�1��T+09��ٲ!�VЖ-���,�?x�k���zE��4~s/�Im4vC���0�z�/?2��txY�pބ�]R�`;�𿜬�Y��i�M2?_�,�k��b��xD&��p����ك>��4�ZM	��1l��-���D��v�g9_��T �*ߩ��G��� +	����R.�7A��Ī�$�N����'<�W���k_�����H�~ΡӠ�HDJ�D�kL��*IRᢻr�$C�ĺ���nuŔ�edh��lؠ��cL^��v���;X�9Ca��T�g����]���dq�&��eZ��QPXR]?��x�f/���L����&�-�ʟ}��*���2�z��}�Rn3PX(��e�p �>5��ۍ�~��N��(��$��p톧/7cHs��T�ʘ~�p�o��X�Q�l�xgH�Eel�*hjn���F	��b�e,o�������6#�3Lsd��@�A�o.�1�y�Z��Dۺ �+��U	��.j�m'����L[�SP�Y�y&ҹ,�����848�NN��p��')�Q�Kd���*{I�$U�J��ϭӭ���r}P���<߃^�(�,!>d��^I�S,Y����%��/�\������Y�������k_$`�l��)I��w`����zj���F�����"��7��!$���CTf��N��,��@%��<�����.���`,k:x0�چ�FBv��{�P!m�?��j�[-����ݖt0��f��5�!�r���T`�#�OH�h��L�1�?�����Uq/'k�� n���S�V��X�~�h�'���}��N������Uf�\�!�i�B�I��G�[!x]sZ����u�jiӵ���xI�!8���4�!�\� ����S!3�p}�������8�7����-�S� '���y������]���ǡ�jC3�����~�PR�����`��X���)�#�z&�6A� �զ��]=����$Р��i3���(�H��m��V���W���������kg�H��@s1��1�>��R�qn��+�%���p��%1T��&�8�9��#�h�L���&��.�I`�PȂ���I���P�����w���,<j��u�6�%����Qgc�T�q8�?6�[/,QO6�8�z�c��oCX���	��j��ƓV�V +�[���B7��f��%�F�q��C���A9�s@��]�
IS�a��ha���H!�0\-W<6rNĎ�I�*3�z�r�p��*qi����3�bI#�ŗc�jXk���>�	2��|\��dV xR8�t�vD�;CO�����,�T���(����MjleJ��'n�00̀ߟfZޤ��]�V�?��>�$1	v#���~e�/�B������m<l�����N��9<�[�X5Է~��O�']��<ڬ��������Un�Q�Ί��&��>�^�p��I�Ƨ(��Gr7T�=�~O[ݳ�ݛ��\��K�u�3�c* ���[u�1�'0�R�4����榟�9j�&;sh���r�4��pX'ȟ5;���K��MƤp�[���N����q\�̃Șg�i�U���.:�~�����7�!���59 �dSu҄���;�aU�,M���\V�̾��753��1�g�>iȻ\U�M)Ʌc|�L�K��/�� Ta����}�eW���&n���"�%�H���Rl�:�0Ef�~�_.�����]FUn+L;h�Չ,�]�����$��ea2/*��D���m�	�w���ez�w?i�9���9����i�5.��eF#�ys�L��/QL\m����!�ܔ!�F0�pPK<u;�V*R«Ș^~ڑ�|����x�;bwS���͒�,5/��D�:1)�W���B!�l����������m(u�cP"���!	�S���$܆�a;5�h#f�9�7S�J�N�_��Ä�f:Dy2�$y�U�#�Gk�P]�䴁H�:���4�2;�-7��J��� ��37��]��q�ܥp4mO�!$�u�1ʷM���cġ����|�[;V��N��(uV
~TU�c�u*�޽�O�:k�tO�����V���~S�z��r2�C�ޖ'[�Mz���g3A���_"�1̖6���M�a^��3��h%��ｔHHaI��Q�|P8<��FO�I�+�<1�	�/�:*'R�� F��B��7HK�t�Ug�x�I�k�:�����,�F����ݕm���6sL��[���T�Z�5i�V+[��Z�wF��A�>�����9�g�����2�ؖFfS��
��8P^�"#sI�����Ҹ��r(���E�#^������$X�~(���|>`�`��w�RA�kw��S�e��p7��~��ʻ�f�G|��Bz�\1�My�`����{E�M[�sŊ(��S7Q�^s�g�ph�:-Z���j��p�K��l�V9�`&� �,6�@W;,4�A�J@z�� x�ބ$�ޛ8���� ��E&Q�R�p^�3����ݦ�8p�f�j�	U3͏m�wHMД���/sCSxt�TxMɃt8�{������)�̩bۤ�����C�ϕm��Vh���/��=�Z�E;B�֟��Zw��Jh5<�M�E"��d>�1DM�����-%Q��K��0s�����99��4]�f�ה�`��դ�����8�.��9�ID�.���9f�
�K,D�D�<����	����8�pn<)nR��9!���kCK\�-W�{��{D#�=Y`�4uH|�Em�QX�@P%�ю���GgK����&'8�,w�槟����A�P'�z����*����$�j\�%���ug�ͩ����BT7M���qA;ƨmU;^g`)�L��e��~i�Cfc�������Z�{.~�8P5�˩G	�HP����~^w�̈́��[u�A�@��JRH�R+�X�\�AEp����ML��z���ZT$#�Ҿ1��f�Qc�ه��b���>�0��0�������xUn���Z�[�]�3�	�
o�I����Lr��t��F��_��f�P��q�lJ��&�.��G���8�~�]�9ʜ{d���)�M�O��u��\A+�.2�;���p����c�`���?���j�`�"��3o�\+��_oL1�{h�n�A�(�Y�c!*gn/n�A( w��+�4v�v�D�2 ���wҜЌ�z<ֽj�i�Q4"b]���0��\M'��@���^k��?����3St�4�e�b��bU��פP��'K\ J�yk�aa�^��q4ydG�V���wN�'�����_R�b��3�#9	���z$�$�Y{pq�ںn�(vS�nn���4�U����3��(��x����RTf�e������&��mW���Zc��
�	��/R��뾿�6AG9�����/"�$�\D�x���\qW�L�O�'�L�}㧑����[�t�3��+�icl�,��2�J�0 z[��6��7���=���!=Qݵ��g��)q����ʰi�Z��x1S�R��q��m��rβ
2����S���Ɨ��
���;�ww������_���S�h�X�<0���?����/���iu_G�)'�b_�XD�ѯ�Ng�ݔʲ���de'�`�A&�n��'9�K�)��~i<���M�0�OC��{�(4Z�/�V�w&�2��Įf�$nhn��+'ܦ�y��ܬU8�[��aN_�W�I�]�l�ۀP�Z"�FA�B��/�%��5wBg�T������  ʴz/�(�?�b0��kN��|���)�$85��ؓcsada�K��OA��>�U���
@�	l�h�Ǚe>�y����h(#���GT�=z��͗?�E�B��2�+�>����P�('`#� �)�,��vC�Q^�r���l��c�3MW���#��^�>�^T-�rY���`Em���Ϙ1���FeJ��Y�Cζ!��	q�=?Yl!����"#���9lz�0M#\
�� g�5�������������MD*��i��b�����/r+	�`LR�w�[G>t�9dX��p_� IE� Í.5�T�p^fǕYm��}oD���-r{̕���$>�=�|�*Kg����|s���q�� �|�W9�+y����szX��L[��vni)r�����k�ޣr��J��˂��Y1>��)��Ԅ�|H\�w'т��g������y��"�g�䠱QY��"������,ǿ<7&���\I�b�ȼ�Z��NA#I��8+�Q�T�Q������Rѡ^b�_����V�Ҍ���B�@[��.a)����\�2&�ϵ���Z��P��>c�|��a�e�G�� ����3��F|��N*��`˪`�u� �Lx� E��%�D�)�t�~+�L�݋ì�ڗ=����i�]�ނ\���m�MP$�n�V�M���a+]�ٺ�r�Zu&;�␪#��A[�r�H�f�.k߰�@2�� 1�����%�d2��Kϫ`��7�ڀg�k�*�PnV��%`�����Gu�>�i�iQ�FF��f��}I�ߊM��i�@_y4�"Ft����P9 
#7^�q����{�&�WjH@��e+BLJ��*������0)?V�ͦ���k��%s����c���y��b��?8ؗ��Ht�ޥ���q#���>�l�ԉy���k�1o�����ӀJ�>¤������yc$��[A_�{�����R���d�5w�T\sM6���>�f|��+FQ��f.�L4�c{^\��H��f��7|2�}X�����G�V�ԧ��{�G�Ԥr����9'��1�C0lÑ�Ѿu�nA럸��LʓM�b��`�t� ������e�~����>^�rw��+C����X�k��Ի���%&��(��Rr�]��L](�n*N~;��}�g�� �-�`����xm��ت1��6�)�?IW��M��ۗAQ��u,���9�wx�0�N[�K��+��M�)�S?�m��ϛ-��SU�tuJ=W%�.� �BQOI�.\�yzK��V�o��g"_>4�ˆ<�v��h.����=8<�u.�',ڇ-�9s*����]w��l��ʂh���IA|r%�&�Y��0�D�&Ҿ(�t���eiM�a{�:ߞn���>�ή�[�#@�j0������}���m'��a���]V��:d`����F��p�O���@����s�����BY3���x]��쿾J��t�O�Z��=�M��-�pl�qG��9��Ɯ]��?�Q�g�* Ku���8���$���	}1&�Y��61;j$�z��Yi���=c�8n���J�3Dq�����Yǒ�^{z�.F%`B�����H���T�z�t:�E���u�tX�M��P-�+VC�mۤ3��l��jo�������.���n%?x.O�<��1�e�6�jdIm۶�������B�^�h:��q�ߞ�^{u�܆C+���6E7�I���1f	˕B6�+ʂ�'��{|d�ßwܺ��lq8��_�+i<�f�d �$ϳ�?����qvi��N<IՐ׏l*؈��|^��v�6��3����K�]�^6�g>�8R-+cm�j���c��3�W� s����K���޾�� ���k(�yk�f���{��r���k���˿b3C�V�����{��0᳤"C��CQ��^�{���l�ޔN	�ڏ[�&�p�w��]tQa��X��� ��Y��]��K����$a��hX��t�ӷI2��h�-����[N�lvv����B�"���F��$?#��0�>!5�s����4�[�ڌb���T?M�����s��19q����ix�����)k�iV<�&G�t���v¶�S'���w ��:��F�Jb�,�S���MYO�+��+�_��RZ��Z�i�w��pT�3�a6�����*�ϳ��e���w��G-��=��>�E���Y�_�2�B=�gC�E��j}m�4g��[��kQs>ί���o2�����:���t�Խ/
?`��߫�$K�\�u}��ͥ���'��	�2��p��̾���	�$������R-}�fR���q����ҩ5u.�o��h�C����<�C��.�4��̔����g?�"g����@�+W_�Lͫ�5� r�
��Bzy� �m�ѡ�!�v�`��<���/E��I&+6vy�|����|+�y^���C�Y5���Z�*��������?u�Px����t��:pQ6}��r�Ti�Ŝ�<ǧ:��z�ѳe�SaHk��\��TT� h��չ��	�F�V^�z��u�ˤ^�~�A@����/�Х$��Mf#�s��톚(�R������|���|سHr��Z��]�zD��x�������"7�xa^�t��?�Ż�����ƽ���w��Ptj��jۺ��_�h����D1�\ru�
`�?���1:���֘�s����1��R����˱�cq�c������|f%4S��'9�p��D>	>��0��|�ܭ.g��ݍt�C6ǃG��&ˢ%e�����I摕����_;��Ϩ�5R���v(��뽊0�KX��U�OB2�V��tCP��&��NHjP��K&�	u@�S�B�����Zզa��7ԧ���~�C�����^D�!X���/��=+y8n,��~�c`��O������ho���\D!ѣ��P~�`�|Gg=���2[�ԗ1ϒ���$�XƜ�b��6�����D���7��q��E�F*-�����P>+d���&E���3���u�d.�^%=-� �v�Vv�ԍ�яK�N� �����1&v�0�#���K(̙�l�O�]����,zA1)�&0%�IC����Z����NE�ܰ�M�u=3u/A���o��>S��up��hb*C�no�?P��q7�!��Y��H��r]قx����9 �t���:z��89�e�7|JJ{.@pq@�\�3�S]أ@�����h�Z��@bpҦ�;��\3�)�L�6P���yK�t+w[=�E��Jm�ߴ����Ķ�<w��Ap�?�X�� �����٦玐G@pϬ����Y��Tg��><���@�+��үr*X�&�ضش1ϲ�&�"���E�v�^/��#|Pb�\6��
�m�FN���Vk��~̕���:�T��St%*�ۛ�sR���ݦE��W�s�:LjBɢ�#!l�2�:y� {:h�	Y�������K�Ϥ|�JCU��s�r�@U3L��P(U +�IL>oV����������ܛ����JJ	���LB,�r���)%�h�w���Vk�����N���r�c��2k"�u�XtD��!�\��O�H�N�hh�)v��
�;4t~'X;ԇ��Ky�:��ct���g��|t|Bd���N4�i��d�K�m���	��&�~��$��G'��Bv�*���RS��/�N��s�T�����$����b+0/��.��<ކ��F�g��qR�Z���+u+&K�����v��z��H�`��Lt�y�6��d��ѽ�)KCY�@.f�Ȝ �oƸP�7,c�f^�����L1:��r��,����Vz����P��ـ����|ǫ���L��y��:op�j�Q���`�o�(��:�1���Z
��{	�����C~��mpͿ��V������3X�I��I�њ���{ޫ���͢w�Tj�Q�g�$	0����/���A���0���]������O����<&.����e�y��
u�B/��2��R��Z��Dt��?�/zI�H)*<�_HU���Vv�9a0ճù�"�%l�� %t�js�1_�ex����Oݐm|p\J��BS�Fͺ�}Z�L�k�D`$+���9�����`����jJ�����s*8C�>R_����A�WD�He�=F?�E G> ~
�M��]����b�>��E8�x�*�h���|��,�g�-{�2b��*�ߡ��y ���M2�IS��=��������fs"�̥_��7�C�%����J�F�F@���$��~���A׹f!�Rʭ�2E����'�f�S���݊h��/ޒ�-��q�f��\��_gO��K�\`��m��`���%z��o����Z	\�M�g@o�u�aտ�_d�,�Q�%����9�'؊B���v�m_��̸ 8�ĭOʩ��e]���BY�oSD�/�Az[�S�m ��0���Ǵ��3G��'�qqx�P��@"���f�� �+�P�l�z]^ƗvP����"��Z�ʢ���A��\�"��g��S r�R�L�d�f���L�XD4�g���?�f�+W�ݿ�Fc��8cG����h�D���R�?��=ڧ7*o�D��8�9bh9�6Us TU�p3O�.K.i��Frlzp�!��<얌���J�%Z9*����5��QC��Ӈì���p�c�>�4�
?������0�qM��KL��{Ah�͜?��֗�}| [E飯Dq��',e� ъI�R�b�"r� ���7�o�����0^�0]_���	:V�}wA��koZt���}�ʕ4~,_���*�����s���J`�w�C��I����;>��n��Ԏ>���QHdu)��@j~��H�+� ��tv͚w����9Xz���w��f�M=Am���40*��$�]�X5��h>�q5ĩ,D^�؃����`P������}��!u['8�B���w�q�h�>U,UZ�:�Y��?H��#_+!��;�|V���y3(�Ѐ`1�(T�8[�pR���j��t���-�kN����vH��<tW��6g�̡�=���b	~�s�4`*�S&T���*��ynI7M�(l��DM\ץI����"�ud�&`��Shal�j#����ػ���`NL�s�)���q] �;�ݖ��1+�c��#A��r�$�n[f�4�����j׺#��y}�Cwڛ9���.K����mC����S�ыZM��p����)X�K�n��%C2M��Vߜ����܈V$���}d�D���>6}wnq��h�[�Mul_��:%�{�M�DV�~x4��h��
��� Sh�S��1V�b_��x��NJ>���4!2�^S�0�Io�KM>���V�O���=�NIA��;1��p�N~�^�>�b��IVR�!��nw�Ѵ^��2���;�?�Mϸ�u��%�i�qP�Xf!7T���k2��$}	�Ū��ְ������Bfb<:�'����N���q��� G*�A-2��@vG'�6C9gU��-c�p�(��lq	�,�+�dP��i��<��Q�,A�R	�qI�,�3���Y[q�fq<���*�bJ�#��}�Iu����'���'3�R��n�^��`�-�.��۽���$��+`��׬&[�Q���B�����G�
]��L�[U�L�9IY}�=ӥ�	�}������i}�p|Xg|}C^�����?~�;�3-������q8R$}�gQ�]Ŗ�6$ʈ�r8�x�qU�}�ܪ������Ny�:����c��+�� 0���F���ϥS�H~���i����N�V�Դ|���Cڹ����a��3i�2V�q����ߥr�����J���� {�4!XDp����
����롄Z�ޤV�;�y�-{GGܜ�Ӗn�O�B$��
��� �ݺ ,M��Q�͔�A�5�`�R�������3%J�3��M\���=�"�O�m���[�|�7�UΫ`	2z�r,^86��>��jV��G�>��(�?K j��=��ⱄL�9*�)۴��^z }vk��kC�Q|�#��e`K�i�{F0�P�S��D��$��Ua���%9p#Q�ULR�5sҥL��.)����֍Q_�*9�:v��~�����&��i��B�xy&XJ�q[��3T1eS6��fZ�����W�TiG'pĮ�'SAm�`����e����F_;+>�fh�@�\���R8yÏ1�H6�YjP߆bC��#�3tĀ^h!K�X��.�#�?ވ��珑�m=�̳o7�)������>Z�0�{<M'���UL긴}=�uj�(ſv��u�#7ô��%�~@P�5��U+cƯͳ�����.�̛�����\J-x�뗩��Lfgz\GC�s7hż�s�q�����O�T���f˰t�����z7$Oq�h�dOR|oA�r~8CY2e5�� ��ɂ�5Y�����iS��)�w�*<('�i�m��1F2�DBI�W[�rt+�dՆ�\�_�����3��������l�D.�Nۨ���f���}��mR�����tH�p�ې�u�dGڧ�����18n����6&f�`/�LqS�`�j��;��q����(����/%K�ܷ������s?��et�C(ԎѮ[����N$��N :}x�"Cl��J�j��l�&{��B�c�9�_������8����~�$y����.�/���|�;�O������X��� ���&�v��(��X�Adnؠ!�)��E��'�>5oEsW��O�K��3��n��ߓ�ފZi���e��#���.s[��
����[�5A�w�c`͡C��v�䉢����۠2��n���J�x���#�����.�yx1f3km�Rk��RK��}6�x�Ts:�t��<1�9��o�g��E#��r�n�J{���+HU���l�,AXZt�c8e�NӬ|�ބ��pW�Z$�YCy�Z��\��:���N!������ƚ5�>T�|a�-{	�a�>.�|��G�.Xf��gm�{���7��q�֌�DG}z]u�j)eտT���̨@ѓ�y�$���#�A������(��jֶ�v�F|䱡��U�5�z�6
W�]����_7|�0��`{�TV1 ���B�+�0��	�����	ct^�K�� ��:��능"%,�h�i���<D�Еx��	L9�ej�����!������Y���@������7�h~ }L�Tv�g�v����jQ�P8�6���p�j�lѲ�	�5�/Ў�H������Գ�p_�$�#�s��7��/g�ZBIdc�E�MB�xE�l?�]��e�V��0p��z() �:ʑ@,>%�f�+E EB���%#o>�� L }�w9w�����!���Ě#�6ř��M�m�>�+3F�f����҇p���5���叐��LGӾq�F����}��A�i��9���{�r��C���d�;E��Ofh�kkA��l�ł��Uj�=F��h.�+���?��)E�t�$�*	G�A
�_R��"��+��4�*^8�H�i���{����'E=`1�mB�U��uȤ��qİb��/�2jl�"�v������^�w��0q��g��ązMq��x�1��*�  
��Z�ķ�I!�+1µ��;��_�*�7ʡ�-��=/`��"�-0t�/�k军�)�D/k�#jE�d� I9_x,���M�˦JɌ�����P >Q���㷡h�eu�7���P]S�t}���?�?��o��}t,�D��
�x��Q(�Y�<���eh�n� R����^�\�v5��+p��0��M�䄚;L ���QK*��"Mo0*�3�=%���R��M��Жm��qXop4�V����m�G��`�]��i�`K������ �=b*^�{�i����l�{���{CCq׭>5V��_r}ld�tWPb���?�ѣ"��x!�R�/�Z
�6�^@G5���pS��cP���;8ۋ&��2/uHik<��<����dQ ƣ5#gL�Ob
������.��=��;R����rh�����Y(Y�Y���j�dSy����ɗ��0w�ߧE���M�qn��Lw�I(E���O��Z%��*h\�AZ��G�k��*v!m�:�a��̖�#̷���8����i
�9a�|FB��h���U �dzSQ&-�BD��8?�V�P��V�w��^{���5!ف�����7T�7���Q9�K��,) � �SM�����(��̍_<9�g��[� �Uq�Os!G�9o��W�ߒ�B����Y����8rf#�7�R6He�{�u��<�q�����rvؓ*+/?D$R��.e���8���E����.�ق<�_��*f>�Ȉ��g�r�S�ړ��o���e���)o�DG�,5�/:����U�7����%�@�f3�0������LR\�.��RuC棯��YB�p��9L�TT���pt�z�Pf_��v�fЉz̖\�}�D����\���,����\Z�[#W]�JD�S��J�t��q�`���7��s*�2�q1>�	(��jkI�8���H�`(��-���UOܔj���˘��P9��!^��'�:H��_��"���x�7a�,��̀����#�=�M>u`�Ԣ�SCT/Đ+{�rFt�>ߨg-�XՅ䝊;��>�hj����e�n��ak�F���I�P���'�p�)5�O�w4jG`I��kK��g���i�ظ,<�>������ �fM{
�<�v�M����y?�!�g %�W��q�DH��t��p"#\��#�4�r���B\�����L��Eo�~Pv9�����c�v�.��\!K^f�H0d��#*��}��BQlW�2_�-��Pj�C������������$8���[����) ����o2�{�TPI�}�&s=���*T�h/[䂉3%�eL��9�� ��N��:eM�D�.pό�q�Ӓ'I�ے`�D�jm�H$ �Ih�=�T�*�������#��5G
�`u�����?6g�qA���SRr�}ea}Gt���=���P��(��5��c�!�_��?h����?\�m>�ӣ���d��%���M쌾8-?��%�al�,�I-��ݤ�⁂zLF|$��J����eD�܏���O��A��<��D�V�wѬ��Z�%�mA�+U)<_Z��W�䍪�D~q^���M���=d����y�	�aN�<��=x)��,"�=ܒ�3��}~�]�QX\T��%�}u�/���m�PxY'���܊|�lu���,���������ы=��I�m=�r�aE;�i�!��Ǎ���v/I������~�mu��T4Wrv&�nq��%�|r�ys3�G��j'����˞`F�� �R�PђY���ay6<��ihJj@�f�#��������t:<�A������>�C�����C1�qaY��P��d��%���D3Y�8<��z�0�Й0�S�o2v��HH+�&H�|9ӫ?X\bt�Q.��a{E��"Y������+��
��I|hW���v��������&��lcoY}v\����e����+��$���"��*��{�N"���7�)���fR)C���j 1Fh�$d��@��ON���ʅ��t��޻��1Ky��:���Ԉ��+,�o��&
>.�ɣC��I�md��/1l��)���j�OVu��[K�2 bv�\���Z�^�V��j�L�p1T4/޸͟2�2��e��/����v�eOX����7�/��#�6��tb^�#��]�<��gR|j~P�R�+����&я�-�$��d18�cR�Y,D�"u��Y�ȤPQuW���6�5�!^�%�
v�3�K��ψ�9��X~3^�}q9�}¹���$³&����ِ/GQ�:<w����u}�&�##v��H������]ӛ�.���-i�[�A�S�|�e�0�/�V�nZ����W��=Vne�v������ J\�E��D�͘!��ٰU��3�HJk�0mF�y��ĭMN��U��+��0��-�'\�RZǿ�o��!�T(��c�$toA���I�,@ce�6�0ox�ݰl�����C���{<t��3=,KWu���=V:��*�-����}�b2�q�\�9�$�l���@��Oe�^�u��g=C�z�m���JPq�{ ��!�;l���z��6��Ҡ�*L�|���~��*ٿ`Ʌy���
mc�W����Z3$��Scrе�
����2�`�����Qoo��)K�& �s��ܑ���[�Sr�O��
,�� ��h��T(}�U��=�/wS8�02�`��r��00���+��(|���/ŵ?YG�.�G��3�F�G�r(MW.�r'�ީĶdXT�A8�#��#��^y����͎�×H<��á'�4�<�ܘ���u��5���,-̛_t�{ak8��2��S���)E{S l��$��M�"kV�p5w~�\p*{J0-�\�Z����St�Im�C�T[tkL��/�¹ƥk����Ey�*E�ꙹT�ǖ����M��;H^#33��Q�_m��'X�$�*���﹆6�����"RF�����Y��0"��ۆ!��l/�0��#��%X���P�Bj���R��̞6��!%<f<��si��_�OԲWA+qr�]t�5	�m�R�ʹ�4U���2����Wꕴ-(��3��\��n��b&Q狉�{<!��˃�1�:�:T:�r[�c��Y�r}�i��zv�7a�����yV��oBqZ��6����.�*��x|P�v�8�cs	��O��#CZ�TyP�>��z�HJ����D�h����F'�e<q*^]$ ��{�O�[]0<w��U~o�D�a�#]_�ʖ��Ϛ:�Y�vgs�����)Ǟ��B�:s{u��fd~'���$�Fh�B���<倚�(�0A�"K��b5�v��G PڪX{G8N;�o��P<�֙B�uR������ 	��&NΨ��瀄��ڔ;|�5ށy�{�9��ܹ�]�`
�٪��r��^*d�a��̇k�q\d8{�hq&\�<��R�r"ęd
�t��{�!����&$ �N��8�]��Y�� TVH>���i8O��H6�B��wc�I���7��Y��L=�u�xy�a62QhR���(E������DE�{����W*2"�S�u�cn3,\q͇��(I��U�.="��7�E��N��	���
.�gW:��ڬ��n��v޾)��#dۤ�ˣ�c(���`�_�
w&T��5&��.&����kѷ����-(6����t ��^3�R�Yʢ��0���Јa-P����~P'5���M�-�������d=;���YA{Y}��S���x�}��=g�(�A�ة進�׀��ѭ�C�l#�p1�bJC�"LZ=��j� y��#��R��KE�fP�DRG�yK��-�*}gmG�IB�t�̯;)S'R�Bt��8��û���/��h$r��� ����AQ6�x��VM�x�%���/kge�#�Y|%�:^�˻xa����eC�BJ�"�R��B�D��uZ�+���(԰��]8j�2��8I�s��5;�\�W*���gg�oa¤5�O\H8� �лp3��]0�2��kd��Vp�br�����:����t��=��%w���f�MF}��)x}o�Oa�I�a<������ G�p4ˡK�t�����d�xfH���ޣLt��Q�-�7�w�6l�X���5k0���7��?��Nk�q��n\��xk�^TZ�g�}��!�2����T��6��6`?�'u�v��#@a�?�WI���؟�-gn�80����_{_�L*�ج�}H�T$u)���-�L	-�����82�V��EU�N�_0 �z�)�\^JY
��!��ߟ���ـx����1d�am)����L��M3��j��$�����y�T��[7��VO��~���'!�N�J�ֻ����\�|�ؕ[g�$l�H�!W�� �
�B7}����!���Z��5gLu9	e�䨈�`[��!0��#2{���f�F&�bTޘR��()�X&CW��2k�n�b��������_���H��Ȯ�x��9���/�f�7�)GQ�-�?��TW��q1��y��~�1�mg�{��:[n��'2S��!X��"�K��^,��5Ϸ� ��YWmJ�2p�V~��k1������ҏ�M�����9����s�
�2^mu�=�����oN��s3i�0aK=A�t�dĶ���㦗��tf�N�� /`�U�^N2��K�Y�0q݋��1�v��q�ˈ�����sۦ�ɭ�G{��CV5K��u�Ko6 ��� ;��ŭ!����D�y�oLa�w�?Ɣ�.Wm�m�s
��ج�C����1H�}g�����w��P����-�==
�NKEҡW��H	��c�C^ r�'�vF���U�����o��I���/^�>p�/&M�Y(�Q���tF��;G�u�ɰ�j*H��O;�wY���`#�j���~�3�Im�M�T�����o�pj��
϶�*>C��1,Y	��ul�:���%�#|���s��ϣ6���O���S8�hJ�Ʒ	x�������)|��D�^��0��4�p�nvL�ߟ�ʞ�� ��l�xF��$6�6c�e��Ǻ�ubtc�S]\�Ь��/ �%����8����ˆ<���5���d���*�u �syBZ"�!�:sv�����k����ʏSK���SB���2�^8]VЎ>��q���F��ա��}��^�0.��_��n ��u�F�N4�Nʥ����ݷ�,:^覫	�9�%)�eA�B"D���>
�k�6~���'�¤d�3�_^��N���m7�a��+�^BM�Y`�0^�J[M�r�(���~���yt�Z_i��q�=S���5U� �/:̓��;�V�&t�ۯ6@��P�����N� �'�XW*�a�uB��D+��H�����UW�뤉���M��S�I�%���hۘ��}�`�U��NL�>.e�j5 $����;cȪ �c�����(����p�W����ýmU���� �d؊��_�/����>w��;��ǃ�3�T��*�s ���%�x6�yV�F.���k�C�
�i�ݍ�aswSs]�F?���e^η	q9��2p�0��>5�B��2$�VaH:L en�D��K��Z��%��מ5!�Z˃P��{p�h��2�4	bӴ�ܘ�����s6_@(����Lrm��%K�LPLJ�tF�&�
���ƍh}`�Ol���s'v�"���{`/��K��Y:�ǿ|�(!�g���.RuX�fJ�w�r.�Q�66{�RO��Bwl�$��'��0��6��� ����L>Ĳ=6LZF��G�	aq�|?8���Ƨd|뜖A� �%���˳��^ُ��&Xj����^"��0��2�k,0y���tZ����Y�w��p���EDt�����Tw��weEV��۾��vs!�}Hd�x�ֽ�ӕ[gG��p+ ������5�cr�T��4GL�<�F#
�=�'��?ޮ�jP'��p+h�En�A���ٴ��Y���g�۔"GF�c����~���P+�����^�|���0Վ1'Lc.]>��\�b�p��VAI�c^� �|�>��E���;�a�`�?a��ߖy�1���D�vzR������4�@��G��n}4�_���'.(!\������pw����s:�%��0R	��}�@1B��Geo���j#���+3�%�Gl��.'�.$�I-"�p��¨`1�-7�	�_	��-��v�t���&O6�F~���o	��b�^=�O&i{� � *��=o �' �FӀ��[�'n�\��p����� ��Q�l�����d��ٙ�_#[��ڝ�0���Ak�+Ae=���=˰H��_$�1x������"~1��v`��:��4"'KV�P^�ȓ��EM�+�Bt�����՛��m|4zZ+���8z�z����m|	^5c�P�4�9��P`���i��v��Oć@47bolpO�p�7�jFPR���Q���u�
N���կm+QOq��=�����N�z���^7'#�i
pkh�iW~
���Ss�j}�y2��0����
��6����t�Հ`������/�Pc��V�IQ���(R���
�v�ё�Pن�j>���?#S��m
h��|6œ/�P>���?6b���O�NOۄqQ��,��*^dX��i�[��kJNGn�O��eu\6��=&y�v������z��
�û�l����8U8i��_<����f���hwE�^$5��u��U�YѺ�����F��n��!�5Gח�J�9�9
��#�g��o��h��3���K���8�${U�i�a^>�o]�X>_�n��1fϪ(�
��5w)�W�T=�O:(/���`�a�xϰ��>Tgiʡ��"2��J��>�VC1	���)Ut%�<T{�ۜ�%ӠT����F���hE���t=���Aqz�6r�#���h��
�Ԛ?�
���f��Ea�_����@m��X'�6�H|��qOE�p�������oʘ�S�K�[iL�	 �9 �y���M�7ˉ0���}U>M{$��R�d��bV����+�e8){��w����\d�X�dvW���'��	@��C���-�j?�/�(�F���LZi�HQ����!�㕑�P��I���M���qx��^ ��٪8���؁�ySD��cd�a�0d@�Q�E1xO�s귀���R���D�8��6E�l��9>י��9L@�V�{"�r��4�=�����X�EG���p5n�8c-6������/�y� "1	@�JE9Op`�J�.CIH��d<j%w�������~nE�ژ�_?�C�}G}���?�5�ɬT��λ����	-��P��t��Lu�pۯ/muɅ�[JCVו�S�y���C�3�_���c J8��n]|�L*��f;k�/�����;��%�e(��U����aQ0˖A��9��f��#�hx��{g6D�"��� ºo����+4���,O�)��G�Jxz8((عX�8�S�PQ�¹-/^"�Ydȍ���H�}M�BM8c�V����<zO��s�&�N�I�1R�ջ/�C5Y:�LA�y�ڡ�SXX�KL���x��C��h6C�W�f�#⯉_-���R/"���	8m�b��i�� ���[�nMFZzU�>�;�|��9���Y|W|����� Q�2*:0��6.��MN/t�z�N�t/%g��i�¾8˥˟_x ڒ�.g;=�U���	ʌ������,�����'*��j��D��C�Z�q�g��a�Ky�.�+t�A?$hů�/٭�Z6b9a�{������X��m c�[�b+cM7���nYo4���K�����X��y*�i/R�2^H��Ӡ�#�.U�0�#J�?�����o��g�?<�����ʽ׼r���@���^E�V����f��1x��F���{`��lneF�����``�L8-������1Y��.�HՇh���H�����+�L���n��5s��{��]¸с�8%��-���-�H`)^�nз�����˾�ZN�s��5Z�]�GS�݁��(��1���>Â�{�э],$�=U������en�5��A5�Y�a���<�yc�~��h5�l݀�S=Iny'm�;�!���j���F`�Z�5���1���iFxQ�&I���=7p�I����k��n��R�	p�Wy����Ź��p�C���!�mB**��֬4�K����Վ��[�Yl�3�4v�M�����`�ղ��^��śи��"�>Ak��z�w�/��R}I�׏�/C��t U$/�D�oe� L�\^�Z�iI�aC{�t��b�ްnf4�.*�'*)�/#/z��Ǜ��)f��̻/�+/�W��+�;�Ŕ194�B2k�%)������j>.R��$�b�
L�ǻA�����YNW�3��K��h��6���Qy�������K�e�1q�*����oIE>�[v��h������Y&o,UNg�N���8�`2�_XF��k��2���W��牗=sYb�12���'�j�ERϊ+���Ti�q��JQ��?>Bh��l���&���;d��${k���(�FZ.�n��~� �{�,M��TP�����~�� h�Ю�ЉHUj'�`�%�1M�}z�����m_��!�v7�,1��(����g&$3�l���0���m����S��A�b���Ͽo�t�O�1��Ť3����>gdyNk5K|�bzx��-X�N�=��`��4W�G��~u��M����LӁ�j��KgPWYվ�`OW;�_}��=���=e��>k��8��SL��,��6���9�h	��YgM��{^'���G�޵H�$��
����;Qޝ{�;�-�ԭ�w3�g�I�lڮ�-�}�P���W� �2�֧�YbJ��i����F�6�4��k�e{�̣#bIL%,��E�������,Ȍ-��B�R�ϖxi0W2�#�RcV���$�$�����,j�,#ᐑM�L�w����$��������vް=S
�vV���ϧW��Wպgc�7���N�Z�������?=NCm5 	:�|�vݟMXX����yCŅ�W��4����(c3ӦȐ��UO�
.��ͻ�9���=�"�4Z]86��f����K2��ոo�RȄ����r���4W�"E70�Yf��q#i�CɭqC��\��ژ�Ē=*���Q|�IyH�+����]���<5��0�)�����W������`�󺪩��S��mH��Ō�QB2��9H�NZ��8�'���^�br�s�e�o�<}*���=�5�a��E�sY���
���d*L��q����r8������Q�^M�G�}t�i�vǵ���Ƹ^U��>U��F���m-*��jz~`]���ɔV�K����� �������چ�\�!a��Y��0XJ����u����7�pR�`��ǚ��]2^��E��:�Y%�m�X��(d���HBe�^^�g���>r����9�Q>ݶ�!�W�
��G<�`���؏����b#�69-�|￘I�<�Πܘ�?�����l0%��M���]�S#�����,tKiK,D���G�\Ǔ�-�CY���+6��Xj�jsC��*�2�>��b���R��ۇj��˚�uKe�t�gf-J��Wg�v�g]]�Z%�M7�2� �U�-��2^Ϳ�N��y�8����M\S��Ey��AZ�ᘚ��l���}��@�#V�y2^��r(�C��A,�gFġ諧��_�ŊO۱2����Gɦ�r&F&�w]C��rn{q���۟J���W8K��`��c�\�����Z�n�҉��pٗ�(@.Jy�����@8�E��#�A�L��Ҡ)�/�6Q��+��%�.���j0. 0�Y��C��D�_6U�O-�������z�Y��ٷ����<�I��ϗ �O���3��[Sy]�E��h�����
�1�i��^�N�&�e+��x�7� �B���l8�
*yHE��7����d,�Z�4��r�gF��R��x7?f"ր������? ��Z7�I����%́V�:����^�z�yE�!�1�l�7�=d�!�=dNIJx~ЌY������fdZ���2��.�d7Ѧ�V�����u���Aq���}5��z���_�ʼVpLC[! �#/X���|�X�*ev�A��X ��}M]���-[��zd$|��	�@JZ�]F.*�n�{�@V�=OO��O^4�U���!Ƭe��M�]<YE�7�.��$��W�T�b���8jbeHq���h~�R��������?�ݔ�N�C�#�.��#��>���|��`���5�c�(?{�q�ֵ@��U=b��;a�7K֢������ ��2��ȕ�,8ʜ�ꋍ����kX!�e�: GXK4�1����T��F�E��E}�!���`:B��>�!����a.�ҥiNʹ��!CvmV5�ʯ�ȑT��?'���Y���ݻ;$�sӅz�n]�|�i)���>��]
��3%�ԩF����?/z�=������pK�v譫� ��]�s��{w���|�W�v1��\ܘ_�vc��a�p4/��a����׾m�7In����%�EJv�-;ıkQM�e(�ڸ���W	�$ΰ��w<Z:`��f4���h�����2؅�8`J����&��0�\�~��ǲ�#�F�������_�ďiu��`���$p�%�xy헓��1��@*nV�8�t4�L��ǚ��Q��Pw)��~����B���3-���Y��j�d�Ps||%L�|,i��-&n��&����^�F �O��dB���G=�5�쬸��4O���类ױOe�Pȥ����,��jy�cכ_��\��"j�z����������X�V���ψҪ����Й�.W	������z����܂v<_�>����-�R�X)��jG�MK��m8Z*� ��;��!�!ԅ ��T�u�D"�ELg��$�[bc����3��jق0X-x����b����3A�#̚����˰�M��r����
9E�o�6��V_D��v%˧���'��^�k�t�.����*e�>���+����Ib��化u�)�"�ʨ��c~g����#�]P?T7�-�Sn�g9d���æs.��)4��hv'�H�%��m�Eu�z*�O����-K��L^n�+_#jA���W2>UM���vpy��?�{�9�v�&�ş��ClP/�h�b�Ľ�]������	`�fN>!O��˒�v$�����ݓzO<��ғ����e��C�&��
��Ζ�^�L�0��7�ٿT���#7�}�e�B�lQZ�0��sieN�\����T��Q䘯 j�%�P#���pe�6y���$�����5dFMZ��p�U�C�9�2���Uy���<[��a�	oB�~�R�.��f�Y��K���
I�KS��LY�����'='����[:xqu%�Oޒ�	��r� �|��Z�vN�
��6�ƖǺ��ѼE���_��M�pM����=m)��+���=��\���r_p"���4Ћ���!�4N7}F��"�@�.�����MaL��k��f�TS��*n�����<�W�lsK�G�;��~w�6~��<��lh :����瑒)�w����v}U�ʮ�P?����ΡrniL���ΞJ(�"�33PP������Fүl%R�,vm���#%�o�6|�opd"a����:��E�<a�����$[w1JY���Ar+z4��.P5���{���.w�ru�G$4\�m�VI@�yMc
ϭ�l2PA����1o�Lpl�Ԓ4|ѼK<�>�@��P���_��>-�U�D-����lD'�1��;F��
#V�Ҩ�Ӡ����Z����1n�Ka��SQm`�ϖ���eĈ'�xÕ�i�9��Q!R#)��	~�i����ҙ�a�z^پ,��#*��@٭✍����Hvq�|���xY�"͎��B� �-��am��:��U�DH��4��%�f��8��lv�V� 6S�����mQ޴G7���Z�����UoZ/0����^��~Ӈ�6��u�ehrŨ>d)��(^\����&�݌���я���&�V���i2�1�JI-7�]�K��+]Ҝ^� ���γ%�����D@D.�h�6���]��^U-f�T�Y5�N�q&r�r�ť��S)�2I��W���V-'��m\O K��"��<�g.l ��%�t]�0lպ��ho�J)/#k��w�2T�?%�������:�W���>�74�	<�R�׻\�7f�3 �;��F�_]���_4���41�֞n�;��7w	9�7\�NL�Uۤ�e����o�_тש����&\��.B��l�<M�bV��vo�S�,.���,��Dicʔ�Z�ᚬ�"��K�qA�T����, ~~-&(�QZ�$����w���j{�kH'��JP�7Έ�Q���Eģ�	�r)�Q�]�5��0Ъ��>�Av�}��]2�?Il�3�IJ����5�`�r],����k���c��0ƻ�5#�)�~��Ǔ�,���tw�I�^<P�w4�,�9jgY��F�E���I��qUTݥX\��r�[�D�ð�wS6
)�R���Q�����D�n4�2�v�R�wQS�P^���d5�q��V{�2��q<�pE�u]y4�ھ��>����H�ܚ`B)=��}Q��I¯*��,p�-�V��)7���	�+��WF��^b���?�����ٜ+i�"�)'��a]��*���8@����O�܇�U���(�%3�����G1��G)�~��_!�:�r�L���D��k�xk��:J�wPB8�s������N0�T)�;���%-�o�o@�/�~
:����S7��� �#4�_u���"c�>�ӂ������+"�^��G�anB#e��**���-��O�ǫ5?Az*��o)n��D�v#ϧ�N��n�%U��0�@!�=��гWн�;��I3U�H�ѺW��Q����# "	�(D�U�7��71^���j�3�2�L5.Lg��т���0�=���V��y_g7,�E��g���o~��I�X!�hv�)��F��dGD����𪪈�Wq��,��o��d��ǂ_�#��a�������S�����y�cxRieD�H_����2�� ����jݡ�
zE��)_3��=�C?g�rH�Q�j�5�#�B���'�bl6���U�`�����=&#i�s@���|���5���)�)G��A��03{���q�a�.>��b�\Lji�S�F��3G��`�%�3����Q��/�L�%��晴� 	��3�x���kU�Yg��1�{ǩ�-w�8�g��)&�L��b�Ƈ[\������,���vX���<5��sY�1˺ax���5�+bo���['��the����B�oZtz�����C6�rն�W{�<�2B����,p��<[�� I@�}x�ʷ�l�j�.��)���B���NlτKu-�8KC�S���˯�V���|;e05M�-��6A�W� �3��{G?<lh!���)��F���wZ��y!}T�c��^�=��0V4�Rjs*�i����[1R�yl|��{E
'q�%�zb+nV�08{Y����: ��E)H��g(���),���ؿx�ܶw�HQ@y�Xd_ƥ��.�쯮��ˁ#9��X�\�_��/p��Q�<Ӧs4Z�bn:�Q7��3�H��+|��s�"m��e�9�Ў��잔�f�@"�'�	4h͊^ׇ[J��� s��jՍ���6Z�f'T���tw����Ŭ��բ&{��d�`I�7>TN�3�)ʚ'n|�eg��&|Kz��؋�6�g��"IFX����:�"�,�(�%��V�1򖪙:�f�d���Fe����w<�{����$h�MZ��D]Zp��t|�:�gf�����}$��"up3�+�:g$6�^�R(��� �}�)�F��ӵ�����_��� �aW?(�}�1]֠X$~7IY5��u2�>��V����tB�`�utq�f}#%Pߧ<L	��)l�	���RU�O���f_&��o� p�_���Sr+
�K�����m��?�E'����#Z"�
�P�B�(0���{؞��@ŇFؼ��<k=�а������Pw}�)�����������6�=$�d ��zb�� t�VbBX`;���H�ܖ�bNE۪��} �[;%^�M~�-Z5�I�3�<�ô��"�SK�yM�>>�1����M�9�L.Y/]�����Fᓪ����{z����1���_���Gh|����<� ģ쐨;��y��!�t�ʝX�F.�|`zqX�p�=�F��:� 	]!�q��n�����T��<�?]l��^���j��.ß�+�1�Z$��\��֓�����y���CH��	�v��΁�c$)��x%T�}г�D]�(�e��<�3|+*ğ��������0B+�Sc�A����@e\jO b3���2()79'W�ËMf��値_/0u���U�Ϲ�1X�ػ8a�������	,Z�_�[6߿�ƫ�o�m�Y���A�b�.�s���ܬI�~�'�'i��CEii k�L��i`�qzDCj�8um�E��G���Y:[�:X�R1�@�E~���QPw�`
�pQxrX�g�-�4�a"�y
��
��Ʋ��93_|�8j���]�r������ׯZJ�)b)B��%���*�o���5��Y����KD�:6EhF44��rVm"Xv�)+(�a���C����t�E�cQh�6�1[Ҋ�m�U������B?٘l��%�T�u�P5S%���Bf[��I�mw��S)/���Ay�L���A�7"��yRS�Z�~�B�o���0Ĩ$wʲ9c�˫+G����߼tV��ZI�~Y )$2�[�o���	�d>[*�c����X_���Ǆϼ��֚g�H ��s��"���i�=bv?�eX���z�eZP�]�k�sV�3q˲�BǋV��K��nr�3Y5�q��%�**<V8��� ^�$5��E����V�8�p����x�	7�ǹ���J̭�,mC`�RRĀ�Pu�7Sh� |���WEɛ�c�3���� !�������d�"ӑ��~�᭎Z�߻0��Bn��u�5���GفqHO_�����qKY\r���+�&�)�9�l����r�Iog�j�{V%>Y��t�H����u:��ڊ�7����b�k�lA1�X�.i?d��-���;20���C���k�Ȱi��{_u�'�7f_�n��:�H�,����1������t��xx91��ݡ&G���	���e$����]�s~*	�"�V�i��'���?�ё�2��Q����&�`N�<2F����ы��Ъ����t�#��+�I��@*��V���"w�"'�-�٣-���W��t>f���A�H���#�� �2����^�S�sp?�2a6@:liEvzS�f���q��|�+�A^o�Ќ��y�� 	���ϭn\N�8�Ӈ�.Q�t�І�_��L���RU�:���(��v�P{A!z�)r��M����\�A>+�x��|o�?��ޥ��Vm[�?��7�������sg���Q�1,�7�m�	�Ƨ5����D~�k����!��:�i'V-��U
o��"�A�{l+��wk�1�Y���,��Q�D��x�� �{]�_�W;33%���J��}�����Zs𫭍Ö6*����{���V�>�K��i��iQ��y���qҨ�M.>����41�,Z:�L���BDA���_�d��^:�م�Su�0�{�$��\��RtY�0r���"��6g~�$9kä�&q�y���D2p� 7~��lDϩ�>��{�\�6����=�㏿g��;�#�^S8���S�c�%��
@g�'}D�^2�7�@ :c�g60wa��n�H�e?�4�2D�#�a�Y�#l�76��� ���/�k�N����~)�j5���'߸��h�?	��D���٢����$�U�5Y�q��%����	Q8g��0� F0&���Mޖ��y\@J���S���+�dALd'�+�W��K�6�OWul*�|?7�s�
Ɔ�T��/I�uP�+���x޻�z9���}����'Uʼ�7��!�����O���i}I\�iX�>��>fX="tg�[]�hw
��1(ȅ�j��%�[���2���'E0c�!D�kR�r����������)˻���91c����&7%Wl6M� ����3����Q�sb�K(�PP�����=&%���u������T��[wݢc�J��J�
��p���Y��·��[`ԁ�41!Ή�� 
"������*��għ� ���'p���\�K�p�Q��3��GM��a��U������U����fQ<mŌ�Q>��p't�X��Ri)�S�+w�&<K%���L]���;�ΆhD��eWT�p#�x��e �,�q+O��]K$Ս���-�FC(Eƚ��FZ���劇ԿDH���Τ��*n�~^���I�2���H��WoS���ӥ�����,����O��J�/�U��#�(|&�?#�+���{�m�Y�=uU�b��ԝ�ÈE����ZMʥ��FzK.�wS9��0p�"^������G�%kȷK�Lźg��/�H^���V��Ȼgn%���,|��ⵂe ���+�ST��)|H���zq!4��r��h}n��!H7�.�7?<#L�x��Fw���N򏮉P���H��j��[LT���G�H��W�rY�{����Y�7��O��I"�$ ��D��eJ���w-�߯E1�X0���h�����$j�mz�aC�f�e��2���\���!v�|VF�Bo�N$E��b���a���(�]�p�39�E�w�R������(@���ɼV-8�0�?}��d'n�"�B��F]������qۀ�! ��F2�	��:=�6ӿ��oB]������ɞ�IO���\V|(0r��EȾ����K@�֌糰IUk ��L���J(��YU,��0��&�(2׫/���L߲�F �� ��Az<eȸ����Z�A��s�gx)�ζ�Di�a]�5�Z'���30��<�Zꪙ�d��Ou��+_����i����N*�Mዶ�������s^�ؠ��8�t2[K(}���"d�o7�� �]�Ҙ��F[��ŊZ����󷜻j����i:��[���W�	�d�,�&�"�s"�°j=n�z��gG/gDuX��'���(����F+���"9����0�7�j������xI���h���+�?�4E#:c~90��;����^h	z��z��"�Bd��>'���C�+4�g@����{8�����#CI3�����Q�0�O����Є쬥����g��H�p�;��N'-��)�j���%���~�����%Z���ov]oKy7��ѡQD9\Zk���ǂ����_���g'�	K�q�G�x8Z���uQ���mRO�TYIXv-�a�d%�(J�����keh=��Z�������'���o��2+Wٽ�0!�]�ʲz��~����L�W�-�2g"�\Gt	B�D*YQ�^��yA�~��YD^�.���z3��9�S��w7>|�!(,��:��U��
�jJ'��mܬ�HZ��U_ �c�#��q>�m�IH
^���؁�4�3��eHS�p�ƣ��G�q2�΢)��A�0M*�l/�oG#��^歗|P6��k��xl�`7vj�/�O���b�In���;�
S��F��o�j���4vM�	2�p�<���{��P�Ǫ0�� �M�bؚg�%��Z��6�V8juc�	��I��<�b9��Zt8)���LS���I���OM���+:�ǘ�0�E?�ie��>,ƍ�)k�=��{jǏ%m�t<G��U��	W�td��j^���>���Y���h<�z�� "�{ �� �-�W�m]47+RvkeN��sF����=eJ�F05�@�5���8�������OOf�5)��'^����#�}��!��X�x�ٹl�n��j))y��N�~}��-tQ��J}����ƇY~:C��
a쩺�>�~��p�T$��T�=��I�8`ys���w�4��I�F�#���,+U���;��Cۏe ӊ���OU�w���e /o�(����)C�S��oɽq~�P�j�A��5��\-��h��?Ő�~�y�0�Ǌ�#�6��G�,�a����1pT�4���.�;�*n$Q�_��R��71L���q;j�[�/�xO�&�#)>�a��y����:'�dKԫW>Ȇ)e���x��D���Xs* ��%}؅�1�=�٤�������D�NB^�ƍ����3츅X���֓D�u��a����;=BE��ȴMZ��q.�	k�$#���r�!l�H~%y�[=T���u�;�v'-�iN;f�,�w�I�Ğ�B��&�?^�Ң�A�s�n�@��k����zmc�?��F��.B���q{0�t%�D�uѝ���y.i�u���6�N��-Y���	J��;퀋�w��aA$��}#�W~�$ߋuie�l*�z��̴�E�Eկ!���؛����KO�-��is���0�a�Zt�^�
fsШf�AMQm��(�\��n?��뒑\lR�[�%b_���8Gc��7�x�S_v�Legh�3�mnaR[�X�%��El���=�A��m��:�v��sO6&!WC�T��w����mb�M�O��:"�x��R�[1E��q������M{Jv��<�)� ʒG/�x���y���Y�8�h����?�
$��
��"�>�UD�z��<U<_0[�cX�qv������~�P({�����z[Y�x���.�	������rX*�m��Wi�1��aOJ��%�~�"���;9E-��J��7ڍkc�����v���#y�J����{�g�"گ�y���p���KV�X�B'
mvF�-�ؕ�?;K�z�L����@��]3��I�a�T� �u�'�{�p��_��)��曰�-������l <�F����iv(Ք�H��~�"�{�k֎9�R��R!�1����*��
þY5����Q"�X	1e�x0[	���c�%�^VYO<G�Ic�w/؁#)|�'.���a@z��ir6�45 �a0
��0���;���9��.��z�Ӟ�k��-JX�%�/��n��w�)w�`���A�f� p�W�7�ܙU���yQ�c7������*�G}��>��/�ox�X�������O7ۛ9���&V��sߠ�,�(���dw��3�阌���[$4ї��"MG�K�Z��B�>o2�J���?*���N�D@��\���0�f��R7
Y؎:g���5!<Z�4������{��\�p��q	?�
L�^qYH�����t%�k�]�7��hSx����'ܙ�L�4k�C�eZ7`���u���.�pq�j��~���i3x�������د�E�v�����ظ���5wcAC�@!!yd�G椻F��S��\����� �a�{��<���.F�"��-��Ӛ�8D���%�0Ѻ�4UϐEV���Χ�m9��:Mޡ�%�k�d\W�o{�������^���������ٟk;�=�o	^"�/c�7�84z�Z��0�}f9��2�A��V8�x���	�y^QYd�'{[����ap�*��6s�n�멎E 9I���G�mFCR��p�ov�=h�υa������]{�e�n&	lOd�er��5~l{Ԃ��v~��J���g�n�S6��:�9�|�+���Ù���A��\IDbr��E��`�^�Pz&�����3��*R0�D�;�`e��<�b��6Ɉ�g�gwX7�?7癬;��PvJ���#?���c�Fy)���84�����W�Ғ���v�A[���&��,��qۢ3��*e<�}&��P�S�� �,"�N�)�d�)��e1By����ph6������~�}6�<ARkE�p�W�ɽ�n�c�GU���$���c8EH]G��wЛ���%��Oi��P3��2*)pE,�����y~��&�`��D���X*l��AM;TL�ǐ.�h�8���B�-�EI*�pŰ�YR���_E��~i�W��v�rH�/=���y��j.@��y�I��ȜZ��iV��p��y|d��Z�ͤ*�N	�>��U��?�V(	��G����>Y�T���{F.wff�v�s:YGaI����qc��l�M8`�cпs���\�IGX�)h����"����{w�p��Fq2M̶�K擝{c�
\�!�n�C�����jV�gmK�5G8��f�^�v�UW�v�M������`S���R1�=������=Xc�Ymƾ<��@� M�S�L�+�%W�ei�ۭs�dC���k�s�R2��uSj/�{1�,�,0�H�m8;�w�K�io�x���\��ƌ��6�$��+��6q>ywF�!# +	��e^�l��^�S/?.��DJ��AT�B&R�a��s������%R�_z�ұI�.˓�0`���A��q�uњ
�j�(��f���!�\D�m&/"�>��|��V�+&b�@�^�
�F�z�뽃=`����p�Y4���LUA)(�T[l�ݬ�ޏ���%.:V���H�^]AC;���5Su����o�,{(�9�U��K�vG;���N�o=���X�4��^�!R��c�{��S?�d,Sr��c$$��[���{!�C	�6)��9�Пҹg�L��F\��0?�&���~`��Y�Epct#� ڈW��0�u�	��QTb�k"���a�魈���GUc�ml٢�ƪy�N���2�J�d�g �QY�KSn~�g���$͗U}.m�ȑ���-��a��ӷ�2�Iy�ƴ*+HSz�!j�B�X��@�;ρ�8W�X-0�]iC+q�q�XH���-YgN:�1~���Ml��K������F�̕��GEKᐯ��ua����ݦy2�=9���㏷U�1~�,.֮����K�T��B^�o}Pt<'w����,83待k��+�����9�������	�c�-n� M<�Ǻ�B&q�Ƥ
�+/��p�󫹣�P���﴿��Dm%����w�o��p�,��ä�Y_5�ACҾ3x�8��{��!��P��2	C"m�9�㬬FѠ�]S�<EH��z�}
���q[�M�K� u�)}���"��@�&Y�H��`v����8NB������sqS�X����W�?�i��&��C4>#��7����Rze;�m��5�DL��}ފOw���??���D�b$��
�e)49ՀW¬�$����3~�J;�ʺYӂB�u�uf$B֫H�"ݥV�]��-��+3�a�s��~�����/F�aM#���ࡣg�B8�[t���YA�Vr����S��V-ޒ��@T8���[%	TQ�14/6NkR�f�(��4�{J�>��j�������tɌ�mQeh>���wzp�Ǻ_r�.gq���,!�O�p�T�j}:	kB���7x$���B	q�Vt�AH�G���R�kyj��� -9D��m��3F��zQ��	������A��qvP��\��=����$0H�����7Ǥ]3�ď����"��汎K&���_;����=�Sn���o�]�a��u-t���|����D�.���=����Rɿ*J��vddU��%݌�}� S~M�\^�	��l����/\��Т�`xj?�����E�ZI>+�A�uO ZV��ҿ����\�O��Oin�J/�Ln�<g�{��=�Qу�Dn�1��^�`�PA� ���2��s�"XlRz�Ӗ�\O�^e���!A��~n<%�g��/���5h^V����@QL��]�S^Y-���/@�*�����K�A�z/��䂣;ݙ/��
�x>uV_а�D�$g�W�(eɩ>&\	�j��?�����St�q�RA�Y�J�WLEv��u��5�W�u�E~^Q���M�'����	�Z��C�;�%���z/YY� �C����D2��G�&���L�M�R��]���3�bJŀI��P�b�G��QH|N�@����� �"�톖��:Lˍ3��_-@o衒��6���|>i5Fɍ�~��P����Ng�(`Jv��m�Sf$%��̳��>
��L��]�vi��B�:�K��PBT?"�3�RET��,�~b��ٰ��Ԯ�j��I���㈚O��N��gF���Ue�$<���I�p��ή���h����ID�b'`o���	���"q�!�Q����6K��i`Π���&,k�c���'�HI�,d�D@�`���l�]y�U���Ĕ�=���'�d����G�����Th;p+A��V_(�nyʧcYǆ�S��⁜��e�TB��I;�
*4�X�9�8�{N��Of;���&��p'�/�ҷD����fZ���o7V��#x������g���,�f<�� �e~�����%�:���(�3��5���G*�~!�����G�Q�,K�H1����B<���
ţN�"�_��u
: �?~%Q��fiJ��)˔�`S�.'�����k�˸ұ>2����r+oS�<5�;����u���jM�~�vʞ��4ZV@���S~�ێ�s��W����7(������n5�7�;���Q]^Y��Q/w�l�U��Z���b��#w�甥��#�_N�Iu�"u��9����Ƹ�g����ih%��<!�Qzmԅ�42\�BFE��z�nl݄!M7է��uG<C���V��Oi��x�M�E2��p�ͻ��3����Cv�R+��"�SO9X7��\�f/L�5<�D�rS�/T+�K�v�y��i�O.2y�����n�.��n�MB"�i]j-�?��}�	!�U{�HWw�g�0���zh�ě�����h�x^�X$���ٜ�SG�Bi�m��E
}�����"�����C�ED�8?*u�b0o{q��s'���~�;��TG"N�wp��kF��"��Ƭ�M*��'L$:����/@N��m�)��3�73�ˇ�%�ܱ\��N0=
Q0�R���̞�G�
���'	�o��LBq�WB�����X��̶5�O7e���igw���2F�"��
���)F�)m8�
�Hf��gkA��'S��e�ϊt^�l�>sX�N�/���$.UI(��	��O��M�n��t20T,D.ϻTH\���Ů: �Y D�|������E��m
���CEO���,�e��9�LΔ��0�
wϥv;�0�m�� O���Q��dܽﱋ��O"1k����r���6�N��=;Ȉ�؊�U�e��ϙt�=�{�o�6�G���ԟu�h,g �nkO��bd��T�	�v�]G��j�9�8�f�~c���5����.s��]�-I��v�AR��5;`z�Nh������_йٸ��$�/63%{և�D��,u�cu����f����I�X(P4��O;
�M}V��X�
��o^�eC���I�4��d8{�%��� jZ��u=�u�����3����6U~��?
7��je��W���$�� {��1��v��`fE\ԟ��4!*c�$+J�k�P��H�8-�P/�K�Z&�F�hFx�<89LUk��y���Oc_�wYڕ��==L�9�'�2Ij�����G��]uЁ��5#��_zn����l5nt��f2$�zQ�t��~=�>����}�f��d�l�=$N�s����I��m�ᜂ�rB��	��#|A�3��oR�ܚjl�D��/��
�ìl�'5R¤s�5cqd�t�]�}��V��ŵ,�sѐ�<����@ˎ����K��0O���%�@@��]��-�Q�K�	lVU�#�^�ʟ4ӄw���s��~F�|��n�^	-�R?�?�J2L��;��h��-S���Լ#��� �x���F�W���n�n4W����k�{5'?������1(-V��z8����7ԙe�֦���� ����'8�I8��l��Ol�^�J �98��S{�����ЪUa����br�F���>�`���4죹�:�
R���Y���uQ$;KÀ��`�'UN#Xsr�0=��;�r�{a��k�y�3E'(E�]�~�X�Q-�3/�r �T���5�%�l�]⏂!�G���V�10�^�}��4����Uһ/}Ufx�SG�!�>���<V6R^���p��d��uZ��Q)��o S���y�h�/���ӛ��Mu�[�o��t�i��7Ƹux��������v��N�qw&Jۑr��X-�:����AU�U�bnc�4%g��,����h�T���բ��]��,�e�C�'	q0����_�7^Y�k�7�g����ZȔ�ە���Q�+a�8��uh�Fx��L��%���C[����*ؑ�M�%1V�$����r��� Rt���Nz�Z�n�.N�lZJ���Q�c8<#�6� 9�*��0�({��1Ԋ���(�{ޛ�쀡YIF/s�!��?ː}v���#`M��:���V��(�{���"?0�ݢ�p=:���U��D�V�e[3�#�Ф�B�6�H|E�>��hG�Z�Č\��&f�����c�Op�j���D��?�	Q��n�1_n��X_n^$3^�5n{�:$� �t��_����`Ӊ���;+�A>I��g�#��O[�j��|���xpp�D�js�ȇ]M
F��؀��z=db�G���m�q.p�wVx"���X'�h���R)@�؟���y�� �ɏ�*�}H�o:��A����k����,�Ư�	�NT�{4R�y�FZyJN&"h�d;c��I�h�?��+���o`sU���CA�KO�Eƭ�
l�I򼢗9 G�&rb?�����L�S*Ew�x�pT��3 FR�~�,׮�YE1�o�|-��#w��%A�J�,(4�z3�;�Lߚ�G@�P��9��b�o��JSJ<��Ѭ�96"<)��������#`��d�B�U_s@*��K����'���q>���>87�jr]��<�F�ZEU{�Ӿ
��v����d��8��/���<`2�D���D�m�� �l��+��˚0�[���q��,�NE �P%$���F�Aݗ�!c��>V1q���k_����l%�帏��+t\_#�M'H)D�#	^��ڴ, ���W�f��C��4��wأ�Mc� 6+�u�[��߲x
R��T"�ҎyLe����56���D!���˺�G���rQ����_����N�p��1��n�zq��~���ɝ@*��m ���x�:nù�G�d�����k�Ͻ�QZ��mst�
�����*/oFw^J�Me�}��ҢFZx���fd��C�v���Y�2�O����'l'�ɨٸT�40G�R��[*�a� 7m0k(i��S5$Hv��b��t��9���|�
։����H�L�����l�K�fd��a������ΰ�9ƅG���⏺R6	���t	l�T`d��f~�k/��5�4M~+/�Wl��e��2�V��ܯ���v�v����m�+S�ddq��K�2��B�l#�UB�Dtw��N�;����2i�IX�R\z�=�1Yf<o+Ğ�{�q?�� �pu	���֠�H��Zc��t�l�_r��,Tn{œ����z�AxuNm�6�b�;��"�l7"܍�>S6������L���ifNs�w[ϒ&��V �,�e��=2����5L���@�=X�<�K�n�/o� ʺ�5t�K�Q��ϑ5 �]۰I��y>Nz�b�bw`����1�T��%>����`�7^cV]�d��=�i�3︸�i�qj��?��DM�1�).L�Y�N�ɖ�(��=b�^�Vt�"��-�°Wy�c�\����T���>�����;���£E���(�B�2w�Uh�p*[&ǭ��G��������}A�&&���_�! >K�9�*�5�p�sPFrY��)�C:I��.�n�ڢ��҇o�D�cnI�;�w�ƞ�TG=�Rn�f�O�d߂y��2���@C"5�E�a�E�z�1̪����-o�Úށ�� ��)_}[qq�\D�"�&���p�0�����~��"UK�h�}�OU����������Q����.褯3�R����J�lMw񠶀(͚6meM��!y٬��ULa�-fwc��usL�6N ����\��z~��SUv��< ��Lb���v�N�
���J�s����[��>����;����8�U�����ȳsݿeTJ���oL�����`�0��)��ꂒ�e1�d�$P�P����z�+�I+�O���� �Ȗ����)��yꂿJ&�a[LP�q�����J�C�������bJFc���}�8o.^��I�6{��"zTP����g��q��?�O�����;8S{mV���Dw[�z��V�	��P����v\&�wh3l�� 60Pfyˣ� ��,��̡mK%/"#r<���?��W!wQ�!�kGR������L�'�����{/H6-ρ�Ю��e�{�<���Fƙ9	Q��Zz� 6���{W|���W���Y#��t�l4�����S#[Y�?�����*��͋���:�I.�2r���C��:��O&�ٌ5�Xnf���y�-���6�u�>:�:�������.)�v��k�[/hw�9�6q�`
m|"ţ��z�M�T���ՑB���y}�e]U�z8#����*�G�_� �H���߳՘N�̠>g��Ul��
0�&Ū�4( x�6s�&� ��Y��C&Ɇ�ܒkM&�,�˵V�5�S+�&:#�rBRf�5�L�'��u��w�|��y������B�2Kr�	���+���ϴe:�Q�C-	��D�ٖ����:�,��=����_�]W<H�l ���Y��������43�W{�7K�� �
L�>�+J|��`�T��K�C8a��b�n�������5�c��S�8܄9�QV�zC�LO���z&�<k0ՐaƯ����|?����>��"n���g��ȵ>_�r�20D��!7a�����?��OS�N2�$V�L)��z^ �R��%O,�7:J�ˇ����;��R���/�� ~q+Q���Vo�x/���b��@s%}i�¹��S���[/͛�*��ݼՓ1�	�Q1��>V��|1��0����c?�O�u_�$e����@g3���we.�1;n2��]����������$$�
B��;���^)��c��-�����m�oНP!6^�1��f�0>.��s|�<r ��$�%�`��/�._H-��1y!��J:|3��	V�\NMp�B�f���杽e*�����������_�ڭ�D�}�ۏ��X6�e����ޒ�&�����v��c���릍|�
�/��l�V��UW�ᐮhH6��(�}Ϊ$3]�fu����j�@X�{�������f���L ��SS����`B� 5��9����
�>�I������G������K���\���ژ׿t��,�P1���e��@��y�ֲ�&]8v��@�&��Bj�FA�m�7>�;Ϋ��Ӝۣ�L�Z	��о��;�5���f�9�q໒|��\|��(�p���<t�;F�j`vv���Ԕ��&&���=�٨/E6���V@���o3>	8wi����7�2J�R�}�e�K	��7���e��A����.'��c�o� �3)�hCF=�
aZel��c����xυ�F����' j��#���l�|(&HͲ �����m�����YE���@/ґ8�g����V	�D��+�#��ÎM�b�3Gw�[�"�?~(�J�L��|���Pm���6ׅ�@��� Ui��v&j.��朗_3��f�T�Q��!xO���>�-J��J�=�<
�ITf�7���\x\<J�����f&�|zjMϊ�yW'ȥ��ܣǅ��%V��1�/�-�Ij�,%��?��0�J�u��4�A��#��Ve�+��~E.�Đ:p����Y-��o�;������-���z�k�u�y���������~`L���2ųtY�*UIH&�W�Bs��B���bxjq����1�Z�I;��=��+�c�(�`1.~���l�w��z��_;�a(�̰��3�-� ?:Nۡ-6?�T�j�f�����!)��+1�����d{Nk-�U�FM�ԝ�n�O,���!Ϊ�װ���D!w%T���l7f��6k�kE�z��|���=�|��`�.Uq:��	��$��8���5���~�(E���2~}�P}�K���SԨ���KL���
;�<Y�`�R���-!�/��D�u��ѝ�+7��HCa�����P�a���}��#�|�����}'��>�������y��ދ��&E�e*-�ኃ�1&	(&kG�ֆ|9c�	��4���E�j�N�p�Of�(K"տ�pB�c�����+5 �H��x�%��pzI���Z�y�cX#��e���eࠊ�8�!}=A�� �!���bf�Q��5Zl9�N��nr�5��`%G�)�%z(�$v�]�+q��>�1BVJR@H����.�o�6n%Tǣ�����DX)k����ǂ����y��V��i����֨�~ͽT2��{��t�0���(�G&;`5�E#�3���[tx�W���TvN#%��jF;	�[?��!P7ݦ�^~�)�֙�-���@L�V������g�	��ۏo����J*g
����ؽ^�$,^� �f�03J�cn�dnT�H'_�����ƪ�;�eR�ͧ��x�P���)
�"��:��S^�@?��EFh��M��q^tq}`��A0��P�	E4_����FΨ𷺻�J�6ԁ��O+g��ikh���jG	� �>>T�����^���{�8����˪�F�i��O%k<�C��k��s4��7���5=P�L:���$ع��c��?b���A������<2` Ag'�H������Qw�	��t����˯��E=I+=Ӱ��_�":�ߤh|���nk���h�50�7=�&�.y]k���L����
Bɬ�-Z����Yr!��b��a3.���b�����+���4[;**��Q�R2��k#�$��`���[�kkA!ʖ^��g�A76���ѣ"�~ϧZ_�VI�����B��Ň��~`�=��sXH�����|iWT��i���A鿡�	}�X��Qo�*�ysZv�pEo���;�XsA�P5��i�T3L6Yon&���!Hѩ���7���N����gfG@�̙��b�Ǡa�6!��9)� &�����͇��X�XD�߫���f6�^�w8��XC��e���p�y��w�`��^��'�]d,���?��\
O��A��l�o8C~k��5ч�u��l[
؛�g�"�����jc
u���e�B�
����c�@B���)�Vz���o�G�l�cw��f��a�aPa�V�.OబaI���;����Ш�_�닷��a~��Ŏ�: ���]��_p�1��[C�m QHe;���ݱ�����m_��[�j^ZM� ��)� �?)�_^�[qm�#j�� }���)���Ҩ��fʸc�7�;��N�F�R��1b����do�A#�
ѧ���k3ۧ�)H7���~<���vviq��ݨ0F+��+���D��ɺ�
�p) 堨l��>NPd$\a蜻�x�d�%�b^��,���a�!m7ڥ�v��Xv����V�:��\��Tq�TD�mڭ�5��(Qmڌ���F�zi�vC�F� NH�N+|���a9X�z���些��J��&�İ�P�$����)�g#��j@��L�{���ب�u d�,������w8Ke@�J��� 0�-�T#�)-k7[wC��j���;�����<��EE�/�L��_��� ��=;��%c�V� ���W�?v��Z�H��zK�Ge���0��JOON'!\,�}!���S��S#��%r�n$�$�5^��˻'Pܟ��Zs��K���0��$�3�¡Ö�^� ���42�K�x��ҚOg�b�����PY�qUK[��'v�V$
Q���C��AK��~��W�H|S�W����ef��bZK�g��ME?S�p\i��PR���<⿆e�$����R�y
1��6Gć�o-�:Zafz�T��2��Jj����)6�(�X�����L��<j|�
���Y1���
Q1O
���� �4�ħ{"8X	�M�>�A�\"��%w�mp�G2����gh�B�Б�8w?��a����Sf�'���nk��*h��é*xD�x�=&bʗt^Z93����}�j~�l��.��e���cHt�ߧ�^㈦��qv��-#$:��ϔaϬP���~rb�L�"d�^L`���C�n�F�%i]�p��e�ݒ��Nh5��~p*���dη�Y8���=�ץ����5O�Ocsk+�-t^��𠒅��n���:�!?i���.-UM�d��FC��̔�i�	�躷�S�"%t�Co�fj��$U��#�� "�Bm��-�Q*�":��m�XM`E?�ǅ��` �a8u��
e�Bq�L������F��uBl�5��܌?gsA��q7N�l��#�A�(h��d�)��7�WP���v!��
9&��PGnx�U��8�~�3�.a췇+����M��O��]RK�x$�G��u���>���d��!�����h��WNH<h]�[�E�og�h�"_�e�TG#0�ǰ��(KDk@��؋W� �?4�v0S<��0�3�zY���U],�*�r��,W)I�� i�CQ�� }�(�0<0-�3�3ʉ���My��w��O�p����n�b��BW}�i����ݘYb3\��n15��{g�bR�t�t�ё̜D��h��������r�n��J/��6]V�.P��	��� Z�^v���~�PoA��� ��0*�Jo�Et�y4�ReZ	>H�z{c��!{L|�0��㒖,�e�z�r�&�:�}d|�S��)����e���Y/s�X�U���)v�`���w��R�ǖc�B�K\6{q�$ �M�p�1���o<�ZY�5?	�5mp�+_ꅟp�Fp��`jޛ��T{I�Kq�_�������U�.�L�QC5��x��|f�`��Qq��2�":#7�j�6�x�c��Ȃ�!�|��z��uZ���ǋ��7㤷o=vww��p�Gy�9��{�ٽ�"��� �+W���7\?���_��;�I��m1q�W�s�1=MLN���_1�ȭ8���]�$�El��`�%��!��L��