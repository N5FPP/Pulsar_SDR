��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VYrF����̝���ySɎ�������)8�oT��!��U�j#�4�^�Cؾ�6�X&6����ԇ���l�i��I^h<�\�-K��T��io�! ��va)[9� }C�B��ǧ����������Ϩ��Ը<O���R���(TZ�l�D�u�V����%�aTxU/���/%΁s���V��������@P�P�@a�Ho0�o�#G������lC��Ƣ,�J�5ci��k�@9��ҷ�Q���n�xQz�i�T�k-�:{����V�Ji��`�*N0z��"������;�(�ҍ�|���dd(`l׺�x��t��π#��s� ?��)WAz+�Gv��J++�D��dU/�}���j���P���$-��=�_H�܏��� �M����k��]�ئ(�pj�}rG��A����p����] }�����R"U��yF�o�_���&=� ���3:�����������,������,�u�R��O�}����Q��[�����D[KZ.���FҽU![�v�Jb���g,�e������*ǻӟ�Qe��dX�/�]�OŞ�aHP��-���xZ�X�,	p�ݾ�1�s�o���P���jSFҹ��N|l�^я�ژ҈s}F�ٚ�-���k��
wW�V��H+J��k���<5w�����ZR<�6�R-�v�6�|%�\�CE���&���y���(:������j&��_m]y��x<�@� �l��p:��O����u���R���vh��Q0�O��V�-�m����G[��8ih2h����Ϊ#��̱��Kb��(7��;B�L��T�?��� e�e�d��q�^f�ΔČ֨�G�ϭ���*!=ȸ9����x�u���+��	��1�g�cW��Kw������.
���t�r�Q���<v� *g)\�jTl����|;�E�1s=��&�z���D�g�7ϔ��c�u��߶�dTc�$�аb���ȶ�������Wbd�u��/P�Kk4!��4(4�u�8P#YiQ0W 5n/<���(���2��f��Q�x��:�*Ch��g��P�X��W���,�B��~!z��r���Ӹ�V+򪾳����,��p�3����@ěaG��"�����I�����BX������.���(n ��[e�6��oT7'VG�'n��2�zǻCGEn(&6zq���g���
�>=����6���Թ`
����C�V�%�o�<�i5��6;]�fR5��(�G��ۧP�&荅C�9�~��
�P���;�@"� 3ȩ�	�r�r���|��[�|����0 'Lօ'��h������W�C��K�N����C�m�����7����ԭu}W�f���<U^Z ��0r|��&���,�.�}��x�yR�%�n����1A���"����'NBl{-a̫�tGM��\�Ƭ�
�_�6	۾����=��;���a戂��-US�ŧI,��P��=+�W�z2��`WϤ��|YpW��Q7�o���wi+�d��s��G|��J�:�et�[vI�+������67����tu�������e����S�k$O���&���4)���Cu�2m��\��&�3^+,'�4�Y��^xܙ�"��O�.`@YuPr��5�����$5j?���&�Z�Kt�Z���0��M)����̥pY�7��.7zӿ׫�|g�d���e=g���$��i:`��k�A��+���Ac���������b��ܷ���պN��C��a��!P�u;`�^cg��44��<���w��9(.�]�3�?�OB��Q9�z���[w�(B��U�N�p8I}�8��b���� ��{�
}���[� ;ʥ�ꇆ����Ƭ��X=6Ј���X)��`���@��6I�r�� ���$���Ql��$�ݎ�t;�;���%��JC/�^�uĭ^ۢ�>N��g����͕9��2������uП)<�v}��y� �����3�p
�N'1x|��?�Q>�z�D��/���o���U6�����sW{��ӈ�A�"�� gY��.+g-�d5��8F����x���ԯ��)�5 a�|C�2��>a���6���'�
�\-�k
I@�l9Xj���y�J�FM��'fß��F����f���M�2���<��Y����^�5�9��$Y�̯L�mdP��b|�5\��q��	NIܧ�fU�Z����n 
&���T�I,�^�+�z���k�'��;c��xq!�}��(�T/3#�Io�p�;�c��%�s 0��E��#}�v��|SdJ��,Tp&'�eL_]�Izp����$�X��6T���h�2]�Fk�[8?u�3�ᗆ�0�� �/���}}F��LJ��G�Ū�$�Z��T-�l�O6� z|��*x78����3^��y���ͬܺR�;���	>�!����?�X�Y�N�V�[��t�|�z�DW�	Z�Kt��k*���������-���*��{]��z}�j����4z+��:����^�=΍%m:G:�Hl��(�t����qH�ҍ`�:��pN|��w�����1�A����<�9��s�t�	�E��� ꏭ_����ɔ��	�;&���	BO�Y��Ă�\N��|��#�)�\�_ٸ=(&�u�jT�^�ִD�'|��F��?�W�o�"��[����X.,��X�Eq�r3J)�ި�Chx-C�P)�q�x����[+ ���߳���f貊�'���g-�!�rh<����.U�z�����ғ
-�fۧ����������M�V����9$���ׁ|ˊ�ص���=F��Qeſ.@�Si�����5�Ѩ�ü�4��_�F��B�"�
���) ��mSeh?��w��g�����@�MP��G�N���ͮ~���QEc���.+nmӐ�Awp�8���,aO�O ���7�u@��Vto�n���8�O�1p��2��',.�E7	��X���֡UU� 0A�Xfu����z�SH��0M��CiA�ʞ�t�_)�z}H9�g���)���ܯUJ�B	f�ڏ��Y�����7k�x�|P&�0�O����ٔ��6���nUf����H����_���"`|��%�i��lƖ0t��t�oK�Λ�e�"ʉاA%w�@,矵�+7w��R+���p����\��(Vkʎ����u��W���pj�!��?�]�����X�0U��L|���m־ɉ��*~�;K�����ݪIU��'����?�JVI�]P����r���8r���O5}PN�� Z���"0y���J2�yw�Euî��XB�.C��{8��w�E��6bM�Np��8ȇ�)���͒��H��f�@je�(3�~f�RN9�=Ԟbu�ޢ�l/��K�
s���\wi��6�����:a�w�hR)Q�N����E��cMze��rvVU �ޗ�L�p!=h���<�v|I5����@�z��!��NT�M*f_�/]�fjS�1�j�PBz�Q	��2�iӥ0�}[��^�����=k��~�3|�?�v���pX�z�)�X>��d�x���ȭO�ж���0F�v[�*
>4 =4!�����,Lt��^t��+��Y2�q��lj6�˶.���֞Q�P&"�V���g��e�5]-�t�("W�ک�W
�]�"�/T��π�mb"jZ8�p���o23 ��H,1��a�^� z"���� }+�d_��k?&�
����a�>9�|�Le���R�����3���˲�O����Хw��P�0��J�V�)�YɁpw�YO�d��������=V;����s��� T��a4^'݇m_
�����ԧ,��y\��m�^��|�<�ɤ���R�<���/k��:��������j�h��H�=�����?��:P-�y�;M6�0gԐQ���-�r]�.��ڽ�/�-T�@Y���
��j�������SaXX�T��,�Yl��	7h\i�u�J����j *����(�=5�I*k~!R��M���1�]?�W@��.�;�qanE���Z= ������vϩh9R4΄�M�܉������m��y���h�P�O)��-�R�����ŦE>\�(5������>�x4���G�Ym������U�����P�f�p�`F��H�՘"�s}3ܺ'C*����3�>*s9�8_a6�����_�̥��~9��v*�8X'�?��F�1ytb�&px������γ�B�}okM�GJ,u����:\�{b@�jB'������c^�i����R4Y��w��7��7�A>��#��
�(j��,��H��&�I	�Η���Vz��j� �PGQ����h]�Y�$jd�)W��3��%h ��ٞ[�0O�&��|Es�w���YC�[d'ˑqz꽐Ʋ�������#�`iS�����`1��u����ͬ�y�@�<��[G�E���)��" �����9"[��O���4�R*~Ł��z$T��x��hM��g�j	ٻ5��cR��}>�Zr�1L���R��W���g9xЅ�)��@�$�oiU�^�1S�
T��w�BV@"����h�"VЃ�!V����R?m�0��0EQ<!�����|���is�En����W`�������>K̨h�����j���r#r �����z)M�+0�>�4g��?��C���� R��r��[����v�c�<{e�ӎ9�娲�=�1�=����i���E2p'�a�L�|�QSe��C�9�~�2�qŅ	,���֢��#�n8�� Σ��RS`�:he]Ŀ�jP��N���	0�hN�(i��,u��gIS���^�R���'�n��h�7{O\۪���Ee�$�A�!����>�D�0�ޭ2�0��5��V5"��Z�m{ʪE�'��N����0�Y=�Z��l���I���}S�RsC��N��:����4$�=6�̌���~��<b�Eo�<�IKq(��v��L��oW������ڱU..3����il[��)�xGıߨ� �����d�a.K#v⑲�|�p���L���9��fd/?��L�C��c�,ת�cS/�{j��"���`���,k�h�$�`���gE�.ϖ'�f��e��bf�SoP�`��l�[I \�~�Grt�E���T� ��Cl�~|d��/�����5��
aRq4c���
����T� xS�1���W{j�x�w�`�#2HdC<
��t��LL��I��ٚ�{��G*�p�H�/_5Q+)W�c�:߽��=�}�!��������ٱ��OP_�zi�<��ЀH���O?K�RϨ�P��e���e��pOM��\I7�D&3z��:JW�km*�;�3���������T�A��.fù
�&�R�CT��x�բ����	$Zv��߭e��Y2ke�O���E�"�����h2�PL��N�F
�IR� {��/��۴\|�#b����4�Ps��A����*ʓ(��646����ȑq�ͳ�pd��*m����^�5��5d��n�
i"���*&Sѭ����Ε�#�5���o�yN���0(�A�+���J�ø�v�~��RD��Ր�E%��H���g�i��ؿ�Uh�('S>�o��3�)9\�R�rmCq�rݗ����ٓ2*����̨*I�Ο�� K�Z)��g��9�t5�u��'zT��p�k-�d,䟅1 U���� XD~>�c���+�xY�/^�Y$���`�-�b"A��{C�Ee~�y���|���Ȓ:�Ŏ���"�i��:a.pT*� o�6��A�^�2�Ӏ���@�C<�KL���?׋����7ת�� ӃO�0](W�R$��(� W⡫��i5+<���[�>�����M�g���- ���$�^f+81�u_�
��ZٌG�qv�F<������!J��s�%��t�"Y-Z�\����*���(g��=�ӱ�S�T��Y����شSᎀ@!���*�L�6^�%�"�}vE�{�޵������l*g��OG��:��<��B�O.!<�r�퐦��Y���*p��VW�iOF�8M�Gu�/��g��ZS����j:]l.Ļ�!\WK�T�9�{�Yt�����C��a/����b>"B~���}@3��Td��=3�݈-��?��<�V��|�v4���+ɢ��+��5T�T�*u�Kw=+�+��6��d�Bi�n�Vc�6����+
���IAG�6�J����Jv��`������x�
�sJd�	�%'��`��Vl[�R1��r�u�F�H0��c%R�W���t��lR���V�`5A�UZX����	/�x�I&�S�Ԩ3n# ���/T�ctOcc�"��z�[�-F�w��M`� ��s��`2�b��2��[B�5�Q�P���3aa{_��WUQ`�j��䍣��@�kWtJ�3B{Q�!*�I];��*E6�L�q	 ����/_Ӫ.�6PZ�����<��w�8{�v�(����-;��P.a�E$��$��͝<=*�������n���k��PMMdκ�g�INҬ鏨�qH�h��Q@�^HO��r�'#��b�vS��Ϩ�`�����8��w���F!��i������� ����50W����7t(��<y��]�W3�4x2�T��4�f�Y��3�=���k���A0���uCٽ�?f^�6�8'�"��߇�K4����y�ySl�g�/x�5<�a |B4���F5\��\b"Y+r(����:>�H�a̠$�z$ R��`�;���r��s9�u-�'K*3�qI
�	��P[@����?�(� ���|W�n��y�T��?s�g�����,Y�*�uN��+��3�1G�1�s�"
%)����^�azaX�{�X�.�_}^J�a�V�}�z9'* �hXU����_�r����J��}��
�L�>�}���J%؎N$P�w���������t�%S��,jH6��!⧹f����Kom��%��+{���;��ܦ_���R�c���<&���B�d� FF�j�q(H.epۦ�������ԫ��f��}��A�����T��)e��Wm�}��G�~tu�t3bM�#�)�w��L��mȌC@��G%�R+���W���->�CNh+�T��{���'�ͤ>�������%i_?Ҥ�k�����	����n!\
�Qw�'�3S(Dq�m�/��T0�>4�ѫ4��Xp=��Hj'�@`�?��I�Dj�-p�;.��/����w!r۞:���g���N�w?�HV	)����1�4y�bu���e�`�2�w?�25=�4����㒦�N�x�R�JHݒ����-7���T&�SW��[C%)|�/���rO�. "@�KGi�֪��qZ�^�UU˂�A��Ŀb�X�>��몥2~��y��6������(���.����V�$�%����e��5�Xd|�'A]���E}^\�e��-L����C�@�ٷ�Gs�V�I����ǉ�(��j�3%@����_�s�3�]/���ʥل�bq�5�uQ��]u# ���uY0��mz�k�R[��C���vH��:w�L�q��S��Bٯ�j3o�E���	i�����l����^z�-zw��.ubx��s�EQ��x��5W���Җ�7��-�1�'#qА}Vy�v��H�U��\���.�*�����E��_�?˂H\ݞ�L �J����Uv~6	gW�8��f��������9b�JD���}��0)�XS?�k�)ELY��Ϙ`e9
�; ?���n#�r.�]B(&��M��ԬYA�~���4����-/�����-�ub+��f\L��s��(��)���v�h��nهq� yt���cb ����6�pp��qJ�$BP{e-���kK&L��U��$�D/ɯ���=�qa~���xJ��'��e�m� ����Ze��F�~���Fý��R�F��s����" dFi�m���\X_�"-Vȳ�v���AGk�(��`�����MWI�Ρ`�JM)b�B��Z�O������֬��k�3�s_qƻ�I���0��)mbo��j��ƿc�J?V�Q�8!F.#����a�fֈ�؈����ɵ��A��6Ծ�3N,<(���k9�+�A��h<�i:�S��F�;���H�>�0�O�G���ZR�ޭ�Q��8�9i����Y�,k��dǔ���� ����`�����w�cD[+h�����EK�h�y΢�H�,1�K�Ә��p����0�$j�Z�^7����f�L�^�Ā�����������j�}�1��o��{E/R|at[��M�/��5޻���L����5D:r��[��Ԏ��rq�3zzďj
����iJ[�'�cn̽���aXym�o��r�,3f ��kLX�w��r !b>8��#r��5��|ȷ(��,h�=f��7{-+�{���PF�n
ZW��FO�l��F2q�@|�<��PI9�<K+'X$�[_����YF̠����D�8P����喽e3	�O�[��V&t��7t��8��Y�OJz���`px�!7� v����a�|�C��)�8�*���{f��)�4=[���"���*G:|��v�Ac��a4R�������ª����x�0�̑�c��R��,�bB,�曪F�� |X}��Z��sHw>�{-}����G�=I&�8��d`�0�Ӛ��4�%'�;��*�����q>�A%���|qA� �֕�/{��9��(a�9w�w�}H6��`��(�fk=�ᬠ����x�uͧi��425�q2��w:lI�ɉь��0�>UF�rk{�e�x&Ud��ɭ�	�.ὡ	r��96ƙꆴ���Z ށ�D�^�􆎷6?�	��#nY��=aǝ� �AG��(1į9�1����I�Wp��O.d[�t�x����`r�U�B���nZ�I��3�d�&��%(+圕��&`�ܞ�~H��D���콎0sI��ᕉ������4Ő�Cͦ�q���������v�.���5���SM�\ � ��L����#�>p� ��`�;��(�xϐ/	U�B���3�YlЀ�iC�b����*� w&(�u�&똗��1_�8��	0zC�������3�^���b���H��<e�#Ð6�HY������2!Z1^L*K����?r&;x'p�L�%LIA>o	5����d��r��fJ��ʅ	c:�k��q��O�����QP�ч�{j���#�v0�h5�$j|3�Fq�	��{�Ku0��H�S��Ȣ��d:��"��j/��"X��	,�6���H�l��t�dc��mI@	.Y�Y�u��Keץ4;��N�����
��,+���� ��<u�߰_&a`��ߨ���r�
��\�X�S�*u�]��ZST{xMhA��Ŋ���r=�A��٦�	%@d7���=��v�����{,��}!���v�z&�F���m7��WPѸZy�I�n�q����a&'��o"�tE�?x$�OJ@�|��!�
#�ް-Xѽ�=*[%nf���w��OM��Hܕ�e������f #�G>����l�o��?E,�����W���]���G3^�����M���m���ٰu����5D63�)sT���#f ˷~1����i���J��K�7O����_��(aU�2c,'��V��Bw�{��T�����fIή�����{��oN�hf)~b���������k���-��O?5�R�"Fi��T֦�V�{gG�%/�@�<-6��ِ����:���y]R�n5�9���š}�(����������AI`\��7��;�y�g�&�j�0YJ����_����Rs��/���s�� �Oܑu��A{���X`�;��rv��L��d�:���	���(�@8�%)�΃�=���nL���[ {~5Y��FE\XD	
=���+1k���ݝ��V-ѱF/��w��#���	�7��2,�g��K��r��ed���4��}�.�r"vEr�E_���G�8� ��ځ����Gr�z��?ǀN�g���Z5��Lv4A�,����?vaX_���H��:�A߯��]����M(q�M����$�[*	�1�ڽldtGP�`Y��4�N��M_�K�Oy�n�|��p�	b�V�Ip��Nr�单�[��PFO�G����]�S����`�Տ ��Vϥ��Ḍۨ<f^��%o4�?��3���v�_L�lC�ch�304��5�0D^��5�G?9[u��1*��p��v��d����Q�^�&�sk��N��AQT����f�=_�&�o�f߿s<���b���3*ԬT�b�.R΅(�eH>B�_�]������t��e<l ��]_�m���U�'j%�^�"p�)���2a���\̔�F�])>k������z�%�[������0��$@6A�>u䩭�Q�2��e����5,���g�1����(f��y��%Mi�"�|��qEO25zI�� �X�ν���"N�=K�����D�L{�g���%6EU�I閞Z������A�	�u�B���J��6���UBV����`�q�K��K��T.ު0r�w]D��E�D��9�~��)h]8P�Y�s~���|&g归b��;�H��q��D*at��;�u�?����D*$g��I�z=����@ȯ�9���˨��Q�з��'�6w�$ͧtt8�$�������6���?4#g�ު/%TF�&��3���C�ͳ���%���[��'�Ĺ24�,j~i�qx%�e�P�X��\�A4v_����;Y^�"Őf�2�o�W��Ү�6H�iY�5w�&�J�r�+yT//[���^j��:*��G��.~f�HD&�"�x�f=��C�%o'��C��Q>������5��0�F�����|���?Z�c3�Q`��md�f��ʭ����zמ#���Eb�!�����w6+{*F�nh���7k�Jt*3Y� ̚�4l�tͶ���SfQ{�X-�7kOw�����m/�X���Pe���&�	�!ھ��^F�+~��d����H��C�ى�`"��P���fR�@�"Lv"�.�:~7H,�w�f��`���VpOdeJ��I�V�O���Gg�*5RqJ�������Z��Vx��=G���F�!\�l�q��룬)G������+�/����gX�
"z����h�a`a��e�|�A�xs�?h��z��x�a7W6��T�Q�s��}�(� 5ځ�y�� �ߕ�	��Q�f�%y�����'m�LV�t�!¥��ζL�T�����X�P7���p��ȋ4���PU�K��M�vmd|Q�^�Ϝ�Y+��/=/-�2�d�������*�	ex� �[�QUKQ��0�3A��M�h�c�������pO����/�f/k���|&���$��qz.Sizoa����yW��c8����je������')��7�O�&��YF=�Ŭ@��rr��U=A��>�3q�Z��`�������X�A.� *t.�Y�g�b2�E�v"����A$���ɯҬ6B}��Wn�n�cW��K�T�-��e���b9|�A���`A�aL��5���#c!cm�O����(޳bJ
A�ˤ�*��2�`gMP)$�w~��߶#����	������Ƚ��pDE ��-�@����*5&�Y6+7U���(��O�|�ޫ�,�Z�ʽ(��Ih�+��HV J�dX�a,5�P���o��0ހm�'N��1)B�~����wL����i���2�����B5\������̍J5�V��)?��؋���mh�=E��-+wH����t�E����%q�y $Wx�E}�s�|{ɤ(����a� ޲��p�����b��k�xBW�4�%��� K+��!�3]BEG��q�^⭘	�8��d�pI�M?.Z�Emʄ��a��bj�52�a�
�*.���� �ʆk�G� �}�î�E�Y+M�准&X���DyF?m�-�\U��/6B���"C��4�� ��K��G�����rh`�G�xm�5����}Ps�L5���f��T:�P�h�Y�����{1��|>�uQ��D�s� �'F׆JV��@O��� ==$e^-���U��%>�O��~���@�|���5Lom�3�e�b<R�#��&��R�7TxI�� �X��|ō$ћGt��\܉�7��C�m��:�g����C?!W���Taڼ���7��?�G��~R��M;F��S��-��/��VI�b��ﾉ�ŵ��TԊڍ�Y�Q��k�	�ڬ�L�.��wL�7�U�Oo4,��D��
�����+2\tXW� ̆Jݟ�YR{`s6~��}6}�,7�Aҿ2�\av��pʹ�����	�ʅ=��~�h�p*���wj ��Që]��O�+��S�"�<M���Q�]��lF�`
Ϯp�����RR,,"���9\P�!^��6W�1���Z.����RYŝj��޽,P�e��Y.9H��J�ۜ�<�x4l^���*���v�KQq�t)���vI �FY�}hw'�
¬y���/� �i��C���Fs4��i!�@���� K�s�����8�i�בsSdfc��*�HΑn�]��AY#��PEm��-+����.Lec'�!���h�1���~��A��3���A����i߲(�xR�ph���ݤh �J�7*���Y��Ga�����*��A5@Plq~r�p�u"���{u���Ey��u�.f}�Y���a� ��d%��Z%d���&���hQ��:`�8ֲ����yމ0o��r#Ӝ�|Q�h��A�ԣ-��9I��q�H�/{%y�n�Z ?$Z'��u�8.\�������(��fV�yJI��6��Tջ�S�h��5��3���apr֚|����m29+�p>N�"'9�F},�W�I�o�_��k�In\�R]�@Y��){��L~��&+C���t�rd"�l��
#dPȥq�1��(�?;�Q���ȕWAE��.��@�V�?��zfe�u�h�ҝ6\g2F��h��(/]����?|[O�%!�~�-s|��+�@�}za��tVW��|��%c)�����_xho�!�-� �	x`p�l�"�p�(�f���O��3���I��i%X�p���!�A9�L,�	Lț
/�H�@1��L�qoe���y2�ӭ�N�T9�0�(3Nw]<j�����2�#�