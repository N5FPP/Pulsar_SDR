��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5o�h?\bv������Zr]�M�wM��a!��6���R�}���h���ƺ{K5I�*�q�p~"^g�3��j���;�ul��:m>s_`�i��wi��2������hL��ۭu�+U�u�.R��_�o���%�t�|�H-�*��I��x���yiI��`�iJk��B���e����O6��k��;�q_�׆�Y+�M���´}��E7!��J�Ż���p��_U띕Pݻ@�݅'"`&�1�`t�z��yE�W�z�Ͱ�NBi�YJ���VM���T�y�f�rf̟	�-M{�>!:D�N�9��!ċ��A(�j8����n[	��W�u#kNn�.0��$�Gݿ?&i�h����0�g�kq1�;���;���D�,]*Z���3�>YɬK��w�c�hx�]�B�d��ۈ�b���Y�C�.�e[�芬%!-�~�Xa7��ؤ=��7X���q���z�(��Q�P
�!_m
��"y�%��z���^�PS��N�T;������o�C$��No�qP75a�yHp.=su]�B^��9�u�oP���Y�VƎg�嬧���^ʑW+�C�BW�52K�?$#j�PXƝ�LGG�c�B�V�s��l�$J����*���1����h� J'HUg�|��P�������M�{@.YT�Jb�#�Bѓ�refU!�7��A!P-�O�Yx,5�u���N�Cي$#���v�հ��.A|:��Ec�-an����!������^�,3�"��ӳMp�T�֜K�� �#��/~�� �gvWRl�L�c��l�\Y�Z�'��R�"�>�<^���?�/3���c�_�]�EP#YDc����5@'�/��r-L�������^e��pH��G ���3vO�)��Mx�ܞT�z̀�#`�Ye}�8���c%�{����0]������ ��Ra�T9Mn<����])W�'׆C�:��$Z-Pp����m8��q��3�#���9�3Tz�g!�����)d|�xW���
^o���g�bEVl�C
3�+�렉+�x���bhN��)E�#e�)Be��|�v�m��ޛ!t}�|$m��rWe�;��4���9��Fpk��C��R�5Y؃"%*�e�J�7���@zC��u�Ø�5�Q?�7�v��k4��+���^���z�Z�=��e��{��^�A��n�k0��g�8�w����	����Fw�kn댴�c�
���"	���?ۉ;`j��@��Q�:'p�I<��w���_�jm�̒a<(�V�\��,���N�}5%�;��Y@�4����x☒�ƅ�C�hnl#Q�r4�tE�Z��=e�rh�s�$`��GAԖ�;�_�ws��r�')\��۝��k~U9�vMu�W�Sz�{r�L�90�w =�%�'nѷ��E�b�0��#`[���z��wg�g�L���>��
�<�����$ڀ�v����AQ�_�p�˽?���U��>/�m�����׽gjV��Q�� uҔ#�2|*,X�+m<��6ӯ-��m�L�$�ڑ��ν"r���S1幯D��E�Q�(x�>�%�����-q9��S�SEl�{uY�30�^��{z+�n#�:5�Zo�c}�y��R^8w��ͦ��;
?m��H�ԂX�������ߧ��2���Rܽ�h	�� ��ꗣ�6��p���?@fa4�W!ŗ�KZ���O7�[��3����\-"�.�7q:h�;���!T#��J�uǀ�N��n��9	s��; ��w�!�����;e7A��n�(r��˻�y�\�{eP���.K]��Om<$ԙ�tejѕ�߇�7��2�6W�r�c��A@��ǳ�S����b�fg���N@A��:_������6��ۋ"8�F�]��zЋ��O�g�Y�Q��/��H7�z�py�_t���I-��7�i�p���v0+C4y���LYa�bW�a�}�П�s���C�;X;�|~�Ӧ�V��t��W!�Q��C��.�Ns��ͧ���L���Qx`ʈjve�۞+7��sE��z����.1��j$�P ��ƽ�p�W`��x�����5��\�0^�[�r��8�
7M��F5x� ���^����SS����qNʜZ�����5�o�D����������Ok�w���O\pG�`��VS/���*�^�m3`8|� l�� dp���R,%���\[�ꍓq���;<��8(�*�C�D��;���^G�_1I# m��P�������i�IGf緷|.�4c�8��c"D`�(�/�9�����u�)�+����;��6]��x��SI�X�C��&��>�n������%\da��N�c��6?.Eja;��u�6.�U5�mį��P�"jZ��@����1k��ӻY�c���$����=�t��+�V��(����ORDq"��=�f_bv�( NX�궢f�I�e��&lHN~���(�(�`8u<�Ic��Ƚp��B!''���I�aX�����~@#xR���)�pԇ�U��9����\�SU|y��������F�:*��7���mC�ʥw�ϟS�:?�L�Ya ����1�?|����)3a��[��L�"�H~;��,;�;�z�eD���Y5]�O��՗z<Q�TSV�K���Gs�R�	�D>Tp�x����7>���˸��C��t����iĢ^��N�4��sx�����%��Eh���Fs�|��|�8��@B����]S�WĐ"P�p%,rE��S�L��mЫ���"2��(P�O֪��~x��	��T��
-��8I7�A�Mk `�v̂��mx�m��Q�����@<�m��[��ӁI�Կ��G��H�;@*5���i�=Ҙ�ִt����f}i4�v���"���Pk��o������C*=SF�����_
��k�̪�c���}h��=ֵs��ޱ������W�f��J�j�[}: ��!Ē-�g��O�=[Zb����{��@�B"�A�']��9�����p6��o��]OT���G��oT���Z� ~C�s�U��o�K� v�Pӿ��qMh�D~�c�>GG�r��0e���u���b�[G��za|��=Ӟ�~�V�YT���jU#'<��o�@��oؒ�6���� Y=�&OAEb��V��(����(��8k.4@v^���m�q*Iu!���m^4���n��*c=���z���e��	�����Hz��a����m4'�_sHN|8�� ��4��0]��:�$\�	:�w���c0��)8:v�[����YQ ��u/���؁��D����g������4���㩣�DX�e���H�

4����3���P�ni�������V�GR+� �ь�J`�L�:j(�w%4L�J,�9����|*?*,������y{>�jJ�?>C�Ă�LXA��<������z^��--V��Ⴤ���<OT9�'����iI�e�ǥ5��j3�j�*-:l�D!33r�lM`}j�T�F��/�#���$��L�U�ǐ�mTp� )'б��&��mŬbjTW�\��<�탉u�)0��� ���~����e�?:�; �w��T(W	#�2�|���h����!�~��sNZ����)����t�r��|F��Q��`��m	՗�p]q���wA1�c�c{�g��Ã�$"ŗ_uqȍ�F���|��R��~\D���3����V�K#���o_3M�a*�G�փ��%���gZ1U`0�$���C��ɸ�fc���Z��j��/M�C
	3�
��qC�S������ʭ�q�������O������0�A�&����_ۧ�9L>�Mӎ���i�H
3��߼�ZҎ��z?�ݸ;��![�}6ܕF����Ԙ�T�$}6&ڲ����lu�sG:	F	J�1�9�E��'6�ДP�l$C�O�Aᖆij�Wjt�$r�oc��T����q�!,w;�u��P���J笓���Q�셆�&8�ٶf����90�ۂ>C��J���N�)il�����O.�v����מ�EJ�I?�ǲD[����o��m����z&?���5��_��o%4|�L�Eƣ���I?�Ԙ��\2V�u$םͅ_	F'4)�j��V9a_e�������9b]V��t�_�����Ԕ(b�PEv�VL�T�k�4x�t�ѐƧA�D��w�CW�D��55����+}\T��l��~j,An�䄽�7�F���K�$|��ag�-���G?��n�~�yq�rq�?��H���>?�.h\�0|a
�FeS m1a0z 
S5	�\�|c��)t��'�4y���W#l����*1ϐ"x���{a���6�a��=f�jf�ak�*�$c��?��E�&ŝ��
=�3'��s���vR�:�z^c�w���-�n���Ӵ�#r@��U�्�k��R�Y��c����D�*����T3�n��2����t5��� 6�G��p���<�w)����J��F`�O�r�CP�G���c�K�fި
G�