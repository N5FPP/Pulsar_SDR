��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY�ً�r"�\��v�hh��PS��,��Q����dTkGӥ(�5uR�6ς�����o��X��|�ك_�a��草�L�/~㬷�^��v�F�����};�P0��0�\c�E�:.f������U�/�1��^/4���?|l��~�a�0�D��:�(�~m'"�G�I��D�[�Ms?� >����}<�	"�{�xi���x��8^�i&��a�"�m�;[F������#%tM����N�X��Nx���A�������5�VCu��A�6��@�aH�q{�V��ZƜ�PR��,���Q��Н�Y\��-L��K���_8��eW�W�)":޴���vI���ƍ��Vi��(Q[��=?ͼQa�.�#�$����v.4� z.���r���op|ε���"��!����h��@��$��j*�_L���RO⾧vp�,fX;t�F���%�"[u��{��P���:�q2-� ����֦��tӅ��e�z5$&��=�;D]�g�e�(�e��0�%cؐx���M:�=�����b�$s�:��P��}�$/6|'
�}\�=g!AU�����%Q�'a)�-
�ބ��[�$�5ý7��\�5�_�ރ��]��������O����çy}�{�7s�T�,�0�$�I�\�Y"���?	�-�v_l?�{���\$9���eی7#�S:7-�����'�cv�|/���&����ݬ�I<�勯lD+���6V4�B.C��6�Cq�2*?ۭ���k�30��=`�'��J���	�J����{�}��04~�XFT�����g��:"-�̇�c���B���}��p�3�;G��|��4�
�@��:���K<V��#D����^��Vab@������~���lMzvONQ�Z
K���!�hا=@��Q}nm:�z�	�4Cw Q9��ʚt:v(��9�G
�o�"��0�I��{"��dc'�\]h��kef(~i��4]͍.TX�W�0�	_��>��-B�d����A��M��j��P��"[��X�2�^�ԧ�����	�=����gy�q,�=�L���zs2Y��l�9�Sz�3^0�A�ҋ�>y��(O�
7�0������{/����V�0����y�9��`v�(����r�)<���?��'׻��	N~��VT~[�x�䀏B]Nﴣ�A�aS*P����
��o'K�;�\�\U"�)n�w�j���Nad��1X�qٺ���NQ��:�=�����g��؅��)�t(���$��]9��w�;м[�S>w��6tf�LN0<�3��i��:�#��r 3�.��ŉ��P�����$ZZd�M��r2V�K�Z�����Ȭ��(���z�n�p��scM9-��e\������p�qØt�@��K�̶�҆_���Gn����ۂ�A2�x�G�����ݠ��Pل�JsV��S�e֡�v��n����1�b�
��C_�+Bٴn�;|w���i9r�<EHwe῾��_c@[�8-�v����:��1��q$ei=�i}�h�� :���U>{�Z�A�tû'�0��&��xMEaUؼ�
�?����������h1 ��k���*�>������59�9���-�
ڜ��P�U_<�1���+�����c�HA�@�,��Wb�`��gb'S�k��J����#{D���G����"+?Q���߲��2��Hb�`-m��Fũ={}y�{�xCY����5kvB'�ｘ�]�e�O�Y�{-^�XL��ey�C�)�BA�I>cN ��}�O����;mef�$b�)�\'o~~7-#?i:��$�H;�����Uo�t����s,c\������^�Ae��`I6�:��p�ּ�� �`$Ͷ[蝌X����T6J�-��~���I}͆v�|o���m�.�k�TO�d5�C�������&1�_<����P�X�ar���7v!�2G���z�u�����(�g��o�^{��[ע#��6�-ed�pЮ�cu��	܆������v���6i�a�wā�c�JV�G����	�u�u(-6��kc?VIy���DuZb��K�x���D�:Կ:�v�����w����$�3��Q���o���9�RMd�BG�u���)r�̋�p�P������у@�S`��iZl�uFi�m`����(��!"���m]��;g�X@`ja9��{��53��r����� �e���T���7���gߋ̓�z7_�АWel���,�+Æ�ݘ F����.$���T�lN�����?�pi�ijB���m���P��ኽꄶL�I�1�m,b������Z"$w�.H����_��<����TA��V�y+�g¶��2�t֢�����ɍѵ��� ����������m�Z���Ic��y�����y���rg*��Ė΂��Qh�,��KHר����T6�c���}�K�A.i_\�P��*0[i����&��F� �]z��o�f�7R�V��5v�y��>~�����j�F=�f�ؽ��$� �e��EZްp'Ĵ/E�b+af���~8[�^ۚ�C�����kJ�7�x|� ����om8������>�k��z���;���Q�+�0��}����2�S�s����#����D�Ec��zkB�[�
3x��H9��#@,(:|Z���ȗL>�_5L$�w=uh}��DȻ�H��3q�DQ�s���9��j�d%]�"މ��Y���k�i��&0Z�,�Gq���l�<x��(�u�LZB�(V9)�Z�5:	�7
4+���x�`n���;ӕ��@(�0Qe�!�y�="�]����ϕ�
"�0P�54ٵ_'�Û[7��jU�:{�/���6A���U�Hu3��B.���ю9yx�}o�������|2��Pz-��C�>�:��$1HW`�^H�;��O1���N��]�,Z�5	Ę�SA����x���ӊܞ�-����m� �� :~@P��Y�|�ІŮ�J(�{f��ML�:�m�'m{�nUZd=����=Y�ڀKEWⶖFƆ��n��k�3=�:a�G��2��4�k<>C!<�����A=A�.k6��k�F��k�-1�N#+�͢���MԶ�McV�G
$e����q�&R������.�dܧt�a������z���>�G ��b�K:$�w}p��~�����|����o� 7�P�4U6�z��uvZR�	�Lu�nh��8��lF�
��D:�9�`���l��p�c����a�p�Va�$28g��.<�5�\��A��܋y�(2���,;9͂��w�iN-e,���Uj�8F)�<#by'�FI��7y̅�O�莒���s@t��	'�3��ڸ�G�ɾ#��%���r�D�}��iN�Z|R��(�w��n��JB�Rj�\���)�.�H�*��!k�Y$\9`�$u̍�6
"<8U�M��;�:��	d�?B��
m0K
Y�H�+(��Ë��7O���
�x����[%��k[leM��Gя짮����<�9���Λ�=�cNI��A��<�I)[��U�Ә꧈�i=�D�y'�pc�uI��,��%�_��UP���q�+�A�nZ�0�<���l�'nǗ6�>�k�-�,^ԗ� �I�X��1S�p����Q���ˎ��/'��Z�(=�n���c�0;�] _�T٩�������R!�/���\�p"&3��r`t&C\9oO��yb4���v@ڪ;?~lQh�Z�����Uـb}aC3� Gk�?'��急s]'�8���a�H�t��Q)�ko��#��a������GM�>4)��\/l�j
��+�y�����|�e@� oneB֤=�����{D�tpK�ڎ-�vȱYbK���E�y �5=PՁ�X^qc�hܴ�X���'歂K�J0��Q2���3�tGm{B���'�JVJ�M�`F.L�A�"T�g�Z�(�&���q�h�����^��V��В(���q�к�k_�L��Jj�i[�Ne���q�S��*sj��<���9���������+r��N��w����Z��k���"�*�h-�Xd��T0�)�3�::�D�G�D���!�E�l���	��q��G^�-O�X���(���qa��>e�����-|w���ܦr�y�J�=�\�qbQ/T#M�'�sHo�����k����X���Քd�+f9T����~�Aj�}����Se݈bN�ۃ��> �/���ewޅ��g�~������ѻU��!���4XHf?��d@�)U2�gR�R����WyZud�QC����[�";h������g�����M�1Z �	�����m�z��w�T̙j>�Ý���Y�%�K�]w'L���v^���B��3�`;.<�\�_X��]'O.����߃�����@��*�N�%�I��VЄq���A _��v�2����V9lrE�ş���+�]�hF���bEK�O�v��1[�Ϥs��N�HVl}�}��3hS/�<0�|_��$�Q�,�zb���W��V���38�P�ٹm¥���c� �$�'�*m�~&���\�/I1�Qu^��B1���h��Q{*S{J�c7�Q�=��h�3���_��?����5G&p�k��y�o�ɡP	��6k͞i��M��pc�r~���W�r�k������DNAp�� 4���(D�\��QE�Fģ-K��@/A�X������%/����Ql&��=�`ܭ��?�<�y
��V �m������[$'h2�k�-�`����D˻�fM��r�U��A��&k�2_KN�8��c�7h'��p��m1�3G,h:�z͓�}�l���f�^T��W��Yї�:/¤�n�z�،�	l�۾�^��h˻x5�n�V�mV��2ˋߙ}m��[���������j��J������ᕖ\Cp��~%�	lJҎ�AH�����	��M��؝t`�x8��[9�����C7 m��%��f�ϧ<>��}��Ư�wO�)�]�i��v2�EXU	�N�2��.f�3�F�!��wSH�FM���zz;uY�Q��|��5[	E_�(lyi��%�8ҹKO�I'����b%Q}HEv>{RH��?�.y%�����>�B{,ښ|@%D[�E��������=�<P1nR��*4���}aL���
�����^pS?��� Y��QI(_�
F�N=��B� ��ٕ�	� }!�8��Gna騌l��/�X��S�ք�ƤD��y��v������B �o4�?�j�ޜ�W��9:�2}�~:����� %��\¯��b��k��"�1H;�l|���k��+FW����˭���>���ٔǶ�T���a�z����Y�q���L�*aZ,�Z\���0ۋ#�H�?�k�����ߔ�F��a'���G�0g��}�y*�܃�PU�����;��+t�e. zKs�:n�i��|{\�I��yV��P��7x�q�YF�H�w��lY�M�c�6YL]���^�.�����d���l�gõ&�x�o/�?�2��T7'��v������"4����o|!�a!��ޥ7��#Xh�h��a�����^����J��7@�vxl��չ	�Fd���;��}��	��aE�gS��pI|�5�c؍1��S��j�ܫ������|�#�K�l���k�a���EG��>O�z���R�f}���`gm-��R�'��3ͶI�DTpPg}:�$�U�D���^�c�ܾg��4kʥ�x�[CM+/:<̫�W�S��~�~��Lp�:��s��Q�Bi3�D@��b�����!�ͱ����E�ѱ%:���y�Ռ15�BKe�l�U�1U��������k��^i��.E�\9�}X!�V,�tP&P8��E���O~-�w8R��gr�f5a��������#n� �>�Y[)Y�oŗ*M�c�6Oc_`����*��p�&W��Moi�{B�K���s<V��D1�>�Uvy� V���KW~ݛn�J��U��=VE�����6V�_P|�8��U0*|#���M���C#��-|?�?;ӓ��Z�B��3����򰔅Ќ0<c�1;�N2��b�6zb���DU�F#�6�NÙq1��!�d�~<��J���Xr��64��@��)B��!��{����K<q�_�U����m#2Ӄ�Y��q�Z���y�����_
/Ne%�!3$�u���XrL��#U߳eI���M$j\ԣ����"��+p��FF�4W�n�3LxPIN�'u����f��A��XFќN�MgB��+)�#��i� ��Huy[&2��$���عY���J&�Ǚ[n���gk��l��.��zF3�0��i�Hv�/&�jv� �A���[v�ݲi�C_Ccˌ��JQk�������U� ;�5t�LGi�`&�6�{
�d��T��d�pz�%��+II�K�������v�6�7������q��Y�8Pr�@�7���{μ�1��\h���1���7UvvS ����y�X��JB�$}"�/R�Le�^�kg`!r'�[����O���b\�T��`��h��Y"t�y�d�kEV=��%h�!���D�,�r�|uu�1�G���k��Fu����J����K�$��\��Bkv1��^���i��o/n� �3�U�B>p7���پxL�,7խ�iP�/�˦�2�o�������\kq�?o��31��N1a��ڙ]`�Z9�]�������M��<��	�13	�&$��q�*�v�X"�b1؞�	��g"�J	��2|fzp��7}B}�~�c�(3ŉmK�oZ���7���]��;�D���@��Jc�|(��|�5	\��ٱ���栎zk�d�i�+f<8��3Y��$O��7Qxr�9�G�ڝ��A>����6J�4H���;� �.��u����2`K�3�rR�e��ϕà�.��U�]#$l�����%l�ɮ�D��,'�5���>�I���NV��)�Pݾ^v�y��_�i�8���{PQ45��XV݁�5)�V�4��	L<LjZ#{+�U�(�!��
T���؍~rc�_����xx��"�`���<������HIqD5�kQQ3;���bK�&g�x�s��Q'��s>�s��c]d(�l�H�[���	����MBt@]ٽ�f-![���*��i���'�l߲���+����%*LfN�C�0��-��7O�����6����N[�ɉJK�@�������^���V���
Ƭ�5$�b���Vpt������� !�"���D��ԩ>�m#���±y��T
�I�;�q��l�hW�3k@e)`5P�������	��	���Ъ� 8Ae�������5乡,�o+�J���}!�zӧn^��*]�+˼� #��=�Q3�f_���I����Х����JK�� �?���QcA;!�~��j�j�
���9K��-5o���ܹ�t��NTa9�J;S�o��LOã�}>\S��Ȍ�M�˥�nLd����h���OA�$GE��i��k'���-oƷ�cT]��kG���%b���}X��B||�MG��D"�L�������"��Jf �NW�?��I|���r�ɼ'���ޥ�?�G=�]A<7��o�1���u %Ʀ_�^Ŋ�����$������_/`:�/�%�_��P��������&����@xn��$�K+�"��Az����H��	�K{�I��������=�Z3��y]Ҁo�g7%�	������9�P�)b��d�?��t$x^����1��-��y�Cco@��)�q93���+/|�]�T`2����i���mQ5w@�խ}��/}n�<�n���L�8��@,���b�O����P���\;��`ٟ�]ȑq�D;ԛ�|�}�����#(OG�])�U�����A�Fi�o�i���H����Ki��i�0m9~�������Q�v$�^����J��$f��},�/�Z(�h��n�H���Cw"$�4:�F���ҋ%�H@j��.��O�῞^�5�`���.�̫����B�y�K�]�$S;��KlFG_B�Ԩ�ᣭr�-_�#F�-=өkz�<V~��| ��ʎz�l$d�\�����n������e�ٛR΢���-�����2�t�C �j��h2�P1�5O~V�z�p��������x��p��.�+���S�B� ����$��`�P��.e�����z宫�[��-%�������3D8>�DBL���)�9~i�j���{�J�����gд���1d��X"�=t�y�=�_�Y�(H���cn׾[}��	�6�������Ă�8��tr�3�l�C̗�7]�<w]�࿙�ҨtU_�F��[��Ηe���EMVa�N�әڳ��z���}P.��bI�Z�Sl��=c�)�rh�fiM��;Ű��3u�#L�we��3��nX�s�m ��V(������JO��D�V�6`�v����m9M_�g�H�7}#�o�����C�O�-��K�,C�RV�ot��W��i������'~v��m|Iѳ"�{����j%��>�D��<���
�(*n�4�Q��	��� �W�o�l�AS�=:�o���|qs�{rr�@
� �g���s�Q�(�E�#�	�t�dXS~�!�^	եB�c�7��][�W�%u��ޓ��X�E���M����ws�'N����]pq|�_�¨�L���Ϳ!�)���Jv�m�c�8P�tU��~��#P��C%�؀	+�� ��8"GFG�Oh�Xo��bmM��Qow����`�AP����֤����0	Q������n�*J��b���?����<Ze�����r�>��������Н�T����Rrq3�cqdi��X�0J�atVJ{���i:5G�a��jO%>dc����w�����,ã���4W�d�,��V�����v�}�Uq�	N�ܟ�,��^�/I��<R,1B�)��������eV�NU(dp�s�)j	=p�?��hFs"�{tu�@�����I<�d�ܑ�Q~|]x;���1��:߅wl�O�(�|���QǏ+be�VC����ט����rh�2�q]Aa"q�)ǃ��|�b�\p1�&s�c}�d+�i?ѻ���y�i@�vVwx�kN�0]��5v�@;6�t����������G��^���t��7�[J���jX����_�l#�^������W������&�W�)��\��$ �D��i�=��7�#�L@��^)FCrWt"f�m�1N���̡�PG����}��Gؐ;��
ڽ���v���N�E0(Ƅ&�_���D�z�<�NC��}��];��v�ݼ]X�O|� Sj%^�|?�����?�A�����GܙM����_b�G+-�&��QԺK�yʡ�BRW2�\�<7�A�Z�8���1�����7:O�B���P�'�Eؾ��2�KV(W���dqͰ����O�#5ִ�%���կ���5� ��*=kRQ����!ݘl��M���s>Mup�y���,%��Li�;�]�	��6�g��7�5؄�?����5��C$�w�W\�AF��d��%��k�
�ok���?�b���C����]�S���!���C����s�s��xj���ٹ�ɱ���RK�W��@�s�����cS�&Zǫo�h�?qD�\.��Oۙ�N76��)��Υw��`ʾ1������Z�}�����y�yS�j�_���vL�[�9�r����6SH��0$������ Mu� ��_��̇5���6z[��6����A�.L3������N�ĳ��t��
<zt�Is�đ>a:�a�mq���b�T��z�.	�upA|}��e��EV"��Rq� %裏tO�>�e�U��m)9�U��Gc�]A3��]rMS������(;0��<�p\^]r�]���R�)DW
o���7l�@�Q��?���N��F�^wL��TqBR��(m�k����̏H&�>�뛸m�`� [4���4�\�> �(6�!���e}=ԋj0)���A>�J<�-;�A��!Q؈��/����
9v[��ꂯ�x����z;I��P0d���^!�C�7�ũ�*f��,��"�H�����,���؈ؙ>�5ϳ�rUS�]�a���moz���k%h
�N�2e@
��`�l�����Ҟ����|>�S�rᮉ�B37�uQ̲�֨,j."�"%1)�Aع;8k�������ρ�%���B�c�ƍ�<��>��[�E��\���`�6��G>+Ib�՚k����5I{��،�=A���32�x6#�vx��?����j^�3ě�Ș� Z�4��C����Ys���b��B�f2�H�qg���u�o�x����U#���Q';��Eb�J�xz�����iJ,ֿ�&m���JWu:A-��K�� ��&��/'����r2_�Jï]G�D�73u��^1gSfL�.~�W�$���*P1i����ˠ��sz�0~INgR�ڱ�C��Xǀ��k��5ߝR���\�=p2>bb�4K��?f�E�9��H��FmoKMs�v�1p��ɇɐ������B[	>ڏ\��t^��g*pxG�u1��7?\�l�f ���b)UN�pbK�U؝$ �QIqmA_�%u�\�A3~\���#g���l�?Y̪P��z�|�JhZ���&m�d�������z1`�.#�Ee�,Z�c�~`NV�%�����.�h##0o��LC@ξ��ɐgS���J����;��(���~dQ��Q(Ā�1��*����Z(Tm�H<d��?9��a%Y_0
z��e����µb�=9ܦk��f?�5�����o��yYY�n�
_��AA��ڤC�h�CW�f]@�2� ��p�8��aTD*>Y�M��Ѡ�C|+�WM�⩒@	�H�`���wH<c{C�ƳJ氽��d�z٧�Q�-ؐ٧h��Kɥ\���3�� ��0XLa��/~K��TE�I򧺜�~{�N]�o�%՘e�����T#�,���v��~�b��b�e�|���?zB�R����Z#��d�{oޤ?��M��3l�ϛ6�zݰ$�� @�o�x��̯����f/���wύ��#E{N��!:ʁ)K^U�%uX�.�p�Iq�[�p���D`ge9���9�!	��q����]nX�/c��e+*��e��!���2����Yn�	q�ӫ��D��i뗛��[1/)3�xl����=ӯ� �����^i��J
R�ߐ_#Q�=����X�WLGRͮ?�@d��[J($D+�K��rD�]&�II!��
���,��p(<�_&� ��Y� ��1��@���~90�.Y47�)3���gK��n�
ݓ/������pM(ފ&į8�I��ƣF��H[u8M�*��Ļ��'����u.�n�����y+KG�K�\o����|\�����' eϷ=o��-.�5�z�	(�-�aQ���<� 2�_�>n
}�hЄЏ�9 �JȀ�G7K���F|���~�:�� �pX��7ȁ}E:�>��9�Č�����ǪCk1�4����A���J�=�-�o�+�����6I'�������7���''�י00���:/x|8#�QC��4�	ڊ��/{���t�ě0�[�\�-����� ya
�J&�����4�l�=��tnG�B���,��+�����
6��M�-�^"r�ɰ
&x�3%n��^6�;I�D��~\U�Y�	^ˏ��t�����~��ԤQ)m���ۏ�o�
!2l�l��dy.'��
p�����ż�-�C� �`w�`��0��UK�)�W�[�:E�Ȭ�UJ����w�.8=t�O���!�U�P]�� ��2�?��Q��+O�b_� ,5�XeKc��[�h��� B��+U�;b�h�6饻����^b!L\�?a�W7�]���:��[)1vBW�D�zy�7�	l+'�#*SP�@7�,O�Ge�f�é>�=����f��dz���z��w��{V�����ɨl���u��u��q��5.���vo.4Bv���q%��\-gn�/AA	f����j&�y#�{:�r�$[��r�ȉ�����s��j��i�[��c叫��S�Pk�o��r^N���Q-@�("B�6.�}T�F�Fн?�ⵓx���͏��E��Ν;���Hk�](����+��4�1���N)��`����&�+����H�9��=0��#L�v�*e���*�X�ױ}�ެz"p��ktR�y��eA�j�.����	R�4�����������Qh�0x�B����Vҝ�$^�팃��f���uܛ��*+O��y����ܐ�4f'�8��oY� e�m0�WXc:`Հ7F�tZ� ��1���`w;��[�N�)��7q5�\�0�ٝuH�䔬[/:��""CR++�k�lF�^KVW�s[ݢ�(���$`��uF�}��j��[�6-c����N��6߲�,g4�~Ӣ�/]�&���IH��G���4J�ò�$1H���bх$���p��mW:b<2<����r#��<j�������t��aQ�F:�V;v6.��G9p�97<�j�J��Ԑ�}1���y
)䏡�d��l:��މ	�!l^���Q� ��__@'�٭�L%_@jH�~FZJ�P�&>���hR�d�"�]���/�w7��l��8�%��Q,��b����
�;R}��~{L�~ƭҗ���"����0�#��COI���ތǑ����ݟ�N���rv��6?FUU��`�O��ø���y�RB���ui�5d#���Se�2�#E��p�B09�xUA���uy�u�e)q�{>>�|�|/�>\� ?և�O���Q�W�V\�ʸ��b'�G�gj�*��������p�\ã��[9�h����i����h���\E�������hPӽ��om���Bk���L�E��e*�����vR�)�P�'!#!a��%��>y�]��:D��V��a#+b�{bi�>�;H�O� *?�/�C���U�>}����=�`���})��Gx��ߓY�sS�����~:� ͟�9Ҝ��{eޣ0���y��ܢ(e
~be˦=C������rꁦ�"��0�zx���v����+P�L8PY�?�Y�m;��Y-��\k��Ԟ����֬~}_�#�MMWJ�ԡ=Ht�p���_ƗD�hg`\7��=υv�-��8Na���n%y35�������%l7җ@ٕ$6!	�j �by���Q(�d�a�`��z#'��u��Дw�R98+����<�5m�ѩ@=2�Џ���%"��α	�<��x ��0��Rf8�3�j�>4:0Ep�z��T�^���]�ڠ�������My�0��u'���K�v<)MT�����n�D�?�K}J�<��(V���lT5��? �O!��b�mih*�����m�*��4����ځrGJ����y3SQ�;���M�)w ?�C*5��	�ُ�L�xv����b"��"���Q�Y����X�{h��N�EY�����٭����hPr����vz�SSGQN<����`�C�CRl�ᔵ�vɂ-Q,�E��Y}��K<�}�7�,�W=�� �v�nU���TG�ʇ:��HK��f���p�����//;v�L�9� �Y$;��g'2���{*�|bDk�"u�II����3�8���UWj�6�i�.��\��WS�Z�8K��`��)fnǴ#�h��
�H�t�3�6t�*`�?���?�Y?�k4�"��@Gz`��!I+��r�&6��%��߷XebH�&�$��5in�7p��?����e5�2+j��؞�2M��b��{��O�TкF��M���{��w��Z�MJ٥��/8 օRc�k���Nt�K��C�&���|mX|�vx��,��<%�j4s��oG����գ)=�uj8�/Kl�k�$���O���1w�ہ ����EG��W�fa�9>-H�v5���j�j�<�aC�exw�`L�,��!�a�y�:Z��I�|���*�AuO�Fx��q(��Y@~L�1��G㌖ӡ�\0,���"��po�4
�Η_�E�n��^�AD�����~�@�r$�$|@­�O��Ř�w~�'�1j�c��k,�H����'ף�,�9�:���,6��.������*�A��̦���r�ӄ���j����IC00��U�ݞ|!��ՊE\8��
��D�D8C�,�k�/����� �Ҷ����j�
������Tݯ�-N.CY�|~ȭa� a��a{���Y)�lp,y�^�)�r�%�	e�?��kR��]��)A��jW��h���HÏ��ڞ���N�.���ǧq�DF?x�s�؂� ����&x��}H�D�]ɋ���3$���,��l��d����s�y3��,���P`�@��+Ӊ�$�+C���Ąu�W�Ɲ"c�Me/�4By/Q&�i�s�>r(��Yȝ:��l�f�2[N4�k�xIO�8�26.5r��k@��qA��~�L~�dmϗbꘚ(Q;�0(<xa
R6�X"�5W�z���%:�����8E���HC8���m�~���*��v���3�q�y0	���7�٤-�Y�g�Z���|Kn��q��.Y���#N@�Ѝ���y�I��F.�U�f�~�%���uA���nf�|5�#�uӮ���N��� �����&4���*�\�^����櫑A��n�k�l�o������ ;}�F�F��R�^�7wJ�}�(o��ct'�F�����y�_�ބ%�&�t?�8�$��[U�A��t�h4��h��&��ܣ�b�Г�e��|��ۋ��$�zu�τ��=W�^�,��A>�;��T�)��7*^���hQMyO�KRt�W�.�M�͙3�Ӱ/\?Pn!/��{��2���H�JM3�vb��-����}��ƒ��!m��v��);���eŽ�g��Wd	eXC���O��k��AD�o�Ԏ�ME#��,�$�S�ʀlF�0�c�ζXf��������#?w�Y@�V�t�;��h��j���"u��R�n��I��@ݘ���u
s#��^^1��4���%��t��|i��G%@�`���؄gȲ�F/P��q�P�y�.�	j�ej��Y� ���d�zc�����w!
x�yi� �6'4�}(C��b�\ooq0��J��r�jX�UI�F�Q���Yјm�z�5�5�c�$O�˗Vn��/ئ�7�O}�� H�0�}�����U��Q���6[�U�LF[��ڝ�pDܲ�Z�J��t$�Y�����Xr|e�f�Zp�sU��B��n���H�5�wNl&F>C�7J�s�3�N����d��L��cz����C�a���g�,L7���N�9��e���j��Zj�!=c��2[����QS�p�E{�! ��	$O)�d�]������2	\9 6C�'��dǶ��_���/4L *�
�}�����`ȯIy-#�6��ب�*����=Ţ"�x\���t�O��2�c�w�>P^2���c{�$�$���U���u�E����-�׊�ř�}�~�vط{E2��WĻ��rB��%$�[/J���r����_�(�}W}wdE���r��&�mG�烷A�j�7~�� A��٧#u�i��JO�.��[{�!V�[��:@�Cs<�펗4瘈
L�m�I[kʫ��ч�N�=�z���:��f9��pX�v+JHU��)ʫ�F��kE Ay��<+&��$�D!�s�Y~���'����&�����9��70` "ǝ9<�ʾ�
@q[�\onG�e���Q���<:��,E�4I��\�Õ��:X��l	�*d-������:��b+�
Cyd��(�!�����$�x�x�Ww�Im����[�zv����;�X����d�ק
iA #����)p�L믥�IO ��W<���S�������1�06�s��_�&��Y�Cy� �M��{�{�[h�L��w�����iF�S0E���,:�h�6t�0�U2E���`f��:�H�1N=>��`�V#��3+�6��9����r�����/���o����b�'���NA�_����rl�}����ͭ�P�-�oZڎꖈ�U(�����\�i��߱<⤹�1��\��+�2}Ϟ1;wV!u(K�^S&�!����#2g0`v��b��Z�^pa����^	�bA�2p�'_Cʬn92�l �]0�_:�-�tT����"�F�j:�q�7:�sˍJ΋��wU$tSTꎲI�������Ȳ]:��0�w���lt��
��HN��+�wіs,QؑD]`�����]N��N�|_��x�&Ï�D��e=��Z�pg���b��4b���ف"W�~���tFJ�_��	:�_)��J�e�U I�!p��)3�k�q����%{�	��oe���D��jjb,����ƍ��`��X��5��(e��t��Z���{z�f�T�I
/TW��c� ���ź�
�d��G�X����"m�H�ۻ���^���@�{�4�M�Gj��@�dyuĥ��V��	i60Is��+?;O��r���<�rb��SJڽ�,��b6�9:��xEH�h�=�둥��l�'־��X:%E��j=&I�{-d��}b�v[뺦
"������l��C��H94z�dJ��} %oް�O1N� '����Qag��;+aVW>�t<���]���P�\Vs�Z#55�=�����0�`��S��a9�*>:�2�� !p�`�S���Q�n�������4>j��$u��[�u�_>�n�*�}kn���!��_��@48�Hd7r�|Ya�������
]�ˇ(ΉVA�2K�{�j4h3���Q}?�9QD:�څQxu�vX-���0*��NN���܈�c#w=�%�cg���l����3���˥��qu;��U(ҏ���ͬIA�S�u�n��C|!�G/2��(��}߸n��c��Z�$~�+Y7-`9}������T�}y���L^��&���)kV���@~H�-,�i���M�N2��ovj7yp�X�m�q�F|�e�Cd-"�J�l��`�s����x��Z�B�۪�t[�W���(��� s�L�H�;�������5{�<Ǎ�A�{�J��|�6k\��A\z.�S�ʢ�ߐ�/b{&� $�58h��K4�6�B1&�H:�=�2ʡ���16YO�ʽ����:�	�	�(xV���Յ˟�a��p%U]��Y�F��4���zΥ�z����l�ZRf1`��� �'?�]P�-]��c>1�>�n����@��t,?�ᔶ{=�$�B��L��kX������1�Һ��tw�p��@ձնI����n<��W%}��>8��)C)�/���E�ʱ��-�ϒ�z�8�� %��V5��<��/=�^�T�D�i�{q�~���C#z���W�I٘�,�;��&�l�RSn��7�C��:b?�Hnհ��~��S�s1��N[w��N�m�c�%Q��1Ζ1����z�%w��7Fl9�ahi��YI�4�2�?�~y����
�yD��K@�p�PU���JΡjV����mz��`YU���e�w?�H?�4� li�<���pG�<\�7�Q1�P�*Zj-x�Mw�8��P���z�6���,��m�x�~^?���tSX�W�����Te���oڊ�,/y�`�0��d�F
&Tuٻ���|{I�SJ��(CWH\Ѐ�Gb�?$�	������J뜎#˲�#�k,���I�k�x5���B��v�^�[Q�}`��/�aw0�+����͎k2gWd�5�x�����VA�CeI�0��;�,T�Z�M�/#�h��� 2���&�Tw��|�6�i��m��@?kt/Z���j����PtL�x�g��{��!�M�^Ji-յD0N=�v��B�����=�,���w5yI_:���+3�fy*�A����#[*p[�ɀBT�_5�mF钋2���SLB���n�6�<��W���ߑ2�+�9�А	X��A�Ϣƭ�^[�:����8��nú�kl��]�oz�˺����[J�}�p�w4��_�u�u'���7Ƚ��첗�^��k�Ă�*��y.���f�=����>Q�,�>��Glz~��Z��7�:nr􊰐ֶ ���(>碢Fa���H�T1@��A��^d�3e��C��IX�=��8���]g��\?�z��e��1�:��K�u ����:<� 1��ϴ�[���p�Jr��r�n��k�OA�2�m�#^-̻�xEv$�\�!SY;�n��^֒���KBo.��r�5	L�~ra����`�[��~C�i���N6r)�2$�ZO��'�rb�+�*�� �Z�q�}k���
"9�1y���M��a#a{���S��
փ+ފ
W<�rԇj�t1���U�������Zg��p.x7L+,v�<�h��g�����1�(�����z����㰸�k����Φ�ͫl��7�Yv�����p��t荪��K4w}�j�Y.��X�F��dg`�\;�����4�)�2t�6��!���ق���:��G�ġ�(�D]��͕b���	�$��F�q��[;C�,���].���LD��Z*.��qt�f;��<��t	�2<g=N�OA�&XzO��|��"ŷ׎�=/y�V��+� ���%�x�[\1saۜʐ���s@O���U[�E؍�%^��@������1f��p;��ca�&V^��B�z��}�bhs��>Ljmj�v4K�0"?�~���1�=���]I$*�1A(��[tQ9�ÍdA��2��ѵ�g�!�bS�"������IGqDŜ6����zxӱ��m^�.��]�|@��J�� �ւ�O�}�ڀ>��G��/�{�9���h]A����Cd�gB3���RBɾ�@2���%�if�pu�.���^0X�<��ۢ<J6$0�˴�[��X�d��æH�M\��h۲&;�𥎋���#=���A�J�gEd�5��>�����N%-ƅ��A�y�P�~��יxع�����bI�+�hc� ���m떑aw8w���!����0�b�o�]`W��)��7�g0%����}��c��2�&��Z6_����qt�WI�}^�F��q�s�Z��	�{���s���;Wf۝�]�׳���3W����O�b@��-�"�G�f����A��J2�e��f�X+w'0��������(U �x�?�������<��:V@J쬢'��-�j���*Xm-y�J�Q�h�~ X�LL>������pO�'Ʌ��6a8�%f�";
��Q��`��v���;�� �p��$>'=$�e�����1�ۧ�H5��av�r���2�w�I�|>�cl	�m^L��.��GQNs�ЛF�R���x�	����-��.�
{������o�`y�9�����ϓ��wL6�!�ѡ��|���"����_}l�
Nj'ҷxο�����YE(=1�u+�d(���o���B#y'O f?�<����=��.���1�WSEp-�m�%�Q���z���n$VN��Ht���2� �6U�1�Cl�&X�2C5��s�G�c��J5��߃�����q	�1�qIj^�㰶��sJ=X��IIL�3 ���G��Wx:bp.���o9,�"T�����~y�;�m�!?t�q/�����+�{{]U �#�Lv.rP̿P�8����M�7#�{����'�55t�frx��fLAX2�p����
Q�yE��W� �y	S��^T�I����� �f�[+��|^ˈ�&�"���8E0��r1����YR"|bes���|���kM�gr9c����3e޷���v�,0!���[OKNqL� �)2 ����y@grK��V�k̴hTϝ�#A镆�ڍ�ebg.� ;
T�0cn��jH_*�S�:�oB!�������^q(�YD�uH*�:V����d�(ɳ�P?�1:1,�ӞH1�O}��5���56��*�S� ���`c�aO���ܶC��ß��v~],U�Wi�{�T� �����6� 2��ɬ�=$����5��<�w+]� "�d���P�"AG���ݟ�-����-7ktfҖ�#��t�}3��Y��AH�PBBf-�asn|u�`��2
�oA�9����ؾ��>��L	���ZM�P�T��:�L�1�5��	�������L~�[�{/죟�B�Y�?q��f?͹]���MUB/��U`�y-hԆ�ڠ��g1B�~�J�%I��L���B���������� ~�/�J׺�b�^�^T���(T-:BZÚ��:�N�����i���@h~�f�\j��]��CYH�!��ˣy/#�Z$PE����������t׬p��y����M�➂T�ŗ��!ܒNeT��z��_�/!#)�*�-�4����Hx���>'C�!�ƅ5�����{�!�h�_����I) �	"����8��gN�@*i�����w���6��\����j�B]�E��6G��5cE�?h�cׂ�;�O�lW�]	QI�x��A�S���7fr�
4ԋma3���!Nj�ǆ��׼o��P^�H@0_��,�}����^��nv8��e��Y��*�4��=8v����#��I��]�x��46��=x��bx��ה#���DQ�� ���q$d>F���|O�ZMJ��~���� g��~�#7�P6d�?eN9����A�6���s�p��/�C��K#���>�}x�+u@�6oQ��-a0�FSU)�ơ�������fB/���"b��}�X�����%5�K?��E�	@�� ��d�z^�2֌��8�I�JuQn���s0Hg|M�GJIY�	���`�8�`��bt�W,ڨ�q>7A�/�涞�Xm��8_��_�+@� ����0�t�W�Og����v	�{�1�.��x���]O��y�v�#�D5ZOh��r��?�dV�
�a�m\Ձ��hsZ{h�>�r Ͻ.�F�1��*���۰�F�9OR�|�8��S\>?T��r�
8]IB����ID0]T��Ħ���D`fS����]�{��E!j�͘o�x{j��!���c<]gԗ]ɍA_U�7��&�J�Ƙ����"h7�\�[���-�X��q�Sbt��2e#5�w-8�I�q�V<��i*"�DV}�7y��-F��a�I���/�Z�`�uV*��0&���-y5dU��ۈ�n��;2��l���a���7�$������L���I��3d�����^��P�xl�m��`?L^nA�e ]� i?-�o��6��V����p�4a�q����	��q92z��*��oqq��ҞRQ�4�LENݡ�E��$�$��uM\V��'�
)�5��qBL-	&�c9�iYrO�a�2��?+ySI'���(�-b�b�k�������6a��UjMp���ɒ%���D�J�������2+���*�@O	ŨG���
�xp`Q������72�ќ@N3�1�}edI�����3��wǀ��6��ް�[��H9��!tvJ2M��,!��XVO��U2��T�>��y8A����wdp�ۅ�K���+�����i�^7x�d!�0�.��|��;�#��6�����V�E0j�t�C(	A f���Tb�J�����PS�,)��p�[̈���P���3�X�� #3����0U}U�5��vm.�����7i4e1��ab2 .-	6A�=�3
J�~�$�iH�_�W��jf�B�x#���6�����[_�x��1�1�a�`]�-���?Ɓ�+�}�cq)BT��ʋj4|�O�=���4R�H�n�a��r�=����� ;�`� .ROIa�q��xg�ܺf���~bf.-ZAı��y�t�Q��[X�n�kf����_�J�١���=�چT��U��UR4ŝ,$Bdѕ��}~�[�K��ݧJ����wAF����G��ލ묳(|�� dwǄ-�4u`V����e�m�k����ǦlÐ��	+��v��b�G$�^��qm�\��i/��L��(]�����٨�A��t���5rH��,j
o���2��D��Jda��W�t����0�m[:۸���4��o(�|���oP0�=���.TI68z�r_O�{�\�5d�J�G��L:',Ρ�W�FeV./i�`��֮l�IJ�i�ƃL�����I��tR�-/J���A�
��;7���m���{cP��
V^H��z� e�Ij�l@%DZ)m�CO�TcO�"ց���nA�5��1����j��+ɵ
���Ӣ6�}8Wbd�ӝHp��[��ҧQ>\n�e�{�7r��=2��z	���Iw��gkRI����F�4h�?���L%�z�_�)�kz����͜(�7n�h�$N2;����3&����U��Z�c���XȈ��������/c�pnnI��&�������'�"}o�� mz���^�Gzd�#�U�0r��`��'��72Z�"K��E��Md1d����]���{[9 C���P22�}��w/H�A��94Q�R������m���h�:{��"p��F�'v?��w���j�5 ���?7���߶�R*����µ�R��,����c�t^�2(�7��5h����i�Я�
 ?�wb��t�m�gu�z�
�<I<7\��������c�����:=���Fd� I��|�-Iq�=�U$	L��I��DNrcǍ���rγw;b�5g{Ӽ��a��~$�w�Ng����:N<ݑ�$��Ғc��(��%  ]zh�Rq�=�T��a����3���a�\�(�s���Rr]e�ͲF�<o�D�L� hk�G�Kv!✼��l�am�ʋ05�KÒ4�Ŧ@`H���)��� S׼c��u��7y�̫S���MwW�����b����>2��ë ���o0o�B���[���G�W�G��
��3C���,��T;tk���5�I�ΖU���۲J��Dz,�?��h���Ê4�2e�|��5&��y��!�@����Ǽ6�ɝQ#~�^T=#|�~+�g:��!� � j�-y�{�-���[!�hU��(L(�����`�:�:V�y�?ı)7��a�4A�{�9y��s�Ñ�*�Pl�_��N��VJvҚ��l先��-.w��n�Ƶ'92;'�K�hB�|`B줝4���wF�^��4#h�?kh�K!zG�l���ܼ��D����(%�0���Õ�D��b��2 l{b��9�2�_a�&?�ZA���r(hV[�j!a�$��G&���ӈ�����W��_O���ѹ2OGE�lە��ă��v��/zぎ�K�����{�<v���g����3���CXv�ҨR�:�0�Q��J������		L�r�P�'u� "�/�B�W���_��mlܔs���oBճQ������T�u�0�UI��i0�o�˗a��\�T6���Ҳ[&��CIE@�o|�u=��h#��RU#������I�`�~�@2?�*#�4j��t�v�ř��gq3��+v���tŒn"��z����{��͠�fK�TWT	Qې.@{R9�S��qv;c�Q� e�d�:׳�
Y�>2��&_}u�;��~?����o.DZjk����L!��rB�YЄ5�'�S���8!y6%tL�s/��	���Y�����/ڲ�ͱ	�7PXѢ�+��"��č%�6x�ƥ��-8N��$���s�Q�߼�]}-�ў�o��l��� �P���>��ITK�{
�30��L�?q8P��#��+Yb[:6n��6E���X�Νo��������UU������0[p��U�ˍ���t.|X�H���?ώ�M����i�mm�\��}���.�4����Ġ0��p�5h�����71u�)7;?��wm�;��c.+���?�F_HYL�Rd��ع+��;k�N�,�'�w[�_C8���!����G��_��Z(�X=;\�ILf9����ﶛ�C��l.Sk��0{���g6eMs.'e L<9�� ,�%�g)6���
�e�����I�4AX����U�ǳq��"X�q��F���s��ݣ�$D:NY̿�a���Ң��:!�c�Chȭz�0I�7V�cm+�'W(��J}L\�o0b�d[`jƍ��x�D�؊����.~�(X�AC���OE�.�X�V_��-�#��S�zxPpv�`2\8"�^5~/�ǣt}"YZ�~�Z����'�!<c�a�l5^76���=����^���Y��{������?eP�c�ͽ��G:���1?8�2I|���*�L�`N^��c��2���!�p�l�\���Y2������m��W}D��;���Ws>��1��W=q�0���R��]�^�{>,�ھ�	�|�� �U)[��z�y[,_�c_���:�r+�HT�7�| �#/��_���OD����B�'�η0s�"H3��zL{�I]LĻ�rH2B7���"���=o�<��������7z�-������;
Ek���Cг,�x�#۰�U�ύq�Odd�4��j?�۫3[N0ɑ�n�Nl�T?{�t?m�3G�2��іm�V>;�8���+S=r�p�q�t�ȝ�_M�Lo�y�߫�-�;���4���hD���3��$�vn�֬�ԉ�q��VX6�����