��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf��4Oᐢ��\���s���(���T��p򱯋��}�w�i�|�typ)4�eV߁�����o9�␬+$����lY0��S�6�ڪ�<�]�Wų���2�:wh�GHFN���Ҩ�*CC�`�CJV���py P�{Z�����a� �w��������V���ѠH���C��~CU/�Չ>�*8,̏��wU0ġ|������CWS�3�&Ạ'"�-y�e���b'�5�Օ\� ����Mnկg~��^dv�{)_v�g���}[���Y�B�O6�c�z��M�����1&dg�ps��~((�(��ȱ7����dN�f3�f¬U!){_̺�䕰�����S�.!I�_�.�۫'�0�	��l�>�o�F9�ß�Ed��j���<�Vo���m#,�Z �DWrA��� G�]�������X�],�T�ѽE�N���8'�KAu$��AAg��a&p���)
E�7���X��|.|9��Z�0uO�(O)"T�w�AR%ً��{�+��?J�e�#b����|9FK��h�K�K���;��(��+B�B�#�N��0�/�b���3��^LBL���¼۩�г���w��> �u%s��o������[�&���&�V&j!ӳ~���Rk��H`�t��D��+8�Z�1`s�8Ə��q�2~��o�= �j���xrI@��9�;1�+-!�U��<;�G�������{*��gL3���^��n�o���M�梁>=��ڊ��i��4Ǹ�,3ȡ�c����t �5����$� ��O��_���	�$�g�L�䟃�ga�������kȴ_�7�.!� 䃄%��v��G/1���K28��	�q����/��V�.����R�����qex{z6���v3��g�'& Y��\ �Y�l4M�qb����?��+��T0X|I$�>������C]$�2�8�����M�����n�2��L�ٞ����f���w���B�fmŵF�l��{`�����K+�d�� 9�Z<�҅����m�F0��j���G�8<y����i�l�w^q�#Pt�\��_V�Ґ$�čT�u#Ow^1�:��5$Ƿa΅mX�V����L�S'\��9
SnΆ��Ԧc\!'oqor��e�7Յ�#~	�_��p|�����8�!ҫ*Hdt�v�.�a���xnW�aWZi����������&�M����$���ΝP1�q	x�ݳ�8�iEE9���n=���L��Q�!�W���~I������>E!����uזg��ݭ?kb<��z�W`$ym�h"
f����X��㺞E-�Ȯ�Gb9!���,�r�C��Bg�}��q?�F�d.�x��%�.ݻοַ5xlҌԧW���X��jJ���R� ���L󸙰0E���4��҂A�j�j�h����yA2&��r��Tg��M]���kv�����3�>0˕���G2�I ���8�55�Q�f^T�5X3|��̊�N��5�ω�IuQ��?��1��e��	�j`���ZUZ�f8z���y�&��EsѲM����"Ѡ>~k*L'v�`�%�֤���ǌ��Q�
��!�f���]�俙�d� e���O��
X��쬲�&���r�f�n��C�{��c�[n�@�`2gu��C	�.a{�ESR����:��z�=�C���I�B�����*�:��Im
?���l�؉�F$���~m)��R��0��Ma�H�0�I�k��g �'=G~,��+���>.1/[��l`��Q,o��Ґ���u~��P~�ҏe�X���<9@���z���Îڋg�0�ގ?�IVP��P����-8�=�V��w�Fho��g�je�uٔ�]U�N]S��S5��W�&��{&�.8��l�|R
ca��2��`��oP���ݫn�UiH�+PC��)I)���+�����z����?mu��\�AB���v�����C<0m�-��(�h�]�ʶrS�1��ә���Z�_�M�ONe�$�g����n�9���;$%%OG���8�i���?�2�ڸ̩G�,�%{�z����4��AQ4���Y>�}�������B"�gƺp�=�����]���E�� �,-
4�`9nwJ��T���Q菢q�9i���1�CSߍ���ޝ_�ˑⱮ�	�y�q�����|*������L��Ú�du� &�3�&0{@�_��ZS��TU�q�!u�1�.q6A)��r\<7 t��񨚅�̨���DJ ���d�q$�S^b��E�m����^�͇o�;f����]�CռIw�3�dB$�jv늊�j�[�p���A?�"m3��/�r���ڄ21Z>Qn���QdA֢P��|���֢�� Q�2O�	{2+	��3�����<�Y�s���.�6-Iw1�;N��!�k��rZ�EO%��'A^�6������+U�����K�8���&,�8�\8���ߝ;��#V������?λl���x�d�F5_	]�v}�ӻ/��������v滘r�T}W-7�#�g�������o�}ީ�I�jGHU=J�e*��h�
,�=0�j�)vdY�c�7����;��\����I�\77�=��r�h{D���4gO��d��أQ�]D���f��%p,�Mh�o���/k���]��e�"W�<��%�|�m�8�)�"��!Ԗ�(j5�7��yW��k�x���o͉��UkrV�9=&�6��[z]:C�m����P�S/�D��y��`�kti�XL�7j��f̵���k+�R�n���	pW��\#ʫh`G�r�dҾ�iiSp+J�	c��kC'��W�� W��A`9�"en.K�X.�$������jУ+Ƹ�s��#C{�Ӫ-�F�_�Ced�mO��<|w����'�D�>�Kr���t��/A�GG誛��/�.U���ifqg�F��c�I}�K`=�(��U,������T����˵9��2r_\�h�N��=L=~���M&�G9R��H�s��(�_3.�����b�y!i��@�k��V�c��Gp/w��o�����x	��K|��'x�3��ά���e=9'�܁r�"R,9�k?�d��TI;��.��Z`o&}ì�4�<y��Q��Ѿ�gC^)<W�|�X\�X�Fv��"��/�6�jo�~_;k
^#����A\NC�D����_�f.ӈ�G��Ua@.���q�{�I��Rb����C���Ix~E1��k���5A��ܴ��3Zrj������9{�����D�S����Ĥ�����<~�p��l��h�����!����pݙȈ�"�|�p�\��oި��n������/&���]��i�C7z�:�fD�H�1�x���孄0�{�p���u`�)�)p�z�6	����	'�&���j�@T�/���!-0L�N�c�Kf�矃�5~�H�׷3$ic���܂��R�y��q谒c+��UᲗ�N�U5���d��RG���7��w��*��p�H�N�%���_��k��e��ȁ����1�v8�(;����{�YH$u�<-Ҷ�L���G���O�S�3��8����ju��3�tVՔGm=�=�|Q���Q�z*����=# ��m��Y�*'��W�ٽNo��.���4������g�y��Ѐ��yO]����g�;���
��@.�q�T,6�"0���T���fsy���u��B�6:����B	�3�P~�p<|�H���e<[���-O�r<��e*û_�菇���٥��y/LR���\LQω��W�0hO�Z�*��XS�6����I���U�*K:��4u�磊rq&|I�i �ӹF~�\��ZP�δ�0 ���zg����D�A*9]�Fon�-M�z5U��P8kߐl_�ǫG*�8<��Χ�����[�?\�E��IzMa�
]1��È	���/�w��dն�G��~�������e[lj?�l�i��Q��#��vd��n1�+q��(:�����/)q)��B��XG�"o�Q&b�qP�y��zXo͝B�6��~?�F�k�vSV�vc�Ex�$�� .f��
����:����i�>��o�W�T0k�i�7h���Yҟ�'��	�4琭�fe�<24���N/�{�sYc��J@C�ÎV�����9l����S ��{\���8�"��>U��}�m6�Wh���}�U,�'��A�OgN�*o𲶐J,.���'���@7k �~o��]yl��:k��z�l�Y8�9��^�Y[�Xh\Q��y	w�45O0Q�¬����W��<ڎ�b��$1�I���P�v�G��J,��ª�4�ˉ��R����(�ҟb���2@r�ب��V"�څg(����ӥ!����05�u���0���5�E�D�n�P�P�����RS%"i$�Бp����I�+�Ͻ{C�Ro2&�(۸�'|[���̅�jh!�xQE�%]�H	@%,�zʊ_T�����$�h�|ٷGLG,����SqV�6_ۄ,���Ca���tXL�q�4o2,d�}��;C\x�7�3�� � oM*�M� �0W��@�,%gak�3����@c�{�N�N~8�+�D-X0�g  �	�d��h�2V�z�G���%Z�Ce�O���3Z�����RM̾��ܶ���vmb͉e�>��%ʘo'� ��U���PG����G��w"�	D�[�F9�=o;K%Q1�fu�=�a�(es�����E^os���=��!3pVO���ȉYRG� 5&�;2���i'N���]����l�w�c���=�u�[u�L[�_q�W�w��W�qk����S��'I����w�����!8��J	�jK �+3K����2D�L���K��h�:�z֋�(+�Y�I����K�R��H���#p{m{<C��]��CjՎ��JVF���P`5r7֪`�7JK1pg��n<�?�闦��̹CN���*�Bk��z��6�
z9#�mU+m��tAlE��w}��4�'ĴvI�_�&�v��� ���(g�(��|������]'(�ʡ�D�ލ�<�Y�ݹ�}�i��k�Bcƛ�绳�q"��	��|��Dd!�Q���<h)I�(���.E�n�dÄ�x� ���E^���<�kL�����Q�_t� �7�
���b����x?s!4�=[!�5T�_9�d�1G4���9�]W,�K�ֆu|��ϡ�	�u$�M�_�jBD[�g�Ź	�ڿ��?D�RW`H���M�l�����-�x��9��*2�vH%7n�;����F�iL/���j�@T��4`0a��a�I&l��+�Ї$�	I���ˬ�M��D���w)\;�P�FB��g��20��rݗ�ڶ,�2��μ�c?��MF�*y�NYcץ��u�L_�������y:�?�$��ډM�l8;ab���K~���^n"`�P7r5�^�p�?�L��u�9�f4Ï��}�L�Ȃ�|�qw���l������u�|y��9�>hs1�R�����5^�Q�R����܇�q��!t}�������J���]�Z틢1������]!]C&�<�ahQiow�ɸY#�&~o��aު��P�Y���_�?����6G����zo��i\6-�)�|L�f3�D�(�uZf���E�N��\L �͞�&�U�r}�>F
toN�'�˛�?Op��BLf��&�d\쬦RN��X Oӝ�~\Y	և1R>n���Ծ)�~2����h����e��ɄG@隺�&h��1d!/�����{��iG����A���ކ�#���&,�(�凯�V�~�?jbr34�^�!i�=/�>%��6��,��i	Ued��p��$�+*�H���b����K�'��m1̐�jcR8�ܯ�ݝ�<0?�i�:�1�U��l���G�Aӣh��AZ�J�⽧eb�R���Ive�1�Ŋ��*G�zgD �
���u�����j1��a���0"�S3��Ҟt�M���{n�!��mq��2-�(c���O02t�X��w�j�7����77�*���5�X=��I4|��o��:�����\���4T��,7��_E4IP\�aX���Dڟmp��K���J��@c�	����UD<�;+�{�X�ve�a(�	Q�$�M=M�k�q�į<�v��>l���^+�[r�e�2Čw��i3�/���ߊ*Z�G�㿣��X�2�����U�|r@~��b?�odЕ�<�c�E��������9βīx|�q��;�892��X]r�J���Y�X;7�7C^�dɄ1�x
�=��jFst��#<�/ȡ1+�$�<�k�3��ά�T�	EҕzK���-�Lk^ ڙ��
�@�����@W��c��8�9�C�|��#��mL�e�WA��J��Z��}�!m����:�����k�h�r�;G::JOY���_�O~@S[��s�oA-\c���tMkfy��O�4*����_�[���U�`���S�G���[v��׶W�-*�
͌�|�l�!���{X�@7O����@׷�����sMX�DQ�������l���D� k(	�<M�D�u����ܨC�3�ϸ��@'d���V�aa����|��ճ������?�p�Ĳ�5	Q{R�������uZ�~.rn� ��6������Ӽ��f��|����k�>��?�j��	����5S�y��l���#�U���Ǌ�i0�\�L᭼������TC*P��܆���,Ú�]�`Fn��5ͫ �4.	�0&�*�~����"�z��+,�������u� H���5����v�[h��{�R~@걠6�4���I��m/����o�fD��r�]5f�6r9�o�۶y�3���_��w~Wi�5`�\K�O�	�U��)b �i�������en����݉�B�#,׎�Q�$��e���YJ*�H݉�͌��_�I��ɮ�*���t�\}�!Y��
���]oՙ8.�S�1�C��1%b¯�#�y&�^�1�J�|�R��YS��Id@3)]�vt|ʛ���g�	.A䃺c�����e����h@+T��&�M������R�k���IF���Н*bd6]�b!�ҙE �Ɨ[�~s�,y��U���{وU�<e@���6G�B�߈%	M���!|�E����M-4���v�}*u��_�����_�J}�d[������C��fr������Q�3ˍ��n�T���Y,��T)��='�%�_��*�Nβ�ĥ��%W�J��{!���'�ɼ�"��#<c�Gg9zl�[�
m�����Q��ӑ\BEx�+����揗L`��V��� c��{�wb|�xR_!([�`WP`��_`j�<G~�0XѬ�\s�K�Jcht��e��!?}���gZ4��.`>#�pDM�ǜ:��EI�nq�F+��(���+4;��XlN]�-/���si����	u�0��2O^WǍ#���Ƿ�5k8/�#�lC�w7|w�
T�`���4 lVg���~#4���0��K7�x�8���>E�j$C{��T�~�ɜ�[���]����PQfB&������*O_#��̍�8Y�PQ��Ħ�ݡ%��PX��Q�$npf���v�"�Y1eC<���k��O�	����FK�=CU�U4��� '� �j�q>�~�����φ���L�����s�*1�2K;��5�XU�����֛�z#p��}孺�R60.����8�|1�C����蚐
�4�4�Ne���������ư��Bu_i�]A:�'����lӠ���'��,"�c��N�Y7�ބζ��P�F�P�������,�M�4Ա� ��X�#�C�f���HFuD�.;&"dMe?���,�Lcm"�a{�E�%���<f)�:
��"��3��7S�7ܰ��x��0��6%��B��J��M�׭�u-�u�ɟR.͍*���y�������������I?(}�8Ĳx���ò`9#�����������4��Ш4�_p2����������'ݏ��mP>=��;:J�aDKtm�
|�@�/b������-�c���:���=f,�x�X�2�$ݼ�y���A~D�r���[N����*��쁚+D���������6#��o^�cO�+����ǘ�r�td�����C�x7�Bbu3?����r0_�p
ZF��9�>oK:����{ݧ�X�Ь�j&E\�qkAy,�v����:C����Fx�-ɑQΞ��
��F�WX�
41��z���+�&`%0��D8�� �H�ɉߩcĭ4�ڍ����S������'4 ez�|����Y����I��S��c�/�p�
�D��o�Z�5�(7�J;��Gg�ۤ9�(s7�&���-��ݞ�S�u�;�d�^����G�І�k�~t\5"Th���v3��$Q��^�ro?�/Q1F���|�~㟲�����n{�c%E-�?��d����mͮ0�%!���m��.�Xږ��Qp�����@#�I��������c�
�����t���)�޼�Bf8�jj���򪴾R��~�T��bR,�|��գ)�q.�e��ml�`�B��M[�eߤ��<[.�=x���F��È��x�_�B1�V�%t�G����,��T{���LD	:�x���1t^��'+��i�ϰ2��Ͻ7ξw�jz�<���ss�a�0�Ɏt�ge�u�U�����^�L��)W�h䰞�ԗ�����ݑ���-��ț�_����Zr�g_����H?�P�[�Z]*	��j��I/���R����㘑A�:l=[���~�O_g�ZX/C��ȇ=(�$N�?�f�`���C��ƞ^��X��0MQ�ϧ�<�Y~������>�*WS����_y�u��#���n���Pa,at�.�����Q����[(|:�l�#���Xl�k?�Y4ˌ�*���|,CT�&�j2,�h_�K���g�#��v/t�&�	Z2��vw0-�wx�7E8�\�Ѹ}Jc�����С|�Ǳyw��
C;�������H�wq������ՅK�0��p[qԭ#O*n"�N��=֚�
��o��s�3�ȁ�S��|������6	���_wڮ��5�����G	�q'u�HQ�5��} �+)���W��dx2ZE���] ���=Y���(z�ډ)̲DST`O��х���*�vl��!f��.B��<:vU�����b_eOV�^�<�3��NL��(k��*N����Aث�>X��Y��Z�)X,�Anl�{@H�^�58�2ֿ3�x��Fr�0L6ʍ�9���Å����͋5���]��][l{^E��h�{ s?_�=,���>��|� ��g�w�K�~]�:���O���q|�Aۈ���%3�*IL$���za2�ꅲz���mޙ}���z�BjM�v;��a+���6�
ȭ����*�F�?aɬh�F��"�k�4<����@���B�\�&��fw!�W�cm�W�X�JZ#7<�\�C���2�K�fg���['����G*�sce!E�zg͊�U��t�ս�B�h�q�J	��'~1
Z��f��(4�12�D���`�67��Ȅ�@�*�W۲1� �m.��ui�> �0 �To"�����H���V�8;�XCi�	�	4��Blь���,L˛�F�ұX}<��lf��='�mm����E����R�>|ON6U����������-Z_. ���%O�$M���A\K���՗Ƈ�lnR�ۧ��-u�\�>׻��Hs>�3����������b�6�%���y�c��1�AU�a҅N1�r��}`��j�������~S$���B0<�8`�1j�*�>Jk�cM!���H��}CT4���*�=�L��+MH_꾃��D|�w�rmw�w$~��-J�́p��m%���4���qI˖Ly�H��Nn�}#M��;@�$Q7���AoT�YS��� �Kr� ���N�y����i�4M_�lI����D��� ���[|�XW�dٳdLi��,�o��k$��`pZc�I�g����;���l\)PB�ֱΘ�1]=#)(*��"�b@��'Y��P����p%�y�>'���$�U��ad`�L3��o�;���w��b��T6�]�������%�3��$�(�]fT-�J!�@����\�aj��f��=;a0�D��R��W�.���_�q:��;5��j\g�����J$/��w��.�4��"�(f`�Ϝ�������ꠑ{��s-E��Uo�}p}��ݢ�{i^Ŧ*�A�N�|}�d|�9��UR{+@x^?'��@_�V`<����N�K\�N0Ԛ��D��K��ȩ���w6���&�?zpt�������=X��D����rgK��Z��oLGbf��� vG��l/��4^���B#ā��u�y<ÂtH�x����&ϫ�>V�:+��΋#P�����f�ԡ���q^���L=L����a�Uxg/vTva{{=���vυ����L�b��oi[;��Ab�{Q�CO�p̙��	[X�
������_�k:�X=��2��:ȣ�X�X����2w�j���Y�+>��P:�����l���(��)��:�<q��Q���)�Z�Br�qk�I��;I��8�C0X�]��{�&�`oa"�K���&�u9��l�R��)����dl��q��%�)榹�S`G{H7��_�و
N��j�n���Q�;�p�0Θ�y��L�_�U{���$ܲ�rwӜLH��fe��cr[��-���~Ipǽ:�Y��Ԫg���������ɝ��:~�[���.<I�n���%V�]b�(��[�ix�͌U�W����o�-���E�#ܙL;gM��@?:�*�È7*x)�b`xV.�~��uO��w�v1Co`K[g�%O����w�3�������c.�s�TFb4�8|eJ��,>��� 9더^�/��<�L�{7��k�_=���w�#9;ud!���ɢ=� ���U�jFu�4 �D%��[�?��{�¸&a�w��VLg.�Q}�D-@EDft#0vڼ������_���n#Fl��
H"'s��:pD"�f�^pN���c5f̟�ڗ����̠I�@��n���{����A+AW���� r!�׭�2m�{�����y�ڀ��9lpTF�Cl��[��~ۭ� �/Dk�P�7j���E���I���G�0�l��wL��2���h�H�`A���QB����b�0���b�DzO������x5i}��,���Ahϼ?J|"�.�3�H�,�[�+����@�\�:�c,��ޭ�����[�x�H��[�� ��X��~��-lٱ��䲖y���zG�$:Q���j0�,mW$P? �$�
��)���=��S`��S����<(v=�X���LdG9s��=��
�x�M^���no��=��s�V��Jn�*h��p�k��[�m���88�z���e��t*����3��B��3�����(���Kv�z�T�i��vp�Bg���*2Bh)�)�j٪&x3��/�]cU:V�}�J���%�MKo8�4qh�	PW�̒�Uאm,���*~�����S�ܙ�?�����.���ҟ��=����c����0h<^��s����ʭymz�����E�ܢ� �1H��J�t9��d��#TS�b��-@�ץ�/, 2x�k*`>����"ߦK�3c4B�9�:����ա��Q�a�E���K��^u���C:/���5��5/%ٍ���>6��� ڵOg0�3��)�7͙5q��)��l9����ͅaے;�(�J(Y`K�&);$��6e�
R��N�r����ev�3��ǗP�k>�5��0�7��oSp�jY�蓉�H����od��s���"��]P�����|�(a��)�:�tFW�><�5+&(��;��=0�Wv�[���(��E�V��n�H�TM�()廑�� �7·p�$���&�f$���}�P�9�c�&��h	�ʠ+3���;�q÷` �}�&h�hw�?�GD<enk7�`�o��vE�"6e=���@㲲:��燀F�2<���A�V��ݏc^A:����k�O�����8,��Q���'�,��|y-(R$�#)p��\f*sKzJ�1�MXf!+�F�0�5�7�]�k��9j��@�YكO�'�v0`C��4���5%x��a7~�y�KB� �!:�s���&���R8��aMþ]9�#�r�%�Q��,��/����`���f�����b�3��g�D���_9@��� ����K��r'Y����>3CIN�Z��*
��)���fΘS�S�I-!Xa�JN����`���}�n�B��x$�o�C:����k���s�8�COH�'�-3���׌<z�@����l�h� J����h~�l��0H��z˻��0�_�Y��tc��d�����+��97h��2^\�	2w�>��
��q��>������62l��.Pr��H��>l|����e�yךwd���Ց5`�.�uiF����]���$���[<M�n�7t�=����ן>�Ӫ��(�=��k���0VaV���~x�?�S\��^xJG�@�5MW��������*�&�� �a�w#3��0P4u��{�vxY"�3/Ѩj	Kp��Nk�Ʊ��C��>}+Lz�v��x�o$5�_�j�����&�WXg�jj�25���wͳ��L��\%p!�T���S��>�9]�B$5kǈx|�� ��߅-�k�7�S���8�;9��U��>�B#��ؽ"|o��YB�h�O�V�����GZ�F�A�bfٻ��S�O���@:+��n-(@�U|mˢη���+l�h'"��yE�d��9�
ش>��������B�=���;����@�$�p�e�8�8c�E`�k��;~�hor�ДB�p��0�(��v�f���Eצ
���ES&s�44�L�3��Z�����@1���}Y9��c������9���;.�MXP�S����d�-Ӳ<w�s�� N��En��ک8��{���I���f���.�vr����cLsXTjҏ��;_����N~Q��u�a��4��%eۘ��ʮ��I�F�d��$�`I[TO�,�}�3	^
'�cNOn��?3W�2��e��e��@	�5*K,&�x�N��?����4�訆$H����y�硁Cd��d�qu���@a崸�"{�*o'��п+SV6�6z���x\�c)� ����\>��k�o�M�>r5}MF�dG��p�(?x�| {Jyx�F���H��!��6�AJ?��h_�
�7K`l��v&53��Ɗ9e���YX2���<�� $�����E��P�@�O/�����޵�[��zTA`K�K��{�@����B��W��u���c�F�`~�֡ϲ�*�ۚt�V6o����1�eMU�7s5Eu�����8(��ν�����0M+y�-� NV�Jq����6�rR��8֚7�FĶ��Ɯ�Y��5��N�}��``��yj*�k
*��P�m�Ʋs�>G��E�I�BE
�;���j���a{X�OZ���|�̦���)���L#. �3TE�r���$*�y#�g��<_Zz0���P��&��Q�_S0����aAm�3�V�o���Jg�ƎEB���}�|�X��){�x��梌�6���j���p�S�~��x��6��T�硅- �z�"0W�k�.^����cp�~zK�_�j5W���eqo�%����'_f���	�k#��2�+���
�Ssj	��-z������<sE�u�ǥ|wS�����@��L-a���:�(���J� �$:\����_�p��6.
�\�p��n*��s����a�*��$2�*`6V3,%�pҊ��![�&Ҥv�s/���r�߅��������~����{b񣃣���qv�FY�C ^�P�f������%��%��h�F� Y�V%����Z�h�0�DF�d���NжS���]��b^�l�0�u�^y��d�g��o�o��s~�Y$cjԬj��I��
y��!kv���5���ek~�e�{�����x����ȳ9 7~b���^��j�y9�;��nB�Pk���1i���o�&3�G��A"4�^RsM*��o%�m�P>��AͶ(&!�"m���cz�z?Ԃr��&�lU��x^��8ij���i<J�����$�yIk���d@��������l��J�O�6||f�7j^���a^�c�s�3��Lم�/��6�U��uk�b�-�
�?��(ݜ�}rօC��v�͐F!)�"8��%KG�\�Ⴞ��O�6΅�!J���%n���x]��s�ʆ>��	^�gz�-��B�Nl�a�!߭�6�N��`�E�����o� `o�ﳃ�@Ę�x�h�W!PĤ#�V�4��.k Gi����e�%�:��;$w��|Zt	{��[r�Ud��V���K�x�~���[�8m���?�l��ң0�2l�����[x����vf�>ԅYs�ϳS�ؽ��/$j�28"p���	Tt�W�D�RvPi��=�p�=�^�#�
�����>�X�h,�Z�D:7��H�8!��n��Q�W�a�D6�5@:a������!,1��7՛��8��R�yi�/x���Rw뽼R�&�_�/�ų��v�xAD#��"i��hqT�!�hNh���`��@�1�� �4�)|�M�]sv�T���m�H�)*�蠷g�E�v��u�&�裏�)�cT���q�'�|���� �&a�/�.�v �?
�FE�&ȯ�,�
o�<�Z����G�Qrd\��ܣ��屡/��j"�W���y�n�!į0^���/q0�b|��C���?�:,slh����7CE��`:e�����d�������h�"��s���ƽmB�ƪ0E�����-��f��	�b �,v�ˏ�^Pڅ��I�-��P�a�W
q�O���6O���e*��S�먄�6�uM�!��u3f�E>8dUaLR/�����_p��Y�jI�Y�UP��
��򪡇�&�O�}:>%Cw$#�����)�`Æ{��)D,��<�=��϶n�HȽ��s��K���ӆҠ�����*&�qK!=��w�S_����"%M0a7��;t�����b�]�+����a���H\�:���JWƉ5>��G�f!���d��Э�b�,�i�qɛgz�[C��P}�Zu#�H�G}b]���]Ɉ�g��B_m�]��B��ڍ�SQd�R|��1��qF1M�pq����=6w�{�{�52Z��]�6���|M��s�>7i����a��h�*ў^)5����0���Q�Eovk}=@9�J�Hm����>�l�@�{���i�e���h�/��ٶw�AB���\$���V�g�6�C�����<y���s\���(��E:HRB8��9eQ'�%�����\	�%�Գ��8�b���b�>?��)s��?�\,֬� �20�ᙩ �9�� $��1A�OjBG�����l0|����&>?�$�fe��qc\��j1K�U��eV��-{���O15���"  UO��>�S=i߈��j��w�p.B��^J�K�>=1�?0jת9
���{�Oi�b���e�C��`�^�w�Y@�X�a�4���GV���[9Mb��D�]��J/"��(V�tx��� �!C���h��Th�h��'6�����{|��-;Ia�����Vw�0�H�Lp�����"��k�t�?��y,Q��)w������ȣ�?Ji|4w|ΦB%��T�,�)7��('�%��X`ۋ��-�9��01oӝm����M#ě�w� �MS~�a�ׄ���1Z+�ٸ����0�&��(��}c5���h9����t.�����j8<`P�$�j�`H��]Mˍ1p#�I҈�Fv��5H�}��(8^�Z�TV��̐,W��#�Cw���$&�+�L�F��k���k_H�*�щ|� /��E�/��Jn4�����~#�ގ7Ǐ��r�u�do!d�#��ӗ�B>��P�GR�-��x=�t-�I�^�-S*	-��m��CXg��{�W`)�A5x�W'�cgD=���M(��Yb����}u8pd���dM�i�j�ne���`������R_y���=�JxO���MDl�䄍�Ǻ��_�h��I��lB�	s��΍�h"�!�tN� 
gk�X?���ZUR�����&�#T��}}L�C%s�9Cw�U�{?��G��S0Ȇt��\5(I��Y2~�@��8uW| x6	kD�:��l��:!�����+�s���^N3����M���}��Rtq���ˋ�]jD4��CyZ+�O�/�b��&��`� Φ�_�N�}�L�QX2w0���%� ����=4:��r�\�c�0�@K��^x�i%W�/�[��X��[BٽU����4
�Jd}O����,���މ%!}��T���a���#�A
KQ�N�p!�#֧=��/9Ld�	��ܖ���W���4�!�zC;�i���aڇD�o�Gt$K�0b��v�Z��t��6��Ϙ�PhQ����B����-��}��L�vIk<8r[:v(?�!�������7�?�
Y&(���[T��8?�����F��i5h��xZ�)
��!�fu�6�P#>�3���|�(�^�Ҫ�V� �� �L�-ϒQ]����uI�*�@���c�-���o�O����-�T;�g����@�ȵ��m�Aܾ�j�u��r���3z��ӟꁍ|��B��LQ|NA�g�؇�G̿�"_�(=���N��x^s�8>et,�"0|��!�Ӱyn�6Ŕ�Y�|7�U=|�i#�E3�ʛm�,|D8���9���/�ϴ<h⯄�	Qv��WU˘��6�`�o��_���9L<�]+eB����d�t����K��yɒ1��`kU�*�c-[
�/�H �z^�&:c�;sa. ����g��H�1�Q����:)BS��UR7�M�M��q������L��sTi��@����U>��4屛i�ã�;xWq�������O}����}F� ���
��*�벗G��z���?�q��f����Đ�	�x�1