��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|e����M`p��L}a�1���mq�ݭ
�:ث+�n���M�B��7�jŽ+�"��Kk��։`��X�z�1�i��J���e��4Z5���C�&�⒇L��禭�c.Ę���\��9�^�+����Ƈ!6A������MΘ���{��1��c��P��w�+�rQv�r Ź�o�i5�[���,_�J!�9�ČL��+�xDM��4�j���ʛ��h�dY���1V�������+:�/������_��x8�=e���?ƭ�øҸU'J�(�#V��XyQ�D�z�Z!O��tr�����$rH&���7��pWEf���~����Q�+�$���:��WN6f;T���3��'BMD��sAPƿ]���(S���T�jX���;��	ib�D��	�l��hVR Ͷ�ed
D�P 	86Hq��L�t`1v�jR1N�u�	�
���c�9b5�춾�[��if���xG�y�WY�C=+/�O���H�%;Suy��N`��4�'��q�ɂl��/��`]�O|�m��?�q�2���B�F{ef�9*Z�+�CG�i'�x4y��Ԙ��W��������@�IP�z&�$���0l��~	F�:�H��^(��\D�EEɚ�-�����U�O)ʃ�v�r�!ޗon@�PT���UK�OT+��[�o�ci�2
)�i���;UW��[.��,2gơ�6��b�q�⓾��844���]��3��4`�,@����Hu��(�h�E}��x����I����eb�*� ڪɵ�6�D�@w�l�X�6��Lm�8�w�q���zG񮞾6|����HG'�!~ӈ�tT'�o��2(c1fj��Q@C��}M{!Uo���2�- ٪hB�m��Qd���k<��A��N`�ˆ�m�j���lﲤ5���L���h}�2������B/��/m�̾��P�E�&c��*����K��|(j��)9�ԓ'b��0C'����� �"�fK��d��~my�}�ׯ.-�T��*�Ԡ�f?����Q��0`��9���p[1
�8�j�)K�m�K�i��#�a����%͜���;��-Q]�6)�Q�o�p�_�PÌF$BQ�DQ#d+��a������g�]?�dŖ�&/I�ےz��MT�p�C��!�U��F،�p?%�c��6`�4o���b�5���Vϓ��Wß�,�rh.YW�ԩ9�6�'V
)��J+��RZ���0�e��_����/�"��r՚���P�r�Dcq��#3Q��EN�Ra���@ʻ7S�o�*�Jr�5�D��I^&c\��0^-��Q�������������P�"�O:��C�7��sH�$!Sb����#�-�æ�{�=tgc�a?��У�{A;d]�/`�Ts0>�f��ۊPf�'�\��]�):���-k)���~D��op�e��\(r\?����~K}�����k�� H�;a���2K����3����O3f_w��2�/z�Ċ,vG�<�0?B��f�a�?���u�Cq���jF�@u6Q�3�c��2���,���ө�ˬ�Y$֨�^�AVNa �l$X��$p8]��f#���"�M��P��[��_aa�4R�ĩ��@n����h*F�zɠ�4�?�<Gʳ��D*�0��<Y��~32B:�=�P�C\�U��^����*
�rԫN�h2m��3f��ɲ��yI
v�0���~�P�[+ ��yb�9�)��i�Y���Y�J���}�M�����M�w�W��l���l���k-c�y��?����E��_�R����e��1�N"�����ohfT�HM
����[�����qbUF#�̾�&�ތ���<��!I��9ࡩ��3�lPh��# �<#C8ʽp������>Y��Pz�et���6�W�?�F���V��.Fo,A�pG!�x9����H�"��G��1����t�2���r��[�vQ@�eIC��+m���^�_����ğrv(ե�슅y#��ůη� m�o��i��� �C�5M.J�b5Y��
3R��;�Q㔏.�E�|���λ����ظbQ�Aʛh%�p�š�]��5�����<������i��U$F�b��H3\�}���q�n9*�A��U�o$�S+�2�B�B#�	.����Ά�hF2*��#��1�n�ˢ/{�椷�$R����O�X�ϑ0΋�8O6�nVe�8ׁ��MOq��@��h,"x�\�����,}y��J˯2�� �w�0$�-�v��Ό�A���s�YXǙ��	ۙC�䭝g�,��P`6k�ox[�@�b����4i���1Wg$���i֙��|�������$(�:Ț	:�[\!Q��WǾ�V/��%-\ӀS纍�I-i�أ N�> ����eLO�����oV�E�斜{�Ga���aױ ����@.���V����_�@�?�#��F� ������`lA�ajlTf����C#�Y�m���~� �c½y���
To�
�����ӕ��i� �q��������̽ͩy���S�Z�Y�(�'Ir�� ]�s��W�}ž�X���X�6$�����w�V�&��!pv�)֘�b�n*�F��������4z��0�Ň#�e��+�x>��K� `dM�l�U�|[������J��`s����+$i��.�{�s9�HY��ؒ�3��q�]�/�d�N��m��]��������l��P�7�`���8�oA�������*��B�-�ٔ�p��e]ȼͦD�闲���8��Q�y��Q��(���0}�an�zX�a�А�c�t��i�WGA��႓�7�33t"g�`�a�Q���r1�{�iJ����Ѿ*D�0��|�<~ɽ��xR��O���d�?�<�'U/*Ί�#��a�]�\�Z��v��#��|���^��ܾz"r>[��`�8³���_�;��h���X*��g��<7,��@�,�<��>�]���KYܣ4��u�^�i�q�K�[�^H��qr�hG�n��[�8�xu�(v[/�J�
Ô����sw��ǫj���^��u�7p�qo����[�vbW�~�*��m_��O����!�>���@S�o��J���1|�3;.0n��EB
�U찬� �`�,��.��W�z��\��i7%�r=q_Ƕ!g$�qIz�T���J�����)�D8P�8S�B��O���5����VN8	i������N=Тȫ��[��D��T	���L�	�y��-� \���r6G7p��F�R�)����fgy�:ioY1�D&��'�[䓕�A��WL�p�:������Pz���lE1���Udd9n�=vU�-�i��+|ASQS"�o;g�'�PpJ긡�M�V>��{XH���D��ITؕ�<��2P��Ӏcm|ѝ/�ͭ�h�lƣލ*i��s汾@d��.�Zsa#��Jq�O0�J4�T@�J�%¯J����3�ٚ�F1u��v�+Y���"�V����V��aL4q ��f�!��	;�F�Z�����:��ձ�N��8@�l ��K��uv���$H++�@+���u��%�?�3�T����CLX�U c_"��R'�.J0�c���N8��kk�n�Ri毞�J�yĿG����Q�,�w��s�aYZt8ב�	��aZ�?g3eX�T���х��F�wM����+�n<%r.S��9:��ŭ	�-�/�`-�j�#N��D���2��p����q���	�b>�@i���2ADX��SLW�'��������)rIc+�����k��m[�^e[1�7��1��g]#I�
�Wir����7sx�ݹ��T�c��ߪ4�a-�4�N�6ηϔ��#|���wFP�B��d��;������Oq�N�-C��n�J;o>�$.�)3q�B�������w�+"��yz�BC��w��_���Q����|FM��8P52F�Y��� �!��ӄQ�T宊y��N�&�<�����nkZc�]�̲"=�Rt�5���$������mW4��{'m�ɼ�B�4��驐 sY�T^�g��VE��q�Q��EOζ���!�i=��a��;��ru��!�-�DMѿ梕,cf��S�9�a�Yj�F�p1n�N��,p)\oO�a�j�gʃh�@�]�Wͦ�%{�rNE~��--D]�=�Vp����
�ܪ�;kݗ�oW�C��I_+K�k�L���m:&7X��YU!�j�>�"b�������)�C��qX0�qi�_>$���T��rp[�B[�5�sS�W�3�����+3��c����<%���b��%t���w*󀧱��d�n���w���(��y\gs�c/_�r;��J�J�Kʺ�JQ�ip!q��)fo�� �-�jODļ�S7W�e�`^�ijv���������OX�D]	��'�9N���	�;,s����7~A�[X�h�!lLhn�E�br�/dq�@8�(���7�75x:�0}�G�F�*�t�u7�5~�s<�,GF���%IJ��/��#:�ox�Ir�����	�za9Æ��g8vh��g
�U�MjRO�=�:��.���å����`��5�8���m�Nn�@�9��g�jr�����R��~�"�O�9Kwh�8�w��NW�4L�a���W�.'��=2;^	�����k��Yz��G�[wk/��ޚ�;�L�̰T~�~��~\�J��W�����͵�[E�<)���Ϟ�E��L0����$M�M��Z�Ći��9Qʎ� ��XE=�މ�ELtm�r/{�������|�؋��S��-8�/^A��o���͔�Z]o��F��w͈"J�<Ո�Φ1�ĆGI��z�bN��|e�񑣤6�x��\Z��9�)�ڹ͠�� �q�D-	�_���Audęb���ƚO ��c6��B��3�ID�_^���tQ�n/N����ȑ��r\����1>.�7T�'��^�_��o�3i��	+84>�6�[O�a'��>n�y/`E����5�k�FZeeCo�Ͻ��!�Ӏ]�~-�Ll{'����6�=HX̧��R�2jXI�4$�"5��9*��e���hd���Ɔ�d�P�7r�73̸G<S &��.�Z�_����?��2��2��K����c1�OL�J�&�,Ls��缱NS}O�;G+R��3Pcvo�wt���v�fQv'�t�j]��"ڽ�`�9D�����
_��A`��1!��f;��A~��Y�.�M���Q9�8VUX�&C���Y_]U�#�s�#E���oEܻ�H�ZW�]���t	ra9D����̥���1ǆ����U�HJ��<L�����_Q������o�u+wt��1�q~��=�Tj�w���1Mwt?Lzc�2o�*8�Wcc��wk<���nd�r`��~M��1L=���z���yh�[D�zV���7 Y�:���7��H0Ė6O����X1\��}�]�l@頍鲗{J�1�=2o���^m�G�ݴj�A;�j���E��}"�WҞf�ol 1�M@�6ʡQ�)#�0>f� ��ӝ�aGz��L{�>������^\
D�0 {�"�� E��%/���>�M�r���/�頧���<�}[/ձ��)�6�	��!�������ǩ�����o��3g���K���Q�|��]S���"���4��S�A�|<�z�
�`�MZ�R���@��p�Bw�˖m� u�>c�\�����)��8�ݳɅ�z�ɩ]����2�C��Y�3���?ϖ(��辝:�������\��נ���78A(��+�70BU�6��\N9ƕ��U�Yr.�h�����[���6�s���)��t:����P�,lY ��㮫-�N�jqu5K*mo\R���M�u��.My�r�`f�#��kVl�v�������N��pG�f�r^��g�����*zA;�����%ɟ�+I�Y^G�Yҙğ<�_ȯ���U�f�\�v���~y�B@���P5챆Qn��\ի��Cf|!Ep�
dwl'� +k��ː�ĺ��x���s+��^1��.:�눤��R�3߽��!1������ ���,���i�H���?ԩ�B<a�9���+ml��6��9~�w)�ӕ�?��|'a��^&R��^��Sb�\��b_�~Ͻ2������U5��_��8�m��V�5���\��qUP�oE�]�%U̏�PЉ��t?���,���nw:[J�S>a��B��!�'��{�,[�1	S\c���X�������F�� v;06a�hoj�]��	\Ο�(��jIo��(��H��1?�s��K�y��)�b✥o���V^N��b��� 3i�KC�Q܈����y�.ə�>0��o��}��w����SDH��8�Zj.����3�>�2��b�*O�/��×�V���	R��ANt��Zd4ĺ6�[�ؿ����H�)�wWK����͈K֜�_��z��?�_�9�'�qG�$��.��K�P9|$*�KmVZ�m�jw!���=�U�Ke�+>6��}��A��Hঞ|>�i��"0\͹ P ����-B�`R��=��ow������\� z6�W���)a��}�-ɲ�ཫ3�x�vb
�T�ޞ6�Ⱦ_3ka�����M��w����Җq�R���]��e�򁁂�I~�	-VJ��8�4��ه=���?�.CRx�M{y����ao�:�+R��E��S�!�W;��
Tt�8t�g�z��jGU!���i��kN��/)"r��R����=<��<��#������e|
�\;���Z��|��t*~dO��n�|�I���1C�W"Y|�#`�h�>9������T�M�j·��c
�)lD�&�nΜom�r�$��&�И�ɲ�)2���vn��yܶn�ǝE�6d7�s�^9O�._��L�Y/�����L0ژ�ї��ި����Բ۳/����\7�1��y3d��PrI�t��?$Y�
	��4��p�ӽkU\#Zx�l1�m�?tzb�J�#�=Z�񾻯��J�.�N�NTF�3�����^��0�yn���3 �\��1���S�%�����gA�c����*o�A;���$�!�9���g@�������}c��r}G��N�	|=�*��]�*��8^Qw�ğ�K�9�9��E�����T�@[�u�!����������P��o�p����>��`5��9^��03���g�V>�ΰqu�w94���q�_����=�c�Aܾ{���9��Ũ[$���\��a��9S|�'N�ؘ�?��2�V6���m4*����k����n��_y�,�{p.�{��AO�6�U�D7�{p��^������z��A��B�;R��r/��YAzF�j����/�+Fal0����v�ER��[7�Vg�q@���^�h�m�UA^O臚-�V�����L�S!�9�Z;<�4F	��%�K
D;+����B���x��4�͓���1+S�)�cwމ\Nj��(�����P:�Fe�@k%��M�b[O�ͽWt��������Y�6I����s�����&��6�ƹA�xt<�>��Vh������"����iǳ�0,�k���Vپ��a��.�}x�'8�RTG-�������ݔ���_?PLA]�{��ۖ�}����GY�&,�c�Q�F@l(OJ�1[w!�XBT�g~c+��1e���� ����s]U/�i ~F����h��G1���`�r��/������R_N�.�o"��Tyt��J)���]�ܸUbZWw�ö���\ܵo��cH܄�����PlS�x��3��va�G_���f��xzF$2W��1�E�Kts��Ҫ1]\R�����eC�$�1�	+Hhf�+G(8��ݟs־�K/��V�?��h=(�i��a{T��b�9�Zʶ	M���e��K�#V�AُcG
[�F����}�.������Ϟ�X@wM�bC/��J	7'ի��L�H�_�t��uƺC `?���S�(0ۑ��S�0�x|h�b��B:�kr���7s�	�B݄�ГK��m�n�sKΨ�<��(5� Kn�kw�1Kq#BĘ�>7jD�	Ād9�.�`a����� <\�GfL���`e���oϩ��n;��N��{�)1�v�4E�c�P��I��\��zeNI��VC�\�C&��k�a�W��"3��#�`�ס����8!|�f�\��rd-A��3^k~X(��[zt��O\���>)������z->�Hh�:f�:1��C(�>#�ae+3�XQ�$F����J>%�Z�ȇ.7d����i+�O���h���X贰c-!K�ض���m'��.��_?[���T�n�����G��w���h(�?ov��]���,Ɨ[��2�;`�UF�@���� ��!�s0���Gs��5<%蝖*�#�,�U�7h�2�S�ו�����YC��g�%�$1�!�:W�6�������8{��\K\H.^H��s%�Ӹ�[�3�����g�@�)}uo�5�JA	E����V��-���YHg�Du����@!�[�����\Ck�����ט1�Y�&ª��Ǯ�F�׈��e&zN�=����ҳ}�T�9��/�+���X77�wic����D�54�v����@v�v�_L}Q�w�o��Yy��z����j>�������bIЮH������qV	��]gq1=�m��\>>T��I���ƺ!�r��\�W@dP����tm6��Q�Y^A���w?���ľ���L��T��
 ��&Un�?⪧�r^���3Y��c�㗴���6���cB˚�G��Ң��𩆯`�Y|�B<q��iҴ�K���5y:��rB�ر~���ض��@�C�0
GX����c n�U��N����f&��Kx?��p�^@��|9i�q&�zu<�x�,�K>��
Қ��y��Y�(G'�V�t+3�	�K��d�����5�i��ZV�ǽ �nqga��=�FT�c6�/���ζO�~��GXN��)�1[��{����^��虃I)��ƹ�\O� EH��S���?�5^RE'���5��u�j�1ϛ��!8bF�,$ea<n�t��"3�"��{:�xބ�m}�V�F��&8�<�������ʾ=�󜥃0 {�F`%hJhd��˵s�Rfk�H�B̏Â�=�	&i`���W�V��ߠf��0�I�`�M����@P(�У�(�O9���GӉ�]�	N#�P�M����i#Di͌�\����h�4d J���l6Z�_�8Yѽ������­�v�~�ɳs�%�L�"�2�^������v�Qί)!$��#���x_k��B���s�{�~!keiH� ��O"�dXj=�F��d��L~(bL���&l6�Qt�g0]�d�`e�u2���[lƼ<�kύf���R�8g�g6�F����k��L�7X��a'D��9����x�`�O��]���$������j���f��YKԃ��vS���,Й0ZUv���t�.+��}u���E��9��1�Kcd�~F��Cӓ����P�j�$���b\�!%�D^�P�ޕP�"o��9�ڋ��}��Κ~z�Z\��d���#�?U�0�-��P��z�I1��������`bWѳ�F��hm�3���®�s�xO��`�u>7�Q�����Nb�:%��ۻb0J�~��[��ء@9�h�c�'tE������|�������L�����깎n���Ug��pT�]�y�4:e�P{��*֊p�wrl�d\	��?��\co�4��a�������;�+}�X�!��x�9\;Օ�&o��qC������BSbPF�8U��_z�zK�z�%p6<{9��m�iԅ��a �@xPi�����_<z����3?�2ك˽�����A��B��oז�ؾ,'��ga������Vm�w�Bt��2<͕��9j5����: P<��/��(W���,�,~w&'T�H�������?W��_wYp���y���h�/�9�p#�7���+�>�*�~��Єܓ�|����&����A&�\���htyN��uG�����$�&���k���9�R�,�޻�2/Gz��/�\t��_N2�e8����1e7?Ы}�+���(Uq���z��K�kV U���Co�'sn�1�$ˏY_�d��1|E��n��+'�\:�ҙ�@с��>���΀ポ[��L��ߝ/f5����b��&	_:7��v�j��LD$<ⳉ�@��cN6 ��Rɻ%QT��2�A2B�j� c&�`+f�����13��2��tV*�N�s�:g&���������V��� R��it�l�o'��^�a[wO�$��$�`[ۧR��pD$lÆ���r�Q����p��.¿n�רt���~)v&��㺄U8��/'w9��9B���Ce����le x֐�h�7LǍ��<�������I�Hg��uңX��G���*��w$Ī8hABJ�����'u����RpYh���E~K$9���N�_Y
}����/4n1~��G�6�PӓsJ�ظˀ�T��L������6�%�*W����*�7��En7�[��T�kpG;�m�S�R\Ìd�?�t�;2�H�J��J�	.I㈋�8VR�0���Qz2?��������0k�v�� ���%r��=�ˡ+'�����ğ=,�����F���yq�UV�n���nWy3�H�O���[6�<�H��J���V��T��h��_��z�-�SX;�]5S��s�m��U�m�� �����>������;�=F�G��/^����VEb�(G2�E������ͮ��C�Wm�*ԋ���-��z ;Ӛ�u=
�bf��W����~���k��=Z7g�_ä6pH���K�"n>�n,3'4��4��r�����ŗzb���H���~�W.�!��]gV[0&�(��r�P�&�tQQ4�8���_�ؼ3;A���aL!.rc�]������r]d��/�Yu?�M1�[�Եt�vӊ�m��r�M�p�j��ѱ�3�ᆎ�%D�773����.SaN��)�� 术6kD{�������I��=5�a@�@Z�V�VֿU��6e6��&9��u,'$$�X��z.�Ҿ��� �~�T����=<��I֭�CKP�Y	���JGݮD���	ƨ,�#��w/����O�[�Ǭe�rug<&f��k��x�o^ ²+'i�{����-f��?����[;�Y����A��O@��I��X"w��u�tM����x)�%��y5���l��+������0V)}�O�;	�_9u[Q}�*�g�1jg���#�0���������)%f���;�u(c_�UE�Q���2�g�B_���0Xw��#s5��t���9��N�6�D;[��
ħ�d�5���6`+�LX!7�F�����~#�#�P=�wf*��=4��\u��pN�I9[�F�ZKn�n�2#�܇�����(7�$�9�H������#�ִ�v��;F�x*tJ�|�W^-[��[�J�0��uz�'R����*& ��ά���o�m��un��G1Ǯ��ù7��7�~�ʄ��N��G��Rn�g�m!u�2�E��3��	�Qi�[��%3�*�Eva���h/ý���w�n��mdd��AL
�r~ٳ�gٸU#=\a�������WS2�CH�62A��ARr�������&.Ë��e�@�f���Ƕx�l��NK<�\��.�KJN^V'��N0��Z}�G�*ݫ�J��Qs|Eh%@�fm�Z�1��K8�J���\�B��`�Q�X��+R�ը��R::6�d�C�/�ZOZ��_۰W@t����0�)8�ҎXq�����K�{�n�	��r����dT0b�_�!��|�)��b��tk�%H`w'R��!��w���0���P 0$V�Ζ�w�|��M����}~iH�|��ܷ���$��"�M��C��~�������[WN ݸ7�m8��@����!cN{i/�R��-�?�ٛ�w������R���ipJV�:^Lꪏy��Չ���*?���2#�Z�+���v�8�-V�W3Х���u��,�?���8Φ���'��}�X�2C�Y��9d�9P�a��0� N�N/C!|}�C~�4x�9�ܩ39�"�'�>;G�>��cy�}T}o���9t i'�K�f�k�Oga؂c�M��y*=��`�='0鬌X�n�����x�	�K�3z�}0�t`5w΀��n�I�@�l�N�]��a_&���E:=h��w�k��~76�ur�jZ�W$6B�)U�O�/�~7@HUU�1,J���؀϶�T<��i5+�#�>����-�)0��j����J���f �ߺq{�T�9����J�G�K�"Ȩf��Jvυ �H�����_	�[��\o�����ϰ�?�r>��:ӟ�Κ��Z��EP��Op�5���ܞsQr�H������EK:Y����G$��OF�y#E��o�V��#�\t���;��&o
"�o� Ȣ,�:����D�2���D�|�\-�0�T��n|��;b�*�\� ��g2��ط��+"�a��T�q-������	�Z�[5 [�$��&�ƤY���e���X�۴Ly�7��� �+���~f�O	�����ѯ�SB��;<W;���e>3mܴƊ T1|����p�,���Ӫa�U%8A�=~T{�@��O7�]�	k(��#������D[�&����	�_�|���j�q	�39�A�}_����
�ܪw��lcV:β�;�O
��o��Y�G�X�eՇS�"��*u7!�`�5 �12KKH�#�2f�!~bYA�Δܫ��r�x'}Iǀ�<šN�	K=1��M���)����\���WZ��hv�V�l�,���>��@P���?��x�̫dɽC8�gj�����mm;�H�8��2Э���|Y5��쳠K��ĽR�T*����e��}�9d�����%ű3
$��kü�G�|D�#7ӼBK�+�B�����k��E��藄8�rEY1k�Uv���lvW�cΪ?�qY�^�aat;m��1�`�B���B&`����lя.�k��θJ��w�p�4�O:��C�M���:���(L.j�HpS�œ@���!��u��e����jzW(C}w����(&���/�J�v���G/��K��	Σ���V�-��-��`9����	�U[Q��Xq☐Ѵݔ��B����)+L��x)�j��6��������ʓM������@�+�v����e�B�F�&Vc^&���j���T|C�HAH��m�������k�s|�4<@�'7��M�E�%z8P-x����l]z�g�w�`��W=��l�N�Q.uv+z#�(���ݰ�7J�|e5Z�����O���Y��m��(E|e���4�����Mr@D��t��0�,�)�L������3Lɽ���j�fTtK��I&UZ=�����d����(���pLX|�H����!w�*��nx��3��[/,�T���x��\4nu OX�K�ls���!e�>	K�?I	�R���E�Q�iS��vD����J:�Iy6nwQ�u�Bh�ʜ �,��PV�z�c��p9�V���j$ab�υQl������89����(��;����,�����B$$�� ��(�����h�,mj����o4�raE@����<)K���%^��9��k��q	���b2�P�5 �]�ι��N-��I���ku�3�/�7�\��n��� L��Z+�a
6/[<�j�7?��xR��'���ψz�$SI���Y�1��??}�F��;<":=%.Aƪ��pK%�00׮O���Y�ZZ%���0����)Á��s�,�1pL�v���|�"�*+���\0G�A0_���e�]	��2���$�������lC��8�m��UZY�wVjc!��z��ATl�;���#k�љ#^w��/t'�D�$��v�Pf�'��tqђ<R���C=�78^�*Dq��5n&:]`���0����S>�c:�����}���hmN(h��H����bfS/�&�r�&�9���µ�GG+��ID�+lH!�*��f{fw��7�f�b�ǷK���K�`��=���d��������SQ���u�W����T���텍���
� \T��c��u�驠�u�۔��k��;�b�w6e�߂$?�s�$��y�3n���3������%��i����f����:�ux��j�C�XS�XWk)Y�Yn7�ZtU?�fNr:wM�M`�Ԕp#�`�Ɵ?��$�� �L��z��P�o���ah9&f��vKN<�~@'���)z:e��}����7�)���s��4��@3����<�Ğ"�nD����A*���)&���x"_����ʞ�5~$��a:d�c1C�+W���0k�e�`ދ�@&�G�;�}�@�S0���
#x.�s%^Ȕ�AŞM�OĴNv���yL�3\��I�Լ�a�Zl�Mй�R�@������Ow��n��6{*՚�����đr��K���x�a�?���p����6i���E%�b܏��;O�s^�o8h FI�a�r�����3#�!�d]���� ��r-t����So�FE��#!BS0M�b<�l��{J}��Ξ�'�N�;�����}���_�r�t9��Ԋ$��%G�M�t���-����c�,��_]W��qFUI���U��4ـn�Zў���b����t{9Lot�y�_�K�ӌZK�Tw���,H�=��[�Nu�Gv��t��!�:��� 3~� 0��ͳ����p����\���-��z�x�z�G7�[My]
I
<ǀ��8V/���+�l�+4��O�����9K�ި�4����^��W�	K�2�J��ګN�I@�Cj8�%0�`>���G�2��	m��M�Gc%Hb�E�2y����B#M�mU�hϧQn�ҏV��K0G�ՃK�����\��P2�?��͇e\��8_�ⵇ�1z\t_���Њ���K^��-3,���=MZQ+��?lN���7��3���z/���Yg:Q`��P�����.�&%�AjI�C����<�R0W�����6Y�������G7Q�?'����S3їS��HPǲ<�@���x��e��4�#�ڡ$�p�S(Wm%�{�}I�@5�TXV�sT��|�����bEq��6�'f��y�����ZإA6�$1��N�"X�G��y���8��԰&�Q	�ꁍ"ct�:I�D=f��H�e��\�����yO�-�f�M�W�j/|c����g��q|*���tٗ����5X����K�����# �M?�ltHB�5�Ku�O3Tt4˖��R�+�ı�kt�D|<~fKW�c���e:��eh�4���t���&��=Ӕ!���ۊTU���RK�2K�-��d9BK몲���u�*MX[46�����t�Ȁ�L�G�ٵ;�n�-��
��D9J�p �A7
���l-al�˵�I�m��r �7Fu]�Cmѐ:�s��g7e���y�mX�\"��Y��B�Yi"�fބl�Eb�Ĩa^5[��%��?Vqoy���{�o�-4�o�Q���Յ��wϝ��z��z��3z�Ƀژ]�暁R@Z��bl���1�DC�B��� ���,�\�����w/����vU �.P3������%W
�w�H�*��Z r��� i&t��w�$�A#�t�;/��O���.A�=B/y�!�	��'�t�,����@����;��2'->�ˊ��c���6-�C#�I{��:�������wK����#�|���[�ң\iF�
f#�y(*vI?F#P���]܀*p`��A�8l�?����G0�����;EĖ���`{�"���1łn6b�J�N��hU����9�0^7�Ě��|(mŪ��[nj�'�>�s&���l:JtG�6��&^xe�IERY
Kn,-eF,d�a��	e��8�2c��ܬ.q&���`1�C����u�88�v�/;��ه+J�
T�l�э���������K��?BT:� !�;`4�d���sW*ک��;5�8�`I.]N9	�$I�뉲�:"�~5�B�z�q�A�Q|ƶvv)��5WJ k�G�n�QApg*�Pc��N2��<xLy&҂L*<��>���u�K-��M#N�&�%Iy��z�P�1k�I�S�ۥ�z益��E&2q��4h�΢�$�_���=��[A&J{��u�\E�HKN��O���Ζ�r���N���!t�5e��q��!kpF���t����2x��n+=ؘ�E�S�9��B1���p�}���#�E�{:��`�Ʉ���u��A�,KI����C��}:�.��.[�?�s?y|��&=�����Kv�������[�N,W��g���#�M�ʫ�F�;:���nK;�_������Y���+�c�����9e(�%�9��S-δ���'�&�l:��pL�V(��,i�Et�����[����	�KaO�m�,�wax0�	`�x�����M$����@�D��!n��K�܈\$�*���`+&�]DjE���Q"B<P1܍\�8d�l�1������aQB��k��h=��$����Q╰��g=ܥ�K{�m,⧖ 2��ޘ�N��ׄ�����z�?۹�B�Zֹ�8��1�yk%�4n��R1Hn����X�0܅W�������#w&ƣ_�A�2~���O�)��4ݬ߲���];Ul�F�|�Pq]�@��ŭ��b�w������-(�G]��vU]y1A��[*��y(���xxY˔���V��A�A�|���N�P�ΰ9F[2��d"���}��1�U�%�)�SQ�΅���X:� Y���1zݫ1�J��̧a�hʕ�-V�A� �3����%/����k6��H�x᧿�nu���0B� i	�3��J� �+	Ֆr���c^�)<2n�*DcDJ�����s��Џ����k�1>��E��B���i�;
����hp��B�`&3xA�urvK2�JEJ�`7��]i4%Z�#����OԀ����N����'�?��&���l�\.�������f$1*���=d�[���j�YI�}	��-;Ԙc;�LB�E0L~�(���p`V�e�B2j�0�7��s��4���|T)�d�l
EȮ�1Ym���Y�a2�l��T.��N�@}�!����?x��,��f��0����� BZk��C�������=�ѝL�r�,ר��R
�����Y�7FA����F�/�vM��@Q7}�=y�S�ym�V��]"�G�U��G��K�+l�vl��rKC��x�S�)�8Tjp��,�3-��������'��NId�_gʉ������,���،𝶾Xt螾�hQ1[��l�޴�����{��H�L�rXt9Y��F�Io1�����Uà�o�Eu˫��inm[״�?�t�Be��+rB�<n�.ͩwM��Pe�7�J�'x2���l�%] �oG�ٸ�&ZFw�o��=NF��`��?���E��(��s�B�T<?7�7L"�����Z��9*G���r(5Gp#gE~���>2��n�G���ї�������69:�z�a*ǪQ��'�����e7�!/��c5��up�I���h�piB���G��S0i�Gyf�K��j�#'��P~������̼�
ɉU���w[�{s�!�Y���X��HF1���������
�Js](7�G���#�OiU��0n8k^�`'W �2ZV$��:���q�?�.�L�d�=��G��N�A���L���:�	Y�uޞ%��9�X�h�;�������P���j��28o���U$�}���m�] ��qS����[H��ӳ0���-R�B0/��0�=����|Ⱦ���L�%��;@8�
}��{t��["k�=5]"'��+�Q�4�V����I�W�:��/�X�l���:��%!V�b��= |=�T}��{*P�(����W5�� }��o�-M�2���ו�\��$�R:-ϑ1�.�'�5T� �/���XY�7��d���:� u��V���!�	4E��<GG��@�4��}
�{ì�p��7���@�rvo}��wi��	��I�:M�	��,YH.#[�{�HTr��}!�9�1��H��%ɳy����TpEo�����d�ꙵ�w�㻪?<��_V�������il�@���q��+Z�L'���nb�3j�� �*H4Fu�չ׀�����u�.����D=_\(ŭ���K�p��x��{��`3=�Ze�����E�~����5R�!=y(�e<�F!ʁ�c����Ll����m��	�T;ߛ�Ob0C&�F�Z�`�to=�j����K��{*�:�D���nM����jF-��,9ZR����6�����K��ٞ}������,b�"'/2�f�jM�eS�"�7���L�/N��Gw�'�š2���~�;&}�K"�Q�[p^oZ��ݚ�Ԓ�.�ud��oB�&?�y	>?d'm�]�ͫ^��ĥ>8^� �rSL��B��kU��OS�-�wEĲ�j�/^H�^��ڧ��S�;����Ix��#n~{��_J4��3��}��ĸdbŐ&��i���ݻ�4uZ�pJjO��\-�����|ǿ�����^�%Z����Q����VSZN�Խ�&�&��
�F RZ�q�k�]T6�V�4Jzߛ��������(�֭�A�q1l�����m��O�l��j�حe*V�|��+Ս|��Q���Y���e��=^�+/��u�
�3$�[`P�O����{�p0�K��tú|@l�50E�f2���b���6�g�i!پ?(��(���s	6�A5.(�Z�V��6����;�:vI��ʵ6hd(��S�3�/���YU=`���͉w�_�^��,����]FkRn��0.��]2o���f$ӒYA�+��9�o�O���C4WH�1�q ֎ʣxƁa���7��0�7�t��S�pMkO�����=���g^���.���R}@�82���t�&q>��v���f���S;�`�,�R�ύ�,+S������z
����}A]�c�u6�)���8-/�7lR� ��	�V��V�ad� �~b!frX��hBf7*{G�E0��R��BDTŴ�?Z��_��_h�����D��8|��X���؉z�+�56-�����Ƿ�&E���#�L�͉��2����G"Hp���n�l�e>q�j�iA�Ie�'����F�/YC/�p����>$��2�ou7vb��D�DѬo<Ioo�测H��0���+
7VM.������V�D��)4,�������t5n0+nN~x���6⁀<��1�r�E5-h��j�ɡ�`��T�lȩC_6K�Jݨ��"
R��KH�Fțe�^d�!�爼�צ��
�zIeW2�*|����@� o0���Ml�u���T�aĿ�/-�����Z�W���@&8����B|�&�'��:B}�V���B�y =��!�� �q�ǧ�J�9�
�$ڜ[!�E���Fj1��̀��\5!جXX�h*��pmJ�M�ee2�f�<��r��U��B�Ҁ���!�����m�EGz�"nB��(�5sHu<�--^�	.3�2V
VTK�����éd����mA�ש$U�M� ��\�Ӆ��X�G����������&�twy����[	�[>��P�W; ��9���x<�����xJA����k����1#ph�T$���m�����Ȼ���Z3��.�l�PD�.:��=/������X�q�;]2^�e��T�|D#_���)�1NsU��`�ޭ���$���|OZ"uUCp�	��&u5DM렪<���z��9I��A,@�[�v�m�Yk&�	���w�D��]����� Ʃe��Fr���l`����
~hiH\�4��N'<��*�,�v��%ډV.� ��|�F#���_��3��'�pes�(7�[�M��R�&�A�g{]w�|J�M��x�
��@K&E� ���1t-墭�ztP��e:�����֙;��h�A�]�4���iн�GT�'�"]���ƌ���Z�0ߞ�*�����3's��L��޺�8��{i��-�<��&��ռ*@�� ���z��"���P:��q�8�������̄���l�'��a����ݨ�G�6&_�J2��NSW�A�4!�Ե7�8?����p�T`aT+-p���S84Dz�ͮ_����疪���I���&�i!W��	�_6U�*�Iנ��	����f-���v���ؙ3���:BaV��B��������:>�����@�}8=��I�)]�B���RH�j�fh��;Z�	WB�I�m:�-��Q�VE?��H�^g�qVz����/j[{c�2�
ٸH֘�Gy4��.�]���OD!��*�zF�`�@�
U��D��r��;ѲH�q������%&�n�ZiXc��� 5��7�`�]��T�rq��!�@�����G	b���F�}�^�A�Ɯg`�>v �*[=8�VGa߯�4�B"
�vFH�
�}\B�����8��fYU�z����d�#��N�����*̅e)�͌��B�����Us�mp�u)�c��^Ԓ�2����������A+GgO��|��$�~�SC����u2������,���ws�n��J���e#(�@N?>�۫X��m�`֭�!X�9��/���F��E�T_s�>�`��D
�<gH6*b���xN�����S��@mq8$E�2�[��6�"��{ �j��O�6S��"�!q1�w��W�G�ʸ�8|��������Kr�RS#�7gX�+�\a���?��v�`��k�>c����䗫�����n��ڿ;��i�Y'[bt;��v��5 H�.b*��U^������q�(����D�HA�k��*h;�d�a�De�2�V�;S``�>�����J���<�"oa7��&گ�y��~� �g[�cG��T���
m!f]�:3�.z����g�B}�?o��2�gX���E7%��?�*_6���iV��7"�q��W��2xK��'�3@��dZ����{���׎�QzN�����՝dg�<V0Ѵ�;9^����g;ฐu�X=
-XXN���Q�I������+��:�*E��v��<��)�ܬ��"���T��L�7�{ۛ��0��'$A�"p�}����3�QRT�A-��5����� \MT#DH�wB�	d������T�gA��o&i�;����.�(<��1`ε������h�6��T���;�i���·�����N�|n�_�1�>�/�\Ӫ����B|P�ϯ��J������>yGA릥��W�eH!pZ�f���ڇ�sub\�4���%Q ��e�;bȺP!���-�&�:�;/��p�iΝ��Ҷ�saN�䴴��`�p2��io�}/���e�iR/��������:@6m�c_\��i�t�\�M�M_�K�u�!2�L:��{l�ŌK�l��)�(	Ƈ�V���[�_y�h	mt4��ӵ��
��bu��2A��rO�i�7�kum���Y����OSH�$���8U�6���O�/�q?>Vŝ��O[�[D��'()O�/�)����mk�����*�����!����~������m}��=��<	��ıy8�+��_�&��#!�XpJhm����Ȱhut`qd��?4��"z�����A�.���X9y�;�Y�G|	ʫ?�~]1�/�&Ϊ��\(w�廂�G`�z����Q'��"��Zv��XU �	P�B�ߺ??��n��^*::�
z�"[�ə3����/���u�P�<ӊȞi(:��\� ߱���:^�Blo��"�������̐LZ��]ƒ�P~^P��p@(�[��?�:6�4�$5��ڽ8q���h���:��2��p�Eb�%������P���r4��%iu�B�!���Mf$��2�O�K�q��ű&�����b������eqNW5����h�d���1c+��&Pq歚U,��姒�㮾V���`�s"Km��d�^��$�F�0&���ϫ$���c��_$!xS���S���6��R<�$�'7E��V-�q���*{;B�ȿY��c��jj��=��o�!1|5$R���M�s���F<�}!i�c��d�y& .`{��5]�t�HGd�~B
����)��GG��4%�u�ى����N+6U��.�ѸջX��V����p���0Lk�+�2~�(�07c:��r���%r=��6u;Q7��)`��rR���~:��lVs�|��L +_G˙�]��b{/٧��,�VuP��%��ϓE�XMi�}�<R���DY�B����[p/(�NsR���L�b��.�<$���vQA}���8D���|���;D�<����$��[��7�X�9�uf]�!��5U#8���e��j-^y��=W�~ǜ�n9՘t����~�E�t��#�m�P�$�R�%05�}��1zm;w����~~�tNP*������D�;��w�q��̣T��6������k'w�'�j�����k޳Fz,m��\���.�S�4-פ.�t��T� �8�N6��mȉ0\�kC.�@/�w������J-�x~�:�zoa�F�-L�L�.�i����1�
�S��+h������v��B^����t���V��e{�Yy��pd^���$��3��]�06;,zhu��dz��}�B��z���`Zc�31)��U nVȵ��(��)FGfn����)�~�r�@��:�p��굻�)��V�\��4�Ñ1S6�~?�փ�Z����f�ZQMbJv�f�Ʉ�����v{43��0�倃�4��7�9��R�X��|���eimD }>|I_H��SH�H��)���`��Wu��
�7lURMaFe�1.�X��w�F��6��E8�ĳ�����{g<���>�������}NO�|o����.�͉�<���i�O�wr�D��� �,����A�Yo�ר������)镒5f�� �L>��i꺽?P�1���,	d�x�S�ܲ����G�IdV���%}��@�^tK�x�Md_}��aA̖/+ES!b���2���I5����[���R���vI�"@�&RU�9i�� �f���	��xi���~Uf˙��eB�f��Ӡ3$"Z�jh ���g���Oy�����Ld#Q���,�-Q-�"��P���P��B�RBm+z�#)���>~��W�ƺ��?�n_�}��t���$UX0;! ���=�Aa�"t����kȅ�j�W1&�n�%�;l6�\kQ�v�܈�����P���/6�={���(���5>���:�A�
8�Z�ɾV��Z�1`@g �8�RS(N��O�����W���V�히�9�yA[8�q��ʬ��U��&�*]
#yY�����\��&=�*� Y"L�o���(�hsoC�9�0��A�4A��ue�j5��_!ߟ��P1p)8� �E���$���}~!u���E�.b�q��� hZ�`+B�{�y%x�)U�������S�S�p�9e�5ZFz]�z���l��q�9qW/�~m�R�r��:xS�$��u?�?"}��PmX6��m%�ˈ��ck��F��Zf�<_�X �Z��_�n*F���3_�G���E���*\����1�H8�[ѿ�"EY�|M$����������l��� ��P�Ь�۳�X�H7�3�uc'�T�R�+3?6�)9dŞ���Bݕ��&�n���c�E���� R2����Q.����_�����n.�bY��R)ՓK�'��Xj-�rWpPßkQ��z7C�t��431�95# �#)b�-%�
zr��|1��f��,uǨű.��&P��˔5��ML�{�pO*���Fz������
î�e}��({ӿ-�H�PB�I��/�����F(@��Z=�yq9�ޛy�so�!+�ȍ2�P�>g��w����ld2l|�R�u�����������`$��{���*P�i�Pc~����/uS�SW��
�uQ!�YA�K���a�in'��_Q]į���+^��`r��?T�x!�曏-�w�e�w�!�](�5Q1�M��?�	��+�KG�r����T!=ѯ�zʯ�����pz�>�Ra�1ݿ�l��y�cn��%�B�j��h,1]�Ek]p9BH=9��{X�v�Q������	� C�'ާ��Or����� �(JQD�:�a���qڹ�Z]P=r/�����3 p��%���T�2z� ��u��0��arT�Jr�Gx��3N�����/Du���W�����%�����(�˳��a�8�0'�w��5&�:�C�@}��΂E.�3/�D�!�U�w�{If�q�oggj���b��BI�Z���D����z|�*�5�7������R�7>���{�G��ve�{�^az?�j�2<6Ǿ�Z8�1%Է�ҳ,! cXE�<����	��$s��\�h��%��̱$
d���$�0�6�=*D��q�G���AL�1Drh;2��ὶ�U����@Q����0����2��fҤ.>c��(��aJ��O,S�ゕ*Z&���V���G1�d�	Ֆ����~w]�Db���c2��>����OtN)�~4�(��B=�ŵK���O�z�{���f�m ƈ��H�= ʃ����j��n�zL%27�~_�Ӆ��N
I��͍�?)���M�f �P��h�1˅��80?���<:�V2N�(p��_K�Ȕ���$�&ڳ+�{g$R:*�h.�G��'t���ƕ]��-�6Eo�&��68s�,>q�knϡ��u���&l�sf6���:��D(3��-1�,~"����+�~a0��#	��$��oO�Z:�kC�<�~��*�(G&Ys�8 �5R)sM5��Y��YU��2Ƕ#��#�`���x��|��:��Y3c�.�C�8�4V�FC�ߕ�3؊��xZ�����- v'�>�@K��+���'�<Р�������o����/ǞH�@n�s7&B��bq�Z��۰QB�����	3P�<"��b*24�Q`v=3Ug�K�djJH��q��`ш��� ��7���ևa��MT)Gk��� ��~ekU�@8������3�p.��NE����T��=�'�+�U����dFX�Cd�Q�������Қ��-���?EW1y"��Ӥ����f�fB����9����HR0Q��j��[x�ɧww#Z�bȸO(��-����L�At���֣+O�\���Y1�1��k{�6Fz�t�f,.��W
�g��e@�d�h �d�IZ\�������Ō`�����r&m��]���+^7,��4��h��TY��-e��Ƅ��$�<!�i�>�_I��ʅ5Ft�X7�d��&l�0�(Fʼ��52��G$�QȐ�Z��jF�@(�Ƶ��)�$\��L%�h/= ��BD������YiӁ>����3W!wBb����<=�J�В��S��qQF�S�N�mO%�oA��D0)J�������L�?%�О�40����}�+cuy9����k�1P�A~�}�;�pʦ��Y/��{�5e	hcw����ʼ��ˤUm��!p�u�*q �*��U�+э��#�U	��<�r���+%���fe�W�ת���Իe���.3$��m�4_�����O���}� ����[Y#�D�r!�"Z�����-rV��������ֈ��`���-m��w-nm�S�Ø,�?AG�����.#OU:7����HV�.O@��p3�!2\��w�!wN�Q��{��8�&�1mko�#�y��f�"+�O���'�ǡ��,���jy|�g�ԉ@Ba�l�<��ȫ�s]C,��H+��s]��L[� �-*-i���-�h&�	81��0u�?����vq��/�_��b���L�B��!/m���2^��n�Q��;�?٠k��EO[�~-^�6�>~j\��<V��PɡT�5`�����o䂪����֘(��������u7�
mD%�e,�M�S�����p�/<�oT��*�(v���Ϣ����k��f� O��$��T��+��}������$r��1�,!�t�Q���;�F�\o�ʙ0>D�}T�lZ�E�Ѭ"��*���N�1*�(B(�x�Mp���ћ�\��ГD���~��˖`�6�&	=�K[�ԭ�W�R��k��=�U���-�Kխ,C�؏�t�W��~���m��[��`�۲T�S��g��ؾ�b��#�N��§�7e�x:%捛��x�_�a��"C�w��S+�R[bJ���
В�xF7�G��g�/i'8:��Ѓ=E!D.KT�G&��cj5F�{�PU	�b6��!k�x��(�8�l�C�%+1�λɮ�%=�D��c�������
�C��bMd���#�ZqM�S6�㠲X�1�i��ЭU}n�w@*(��g�I��H��'�2\Y�;�@����g�����OA�Q��!��.��ᅵE�/�w�#��X?w �n�~�RhhQ�˙���K8W��b���lZ�g����P�y�+���+S��Z�s�e�� �
j6��r^]l�8�f���ELy��M��dJ��Y��k�[,��h���f�Y>�����S|`� �u\~5uQ1Y �Rßf�6����I��
[S�X�5��ӄ#�o1Ӓ�.��F�x��@\��k��\N7��g���L=���D��(�6h���,���R��ҭ���1YG3mQl�Yr�ru�û��	a�����w�;�m �lA�����]�LL�����q�����-�3��Vdp���&2}'��r�	I���t��g�ې&����q\��ń=LT��u��P�����Yˆ<���ʑ�X���Y#�$��-2o�Bդ˺��{PZ�pHO.b��.c����=*/ݕn2���=�d����*3�@�M�x30Ց�P�a��2Ӻ����Xq+�e~l'*L�\\r�*�l��6궩�^�1��Y: ���#ꢸ��F��Bw���Q�#U��]�b`YK����)��$m���ݯ%����Bi��D��Y�2��]t	f|7�7OV�wG�|p1e�U�̎����K�g�,hp�"���Ƚ!���?��h�t`IA1{�����Y��"j{}�K�F5�Q�v�l}��L�ֆ�b�A�/�|$����r�T㐍	�+�ؿ�9tD����t<��
v#�Vѳ�)��Ȟ�e����T�����E�KIa���2��kS٥���;3w��%�Fөw�wGCR�s|kF)X��X�}���k.���[~N�W̟;���G���p}w&��7�a����s�� ����_э*E�ƫ
��!�����;��#��	Z�+�i-��-^�W���L�f@a�v��Rs&�q��+�Yg8����m&�H�u�<_��S��oPǵ�H��W�H|���,��D�1B�[����yh���01Ռ��D�����<�9����$�2�` j��/�(M�O@��\ζ׉�x��d8}h�ߤ�Y��l��1đc�N0�4*��e�s<6~�t�I?l�1��s;���2�e�â�@#֤�s���8�_us<�7 �PH�����t�u|��n�W69�T��
ۥ����iG�w�=�LT�Dr^���,Nا�7q0�~�ɽ�y�$�?I