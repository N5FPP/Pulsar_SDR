��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��e�ik3�������w$����g|��J^]�,^R2�D����د,��D� �4B��|۠O9\�N}��?�N� ޠ������<��	o�K����p� ����H��''���"O@]�U����������aMϦ櫋��H� �z���Q��勱��:Ĺ�n8X?Qj�� *@��\�D�/�'Z��^��rw¿2X��o�ph�Gv�y[�A�Q����FlFL�)Y^�Hӈ{0ܗu�^)9,o�竐.���&\@��*\�0�qޣo`�}��|������$ݭS�"��}Uf�]�
�I8D���X��Z�Ⱥ����;����������+i�����Z�CjE�JG�_޳�m�L�C>�f[	XʶF���i�Ryq����O�'M'y��k�Q9�Oѵ��-O})�����!�٠S/��<WU�c���q:%U�]R�&�#AϢ����< �t�B�a;�P�>e};-�([���� ��ܨ#��������Z�۟����0V� آZ7�Ju�#)~c�_K>|�Cߨ����`2|�U�x�p�d�@,�,��O�
�W���¬9���|� �iq�oSP+����������*79`��h��DH�E��U�G	hٸ� �I�n������_�TU�#�m�7NGѤp�S�&�s����cW���Dctd�{���.c��Zr��f�Ͻ���Y"�_����RJ�#bJH���c|���οW̍�ѧ�������ڊb2S6�d�B���=��2���PN�L����͟<�:,�J���0�M���5͋%=�Nn>}iο?�5��r��3/�N2ϒT�Is��C���>�@.�{m��
��ѲZP⡒��¡����`}1Q�4��t�����(�`���C�z{å��H-�lǩ[��C=��IzE.����9��O��z�R�X�H4ÔY`���A7�0��J�]�<r��k�1�L�Kp���R�~Or_��VW��}m����ϔ2N"�͐fq� ^2��?;��S'%����h����ўL�*Lh���r��i�f�@��(��}KN�G��3�{�A+��ᒫ�Nɞ�F�!9�C�B�	2H���%�|���`���)O�+�j���qe6lڅ�	�a��I��m��?�qM/TU߅�N�0nz���	�Sv��>��'5C�
�
��h!��O�ף�I�"C����=l���-�ߜ� �$(#�-y��X���>�V�])�(����|]$g@e�%��<Q|��5��I�Q��BD�y�Q�e�����3ۚ��h#�z4�{�9�#;���s��0R�>��Q����G��u���^���wY1�|�Y% �drFy?~�2�QWQ5i��.-�8��I)rK�3 pe���&;qGFߒ�H�7!	:�3�y��y!(<��
���Z��P�����،c��J�������8��,�ʉȰ��#�q�/��t�B�)q�C��6m=/:Y���f��G�>����,�f��F�:�5�Qd��3i�n2o��{��|��|�{�N�rf?�����Y���0���,���'X��/F@�BP�H�8���gJxM�i�9CMMڮ ��t� Z���ڀ�O-Q���u+���p�dדk��$�z��A��jA,�,��Jh��j�3�.����A�g[��-�f��@�N\�E�� Ѓ���S�7�p1�\6�5�AU�:��x-���˧[HT�c��T�Q�fj�d�Y��N�.��4J�/���Dk_�G_d&q(@��yUim� R�=%nX���Ő��������\�nX?�Z3�s�b�aK�H�7Q{@۴�V
K�o]VԈ�b�Q��Cs����C2ؐ�в�k2�  NOA��ǡ���R������r�Oz�?�aX��4�EȲ�X><�l+���)?MH��f	�����Ǹ=��H^"�l˅@�4����&��m_��^A�g����a�4U�� ���-$��c���X��F�L�,��#g2��>���ճR�n;��C�6��y���	`S���jc�e1�Z��oӿ�`/ǲ;=�܆��7�/<���&�7)���c��������s������y+yjrYyB�������]$��]R�8}]���$4&�Y��hsO��#~�FxDU����g�.�g�xò	5�N�����)=&R�I����-�;)��;�%�4D�U+������/��"��$� �L�M	e����!E~���P:n�t�,�Oc�?$�?;�FK��{v����"�$�0��.,����g��E�1vIݻNl4���x#��	�C�­A�}�2�ο4*O�.�͗0O�{7��b
^��%#�p�F��Ɯ�c^�4b����Ȩ|�6f38/v�j��2B+���aN��HV�G�79҆��]H�9�`&��S��{�7W�Xq/)m���!`$�<d���rh�Įi^cl�d��e��ӁE45v�:�^G:��w�pD��t�v���|��G�ml���ń�P���DQ2�������RPy�.�Ac�.ք���xQ��y'���"��� �؅��-���l]A�H�K(��u�6���k"h�έ�Ч��G���Vju<�Lko�d�i�Zf����w6Ǝ"l(�v��u�4�<���_"�՚��Q�i�/H����ɡ�("��j�%���.j�C������@��)�V���7(?����:��l^{��y���O�\15�%�'�N��H�rg����WL���������u%�oɉ��:3bn��Øb�U�n���3G���B �XB踣�/�������(,�<@��.A��qp�_�Rl����x_�]����rE\�XW!�s��;P�c-4cܟt,�;X(��r��-�޳�O-xN-����B#�f� $i����k�6+�����z�Je@L,Ô�jD���|�^��j��r;�@+2ޯ��"��В��5ޏ��g�����^�#t��i��#N`յV�k����{���a
��Cs�1⬀m�����%����nd�m|�:�J�/v��L&86�䔲£��o-�^�h�S�5Rl_�}��������;˱G���حK-�]$�6A�7�m�i�d;�8�2������fm'��N�A_({�szi�gj3�4Қ��o�!���J=43	��}�)ޢ����/s��q�d� �}�yK@�L���g�lI��jz1��5{�`��Ą��C���j�A4 �?��U��Չ��yc;5ϐ������؀���@�Mx�����1�j�W4�gՕ�3 "a l��� D)�Ѹ:��.>��o��{����;�M\���ޚ\�}�F���x�ޛ���.��*�9/��Vβ.����%�h���Nu��z?_z|(,�@ =a�2��A�f��n��`����#��g�U
��5v�@c�~l��Y��;�㋄Qץ��Y���u�5�4��n���*L����مع�.���5i�y���MS	�A�'P�����7R!�z�J�%I���+��Vw�|nz'�,�w�\+Z�jP%�*F���8��m��t�&�1��o��D��������ll�Zͷ�G��r.4"m"���c�w��C2���� �m*N��ԁ�k�$�AK�f�z���jM��g�ĵ��E�n���d�?j�BY	m��|b=Lb[���X��oWKL��a�
�D,�EE' U����J��,��Y��2�V��,E���X��/���Y����`�N0ߓ\��� �0�X�{� eЌ��:h0%ͰÚ{aPYD�x��k��������K#(Q"���gq
˻�	�~(\���y/ކ.��#$q���(�# ����2�������o/%�-�Š%�Jԃ
�����g2�Z�4�c �����U��W>����Z!
�s�O������"觘���I2(��{% �VS~2ZC�3�/��f\fNrn�B��U�%���_]�aP�L��V)es B�?����i����S��٧~��s��H���=[�b��;-bS'�ҙ*��kn~�(^����P8/��
�<��C=� J^�_u�.(SW�����[��d�2)$�ƽ"�y�dc(�>;��Fd�9��w����nc�k�|}Ic��ª>�ax讣�fI�#��D��K(�tT�S�Wf�9��~o�+U��LX_VV�n�n�M�?Մc� �>�,K��:O'���l��[��:4��^	��$�@ž���' �Ns���{!��DX�ƛ�S1��
��j�H���j'3O�nb�a]1tZެ=�u�}�a�͸H����I�a�Ȟ����,�?��<�l��G�(�4�5[�4�G4Q�
A�O���v#m�-9�K7V��+�]r��Δ�۫��l^�-JM��I���\�7v�'\S��7i�6
]�Y�PZ�����Q��3���T�u�� 5����R�	�l�kZ"�W�����|��(��&Hv1�W
N�I�i'��,�cj~xd]��-I�Y��ʭ�y��BQ���u��m�M	������ڑ�f�b�\�2��h;����W�z'���zߪ'gF���P�g	�������2��ά��0�5M�}NV3�bh�w
�Y�0�|q�>��rC�m[@n9�g+�f�"5_iޕ�;V�dɟ;\*�"m_�/q�;Yg�9�9����P�z��S/@�Ti��# ��o+4�|;�G�d}�f�eP�qI���k��c�`ġ[(R�&J!�i�IN�iv���/��5�m��]a�L�	��З�٫F-֚�]5�	'��O����-�"E�#Cm��u� Nbh����v"?�|k��~����@ώ�X��d�4n��(���/Ѩ+�}ߒ�E h�ޠ݄"�����
�K��-{Hdh}�I^G�*I�e�ǳK��o��N�Ȫ�;��P$��J-�^߶=���[�Ƽ�)����lp9�M]�Q��u.��!�dǘ+�Gw������� HM�����M�~;n���N�&�j`(�y%^m\9��
|���5�������bo=*׺��3�5bG{%���Rv���Ȝ!�� ����ʏYx�`'���!���D��`\KV�$`�G��t��7�G�����*�T���=��)=�^z%�Z��W0����l~S�gE�1�!�T\'J96ϯl
G�+���s�~;@���� 8hn������
��V�dUYi�����]Mv��\~�>��!9���ůEpr/�hMl��iB�w�)E!���e0
�W���%n�ᝨ�2*T��C�k,&�M!�ʓ��pR���y�-,S|�` ��޺./x�K[pNw<��Y�u���p��<6�����{RH,�FO͟x17n�S��u�=]'<�"�����]�Q�>D�bZ�i�9B{�u�q�4X"���s���@���2t������j���f����Iě�V)"���J�I�㭜֢��6�"����D*�wF�q�( �f9������8���#��H=�teڷRj�����aϺ�˾�4^����#��hL�KU��5E &b�;f|��f�<��@!�7���Z�Ղb�Y?mE�Ĵ%Y� [{z2tr���1Xj᤼!Is�f� uz`l9�\�e�ŉ��I�����������Zc7�-�~D:a��m&Ԅ: ,X�A�}SDI'����&K����.� ���N��(�{�t���*s�^��t��R�z�Φ�F����Ȗ|���OV8����[������{xyD��5x�;y�S�->px�x,_����[�K�"NVM=��g�a��s�|�n=O-Q���5�`��C�)f_���q��������X�T$���>�f�w��ˑR�l*��"���~��~$XʑLn��Φ���!�U�t��Iţ��ڂ�&0�:�=�W*�`C���'����1S�<���.?�=�-#�"���wT�tԑ�"��v�F��(x����T���@-=�"�?�D�1*Y�*"�c?�x��Ln��>�Nl���C���J�,M8�p#s�%��E�(��ݟj�a���.X�+��<mQ*��7���jq-~�J�[���vu�^��J����*����B 4�YP�|U,�a��4@Zd1*9�|�йo�` n��`0���P��9�P�<����2�?шFz0nKp��]�e�O���>5�T(H!�kxzp�bcL���]���)�>��x�P�P�V��|3r�D�|���+��*�l�EK�*�)
���ij=�(��,�	t��v5�'���4����HA�';���yc,�aq5,���؎
��&J�A�=%Ҡ2�<D�\�%7:��u|Z�V�N�9,����	�z��mT�L��7�G��8���CT�(4%��ו��4ʲ�Љ0�y�3},�z-Q+3�b�*a#�'��;Z�i���sm7UJ��ͮIMi��5�U��9`e���S�P�i���|�o��iV�����5J� i������el{%�ɟq½�aWw@NEj�k+i�}���b�7�s�ĭuGX e0���D; �-�e�¬����+����3���i��؞��0w2��_�qN��XR&�zP/� SP�T�����odI%�%�Wf����7�	2�6#ikv�Zp����%m�3�v�혖���i?�	�+�d&=��W'�E�t!p?}�k��M�0��@��d�:�������m�;�ǵߗ����x�_����Avkɛi�7*��	���-#�'��ݒ����Ӓ�hΪ�驶؉�Gq��d�����J����o��&�b�#R��(�&k�2����4l��ٯn��j�.�{v�2;w�OL�=��S�eB
��r��G\��~�z�I�o_�)�-�������tn��S3��r�
�VF�Qt�R>�����R�cJ�тa*�,�	���4~�C�F�z# jz�dGn�g\����d_�l;s)^s�u-����t���v�f��-�X#�c��l3t���3�E��L�۝�Ϛ����6*��v�Ĵ���n�a
�U�U�F٭9��0��V���Aj�AD~0�^���2�PX�Ʊ#�0@w�8������x?�����r+��ƙ"����#�|�LX�Tw��1b�K��}yU舵9vz��P��v죰��͵&�{�I\��6�r|�"�b~l^�L[���RܴZ1Z�h�f)%�Pʯ�[o�at2����l�);���H��b\L���0�m*9�߆[�O�4�~b����o�#J%	
�(�6do���z�׽���*�؄��9qd@-p�mKf�`[v��/��u��:jF���#V��o%�>���
�l�H{�)$k��C�'?V�Wq��D@��eA�Ύ%����=_v��¹�&�\njh���8ۇ/�3MN6�[��g�tU�G�����[O::1#y��O.��Es6k�MN�X�33.4�W@P��]m�EM����oB�Կ�`��`�L��$7;�yZ��rԪ���S���I�?Dh���ߒn�~�n}1١P�9G 9��FU	CdR����M���p<��U��SL��EZY�p������=k-�2��hm�u����f �qlh)\��̼P��E]�����	/��ꅐ�'�D��|��-ѩ��8���R��x�+*s/W$V ����ɣ̆8�<ݼ���-M��V>Z8�B�:���?ۂ�ٹ�3����?�h�
��.����o�/Y�5��9��Dbw�u�u&Z�--j�ԻQ9�Ia�����tk�	�4���Ȼ�¨Q��IW���
ᄞrhejA0kY=߲�{�y;`Ȁ8$Ze�B�u��ŵ��oNm�#u!a��f�����=���p�DA�dF��-g����U��]���/�y�Ԓ�.8��ieci��>�K�����Ww��$�}T�o���*��S1�뙬�vo�6�Sٟ݇�N�O��G��%J�]���窻9�ʭ�I��a-ҟ����Nrj�ݢ�{Kg���`<���;[9�R@��Сy�,$����-�܄#{T~�򉰺Q�t��Ok��ys�ꄼ��)6�4t��&�Lj���,}1\��&�%r70TN�a���D�&TΈ�#g�r������O3R�(�"�0@�|��&��<�*1��غ���RQ����I�<�����56�\)�ٙ��������!3J� ��J�?�֩�	�UO^�$AC[��  ��,��a9k�(lZi>Q��h�`O9���6J7/�ze��m����S��un�i�z�cֽ�������Ըm1��@�&��*��r
ꖉ?Eu��S�t�) 4d�T	�x�hb����锍���P�X;��7���K��~�=~�����D�kGʖ� 3}��n�:��$�j:^�{3�A�p�z>Fj�̢�W\��4.s]���(�2}=�H�EzpM�� �x���f}��f��-����l������g[�JEK��9�-F�:E'6=�#.��u���gfd���)"��ϻ&���T]��v���WD�]ft��?"0^aי�='6�o`��V�� ���B���q)�$-H�*�H<�/wX����7�g�r��b�3\�_��Z0�ނ)�g�&e� p��.W#��O�f.̈́U����(�Wq-d�cgS�uL�Y���".�'��	�z�X�/8炤�QX٫i��<��鯯�p�/�RػpvJ�������ԭ��.q=�m�-O��`Uzp��{B�ު�`~{n�( ub�2�)��0��b��v�x`�O�u=O9���C�>�=E��Ց[�i�����v���4��O��Dؗ3N�1U�#�)��k5���]�;�*qW֔��7'�}[��(D�}�ǩ��>	B�-R�Y'�)�y���-�(��mA8�4�η)�}��G{Ve;
��3��#6��h�0j��_�#Q$fF N��G�(;h�m=p�
l6+Pi?[�C��
=Š��
?���2Pa_bi:F ��9�;&l��:je+ ?TFb�O�E�X�*�����2F�#�$\�['S�nn�0�oi0QN���q,��w�E���ؖ9֬V�*H�NUg��[��GN;[������K�9�od_���L�o@���	�H�� kh$FS��D�f�j9>o�FZ�p��Z6�yF ԗ^�n���ȥO7��1��v|��=�_��K�i�]�LF$��v*���!&P�	���������\ )�����46�>I։�1�Q������D����w�ͮP�
�W_�?�Վ��~;���ca�.���m�=#N�i���KoȋCz��M�;�`� G�Fb�Ӥ�A���l�	����OT��>�	i��t�8`���͈-@^�!�y�^
��?yR�̾�@l��,�)q �� vے����*j:�mz��/��WODd�\���q��W���n��Q�MX����$�`£2mp�f��
��af������ͅƢ�����F��=�s�\�$�2������������r����ei*{�4�[$�
*t/p���
�, �a�(gֶ/�*\�y)��,Xi��t�O3���h>M.J���9x�%�����^o�lv2��!�A�R�A���?��"���1�/�'Ҟ3xگ+õ릛.�oR;Z�{�� �Xz'���܆�ca�I�z�U�/�5�g��,s2+ο��U�HTÈ3�|�j�s�زQ�==��*9�'�jo ^��ZjMPm>DL�r�mo=2�F�U+*���}��l=�К��$� ݺ��}�׮9	V���?��`��m���ȴ0\@|S*��g������v���o)�u���+������7�Tt�����
�4�!�$X�2�w8�E��X��)��h�z���h�[����(!ÆS�)��7�`4Y�1i�W\2�!������8����0���x܂��C_���Q�˥D�$6���)v�N9KtH����	�FA�5]�R�F[
��;�L��� ����s��E�;�a-�ѧ�S���zߝOT�����u8�i��o!J�j��]�I�q|��p`[��²W���:�t�5	���kS�X��w2������_JV�&�*G��v����r*�l����#��
��8����K��˗�\(�WUL̀��'�Q �K-�\��R�v�/}ޣ,�s��G�)�3����1�VФ�|�#�ۅ���L���N;�5Rn>���l\�m�7�w�zN�:���.�E����y,�\�ٕ�ԡ2d[���^�#�7<��Te\ҎO�Cd;Ǻ�xA��2��]���g���淉�/��4_g;�A�75N��{�����������x��i�F�,�,Nu����D/@�����U�⒯����/����y<�[����ξG��p/6�(��I:E?��L�#�n�O���3���&;&۠f����φ�E�}K͍�.��x!i�4�4O8_��_`�UR�O�Ȅ6���P�^ܮ_�PD�	R3B�r��N�b�b�r]��_�N/��`�Yv��ϭxٛΜ
 �ژ��5�Z�C��d�K�����E�Tި�`jOn�Y��R����Qu��S��6�Ƞp�y���B^�!�P�XZ&v-�!U�6��S��-�o�ѿ>fڋ�O0Z��
���*")W|$fr�\-k���������P�x�s��f��K[kc{�����5�$�(�.�*Cr@���
B��k�V�Vlb�ZϤ ��nX{���o��b�P?�(�w�9F,�O6�;˰R�>Nf�\,Ti�/١�o�A�N�����X����y�+���t�+~1`N��^��N_����,��.]r%�p1�`��M"k�!�3�#o�C#[�	�5s�}����bt��LjA�ʨ��|�Z~IB�����?^���g���^��ɶ=]b۶��Jd���i�=����MN���C�9 ��w�Xb�p���p Wv�S�(�����o�@�B׋��6���!d��KQs\� y �������Ԑ���q�р���󋋃3Gg����Ě�E&?�L</�,::~�g� ����Mh��b��S�|�z#��^���|˿��g5)z���싄�Pj�KD�R�g&�p�|�Y�apdBMY���{�S���B{�U�TP#9��M���^��R����n��4�)�Lfc��z�!x��v���)�; ͣ����v=i/�����VUZ6�9�X+"�mEt�S6�\�ᥑ?����5���xۿ�ʏy1A����_3E�T z�H4su����Ō4�֌;ۺ.ϊ��cG�R7�U��[�{�����@9L�����?� S*���N�[����Î��sv��z�܃�q�;2�x{��h�t�/x�u�gď��`|ɑ�!N� �|G�'X쾔QX>,OA-�+�c�SGM���q���Z.�G�o��+�u3�DO~�ׯm���q�XkA7��_!�'m	���уNDñ�p�z�,�%�NC�KN��/4�Qz���+ZJ~�%�йG�C�	ʘ=ti>�W���d]��^n:Q�'
��[��t����S5�#(
��1�6���s;�n)�Uk��x���T-���@��k4lt�q�=�q����!�G���j��4p��f�d���i�4Y}�rs���e��U�V;�^��xu�f��! \l��N�\P�ۆ��� ���Kd��mr@��~�J�\���/�G�?61��mO�_�VF��?����=�Ije���"�z�
!7��/�r0���x��۶%Ѱ�怌v :eQ ���}�ݻ���~�u���8y��KJ�C���߀�:��_[��+���7��j���H��� u���u_��{��ޒd�,��K$��(��3S���t�ɸ?E�!�
�<�/?�g�b����5Sk%c�H��u �'	�դH�đ�$FG�m�����W�2�iyC��w�Fޤ0����r񻵺���9�� H%�a���W��8�Ȉ,si��X+'!���F�j)Y�ߑG�p.�fH�t�G	J-*�;6?�� %\�z����2���խ�$��U���SPc�v&of��hZ��s� �×�=l�T�X����9
�P��$�qn]1D���^*/q�s��ˈ����hN���:��_:��9�Y�L ͕?N���b�4�ܙ�6!ҷ`0y-2|��8$����6Ƽ��!��Z�!�Vܹg�"x�v�(��P�_�;r��փ�/�'�����(�4��;������t�O��~mܣȧȿ�'����%��u��g��>
�#�s5�@�o��谤!���d�Y���ސ�6a����M5��	L�*p�]ܨ^d#tf�`����ܧQ\�*��7����`�l`�NJ�&CM���R�PGM����s����SW����G�I!����Iazb�$�܃����~A�>���ވQ�[qָJ���$�̵b��
�G�����_��cq�2?%c��:|��C���|B�_��Yj�#D�2#`e���\+� ���V2��&���o
�%��3��C8���⿗[+Ar�yd�匸��� �l���&�������$���R5H˕�ę�r�HH�NS��k��I8n���--py���e�MR�2!7L1?�3i&U�/.�`�`r��a����prN�[�_��a��.��l���O-��*hr���N�8#t����"	Ц,�S�[h��N5v��#Tw%JZ$ I�~/T�,�Uڏ��VJ��?EQ\����O���ՠ��D�a�� ����i"���
>��|��}|���Go�����*��c;�.���	�.��Y�|��[\RJ僲������]�B&�t3��p�	(:l�8�̩#�T>�'��c<k�����p;o�����S�um쏆���ݵt[����춘���c>������;��1���ꕝo�&[<��<��mP�]�bNK���?��w�e5F�*Zт�<��Pl���� �<eC��r��K���kt��_��P�Lc�\,{�;�z�y�-(���i^�#`�ch��t A)�}؂Z��A���^'��'�Y��<���~̼���	�����o6'�<��".䵆g,!���@�u��exR��ئ����=2�d���"�f�<�;���k䗞dΎ�$_�Y�6"]��/8�.�����*5��p�)�3,)@�"W�l`�\���ΐ��*x�V�lQ�2�B#f�e�%���|��N�ղ���|;�u��Bz��6���䴳G�"Ц��U�<�~�i�%���Q[&��t��n�g� �W�A��h:��#B��R�C$e���������T�W�����(���C�Zs���i�? �荰9�����]�Vϒ�j���������5�CZIZ�,�.NIY�iZW���7e�M��N�M:�jd����W��FD��`��ƂC�����y���	�8CuP{��cޡ���&2s��@��;s &�9)]u��B+�ۍ�P(V�����+��_hbP��ھ��fi��(Qn���A�+M|����^\�`DF�;��C�t< Fj�c�����({S}�5$���w�Q ���B}43��)��5�4Y[4���"-C��)��D��t�qVK��B����K>�b8��}�Հ71�߀Kbl���S��D���4����d���9��S�i�kq�I��v��d�E\:j���f���SM�P5m��+�DBj&{-c�A�o�j$���s]����;-D���c��}�WsWv�3 ���!��0�HN��QYf�ᵹv��i%B\�O�%���#0�eC\p������P��AS��ėx�D�x�R�Ў�Hj�^  s����c-ӱ2��b��y�r`#nsS��<�*|�Qt��(?��`}�zsJ>pZ�tu���{�����IC����o:��0�t��n�5U��!R�V����#����:��¸N�JDG�L��tv�6���c���D���h&F�j[�?&V�=m˝+�RPD��N�A���be��,��1ǺJv�qXX�����Q�������\���?��*�����Oe|�e���2�*���V�EKY�ದfR���N�� �(�����ARR���8��߁�Ѝr�jZc*�[u�Ŀ�A��r�?�����&*�I�JG���|��5�`���`X���٬4T���b����Ծ߬ҀXR�^��N�w�1P���;��U���^,�p"�-���@��n(}����&x� �u�e�c�8�)��a^ڛ��"��t����fs"��F0�'�����\��b`@�XR��+5��H�?�6Y>�u<���[���=_녁�����6~Q"��Q��v*��	43�%Ʋ�s$Je8&:���&�Ƌ2g��'��7�St��9H��
s�������s8�2H�����wP� '�@X��!�R�)��X���#�v�V]!r#��'|W�PE6�"/�oU�}�_
�����Ku�Y�I�q<qK��Iˑ@�p�:�&�h>�f)U�.(����C�0O�DM�>D�7}h�mk3VL�"���,�N��ȫ�7��� ��?�.��
�2?}6���Gm�����ɗ���G�~�J��k+� �_�<_h�)&bj9;$OOz���ѠFB�}��`��3����O�⫨�'��H��z-D[:�p�Y4�n��Û�Jb��9|�����l5��L���{.!|ݢd�t¡����H���:���;W<g���
O�afU(_������Cf�@q���i���c�ͩ�F��:_���+������&�[/�
.�_�l�ˍ�q=7�e7��5���F�7���O�["I���-�������ZHA�.T�|���.у�f��c�˷���x�N��{`���By5V*B���s^I���vY�R�단�H���EY�7���N�v��}ȱj��x�:Ԓs�0���hPa�ܖ�u�N'|�	p�u\��~Ňݽ��_P������`^�s��p�}nyp��+��z��7��=�.֔��ձ��Xi��	�HlF�RJx�^?�c�h%?{X��@��>iu��4R�4���j�\6A��$zd���|֑w�bLȈ$�}9�e�@PL�TO�zx�Kx%�w惀8�m�=CNl[��������@n�j��G�r���}�^D3�4=y_�Ō������4b�������r��������������v�5ɬ�U�*"�M��plG��դS�E��n����5)�"1��î*c�E)H��s1��� `�P�9A.oę7���ۃ4��rJ� �n�q)cCpM:<��
��6�!L��������{��F86DھQ�g]����g
�����ԅ�U^�3�4����#��'|� T?O���A�Wu�nN�f�%ӗ/�+���z�*i ���r��b�)sޡ@b�.��U�N.ےn���9�D�~hK���2��'yV�-J�F��}�Cn K+#�-N�mAU�/;�-%�VȌi�1 �\_.t�����4ע��:����>��ڭ/��K��,n؏g�g�\���Kٙ��K���{);}��2��0��`�����@��8��fG]�F5��P1�Fq��e{�}[�ޞL�[��5�@a���6�^��Et=/V���a�\g�fV�䍅���H#ZJ�W��_���̵;���-"�:Z�'R���c.!��g-S�؂q&f-t<�� P\�E)7���E1`N=�����g�c���t�RZ�[R~�<����5��q�X�R��#C@��F��+Ay���S0����E�U����1T�󎱣	[�)z�``�h�C�8�;��~c�G�D��Ry��&%m�EIoZ���XFxvG�����%�m2+nk�+�>r8L�V�kVN;�T�U�0����7M��j�℥cT7�g{����Wr�&v�6G�e3:3t�1�+�a��p����*�9�>����E�Ij�NXI!̈�aa�`�x��X�������\�޸%���:�B�bX�rߧ��A����T�=[Ͻ�G�T����%�Y ��E�s�4>xE��d�~���7�5W�Y�9vz�˞w���$j��k��[D�~0^ySy�lف�|�*6�z���+�MK��#�����zR�R���qp�U��S����F*�F?rsOSV��m����sN��J�f��Κ4��,� �T�a�~mN��
]�&;N�]o�4�:a�x�|�4e�����2*��P����yP $&��.�=TC%V�o�K���.�!g�G��˦l�/��R�-�7�7vf|�P�I=�g@nPz���I|#^�,��Rup�{X�|��ԕ� �6�T3�ǳI?=�h=+""#{d�{�^O�j~���SO��{J��� 58i�����:, d�Z�vZJ�x[b��d�=o�f6}�o��wct��`mek)�Y�[t)ָ�?��&ʢЯ{�)�vYL��%�U��M��w�$j��|�(٩U�A����U�Y��<�UYq�Æ.Mz�1��4���%VYan{,������+/��	���4�ʋ~�}t��.���@���A���-�'3�6&����P~��ȏ
�����BE�^�6����OIm��?K�q��.�"b��� `Tļ0��D%���-��������e���"q㳺���d�:���5�}7҈���\��fTah��+- �q��P%�hk�! ��� ǹ����v~�R������ao�Gbl���K�w��
雇��S�k��D)�>s<1�%����j�ʹ���Hnʩ�{�tf���?�cy�iG��8yA*]��Kz$�hQ�{އl�(q���$)/��<i�C��t����H��<��,���/��雑��F��m��lHU�
Ftب��=�J�i���G�kB�����
�L]�=����*:FF��)��d�;iIV�Λ�k�"Ï��n�]^P�ݗ�����E�Oo�~�?G���������o�2S�އ��/w2����f�����~d3Ͱn�n��C�y(=3���n<+�qd�y*��� ������Rs�Z��nxc����l�j3g�r�M^��'���FM��eG��Fe��>䠹���3��O܋�(+�h��h%���?�n��V��p<GxV�W������rW<��O �̀l�F�I�K��Zت�A��>Ad�ےuv�^'BBo:B�v�J`Zn�!�-ܡ��5
��F���nc����dn��8�3b���??|�[yTѯ�X�՝IJ��/���1�*X�n}V�Z�Fh�E�\��Sp���9���P���}4㷇�q���B�+�

��.�oO%l�,��h�����"�p���3�*O3�Mө*ҍ�fe��}�p���O<-U��o���8� �qˣo��K`+eux�
׸�)S��d0�]L[�5os�@�㋴������V���4%p�>��ѐ4�_����жu_�&Up�1wb�9�7�S}���	.��qEO���{g�5���q$胺y�H
�&y��:����1�x�h<��X��4�>09X.��v���~�NPi�;G*��� �bo
\�H1j�L2�94U�����^�c����'r�%�C̕������ʳ�X������A� �j�����9;5�����Y9�Y��1��<�r�T��*t/��a�@^%xqeKa���l#���<f� �i7����z�m�0����r<�uJ6���OYQkي~��ݓ��
~f��vUt/�д�5���E�I�Y��0`��4W�������X����e?��a�|X{9E�H|K���Ql�_ VO�]d��MF^����?ƽ��"�#y��$rq-���Ƹ�)��"���s�t\�E�46>�����S�!��8�����#d.р ��(�� -V��מ�
�NW�#_����P��}���p@p���$j]��ᆡ�0d(��(�g�p�������j��F��{�����'���(�N��2�Q�ݏ���3^��^�@D)BM/�h��~�F ���I��z)C(LX��_d��ZQ��_��EfE*I�T�����)�f5��G��ܧyK]�!R�K��M��n�NMH?���tG��ד�f�S7&��:�C��������Z�J'���~_q8͌��O��i���'<h��^ov� ��ǢY�8_y T�Ǹ~�?�I��� ��V�N�b�Jdþ�X��n��1��Z�'ܕ�K�>5��LNv���8aOd�E ,������SY�e#�*D<�������	7�2ͻ�P�a�mx�G��kd���2�>�yz�?Y	t*�@_�P5�w�=Jz�(I��;�� �3����ɞ�e�'ӺE�.q�F�pZq���Xsk1o���c�P޾=��-E�d�r^~�vǨ��
�(�C����@Y�$\w-ym��b�J��oGE�*M<�f:�Ef�5�g�o�*�c�S�}xA�{T��2�a��v[�d�w3ίh#�9�#�%�l���S7�L���sGt m)��C���H���*պwt���ބA���2�V�Ơ9iT�b@��# �5P��
r(%������.1��
Z��+,�hh��;s���D��Gf8�?fɣ��;�X���h��lF�c��nۉ���;j�6�����oe�wY�7���f�T6�4�M���Sb�7�P#�u�2j��n��̇�oj������?�[L�-���[^�J�V���y:��$~	F�:������ �w�[��U���q��ƽ���:��dH�9�72M^��52��N�Z�M�~"�/D�0?)�ת�A�\�`���V�n�(��"p���_m�U�J~��l����?�W���OmU6~W.yfz�ǓR��h �\���!���㱧N��T��o��U������8����9MЍ�٧O�e��̈́�!E����G�k�8�M�L��ي|=��q���^��+c�.1���GZ��ĸP�G����̚I.��~g��B�˕;�y�/'���%$_�w��5�R�4iJJK�x=Z�nOP(F�216x��ת��t��z�����ra;��&8���ZK���/�R���T/��c��ܫ=e�W�x�+��7�v2Ȧ���ށxb+2�� M���\���F�N �/�Wo��z��T�О^I�qi��Y�����T�k)����o�߼�#>���(j!P��Z�xе_ψ`���޹������"-[�[ު��9����H*0�-Nf��]U��IN�n��5:M~+Q��j=jl���]��h?�#��� ��]-���1D�	`�`�}'���g�c�C�����LQ�s�|�_ >���4�R�t�1��9����`@��&C��%�/i"Lz^Is�7a�`QFYyzK�Y�(�
-����hk���o�t�^�����R�4Q`�,c�@���))�2������h
��jH:},����. �S�>�������SI�Ʈ>F�����n�g!*!ql����n������������4`�fr�2/���]~���齯��b��ʱ����[��d�Q�	���>���auT�ϰ�a@yVg������>Fȸ�+vK`�h���_+V4*m}�^a|[�3M$ڮ=,�ցO���� �z�̮0�G��H+Dy�r��� ����&<�,�Z  1g�Ө.i�k�_oy��HW(��?K^�T���w����nm��o6�f�آ��M�Ef��hw�Y�Msvh��6�:��݆3�>�.t���~ζ1�g%$4=JޛFUy��x���1@���ː�qV���GCz�������w���E�*m���P�^��\P.'^f�11@����t��'�f�q�O_�=\�~�!��4��*�ꠘK���ExR�Wτ�T�>��B�M��=��jۍY���.����AP-}a�?l1�[(���ʙ ����D]�^��Z�v�]R�ۙ�tA�*p~��Jl����������?Hu�����ǔ�[[�kR���o;C	$R�!؅Ls�lK����Gu��ގ�3�E�H�J.�V�^<������xlj�����fb�g-q�EL ����!�d����o����&%��|Nln� ]�x�P\�'@��j<�V�X���o�RHc�D��82���b���%n�M��$+?���4�������0�x[5"��ͫz��gu����1.�%���2������� 9%j)<�@�%U~���/���.U`ҘAӵCi��I͋Sijz{yK��8�x� �i.m)9Er��A^���#^)%��siy &�&�l��6�p��޶ۿT�J�)hx�>IE0���ݵ��!���L��KTo[�+P�cy�w*�s��0+�5�o6���&D�����$dFl����	{��Fa�U��#��y����[�T���7xLa��K@���ꎢ���ɔ9|����g�|;|��>�3���M珿"��U�3XΚΥ�>U�q�����S.?a�e�Q�.09�%��W'�p:�-����n6>��A��ݴ��X�)9Pm���0�_����1p?7��2(
����t�f0�X�������U��CO���>��Ѣ��~፳}+�nV�u�� ����z��p2t+{�ޒ����M�,D�=��е��:�g\�a�w4�fʥ�2�_�M��c����_*8�����qwp2.
��	O(M��C�b!?5ZP%:�L��!'���$��Ɩ��,$׬3HE�3���Hz?����_�D�"�JA���|g)�\@�B�V3Q��e��(m�
����B(��=Ba�g�}S�&�«m\����5���@��l�D��.�$�h��#	 �kV�FS
8��ap%Wd$}����B�Xɬ;�7�����v�>0I��p@Ȑ���:!R�&_�҂�I�~Kc�����P�K'�}�*�h��af�Lo/v�=J
q�\Yf�A��&�ZfY̫�-&��7���� �P�����\�ǎ�=��R��!��!R�"VĬ �a�)��;�c��9*#��p���|fqn��c���*����}?��8�a+<A�(�Bm�
�R�OfZ�y� ���旊t��rѐ���n'�@�@;�y�+�0N��>����eQ�آn�"���o� �&���"���b�ȏ�I��#��;'��˒��TM�+���7�����0�R	�L�⫧���)�������.�&���a��׃��q"������l�ϥk2����@q���P�D��/nw[�y�\B=e�D\���Ұ��Zt��l<�����Q�(��Eqf	~��ض���Q����WK��9qK��G�F�~�}��q�8�b�s�LFb:^%�,3��8:�c.���7�E���JE�GJ��b�w�6-}-	�V����k�R������PZs��c�r�6�T��`�>\'l�-�IL���T�H����yj}�������}��[X��\�
k+uw|��(/�q݋j@ 6�*��lA�"<�(C��t��Z~sQ�L�Af�-4��wݚ[�S�����,Rw H{�Ȋ�s�l ���#��z�����6����2���-����\2:>]�=o�l�@�S��c��A��KB�^1+��=�g��[���Ir:�:]�9�3���A*���5����%�} �,S7��7dz�L,c���kgY��&����5��/���++K|�=�l1k���T�e�!=Y@�c��S8�{<:�hN�l�� +L���̦W=N�eO�S_���^�Þ��=�/ɜ�2����v/C�˼B��Y�~;��ud?�Q�
�_��*�������c0i)]��hl{����FF���z��*Ĩs�Y]�l@��E�۟�/���t��bw;+isb��A0}��]�-��u��І�\���*@�=�*t���^Eyc��%�z����8����`��ѽc"*fZ<��O��y$C���1��į�['�ꓷ[;���t�����=+jǏ�kh�������"�lM�y´6r��W\#��������YP�[�ۥh��#�9$f�x�4>���J�[�P��M��&��V⪽�헽�0D������o��<�� OQϼ����%��XREG��c�E�0�A�X}Z���o3�16l���e��o��g��K)j��;��A�� ����%��_��"�>��ް�©:��kk]��Xxa@"�[����'c�` ����&aV�3�!&R�hq\��Tr�Zn�DF��.|0Z�ת[l����RT��2�Q&4@�!2����B�q��I�?0Ǽ�` �&ر)D}B�����`�bC�R��Y����ɴ�i�|���dX��9�ΰ�cc���ܩ��d��:ۺK��d�a�i&��q�/���f'��8��ïS��(��X�k�$������h����d��D˩q۵���4	Uft飧�k��@S)uF�lGHo���|���?�?y����<��l���pײZ�f7b��X��r�kA�⁚1afc�� �:r@)_����%_�79p@U����I��CM�J �c�UR[R4qVscm�p�#0q���sҫ/���AJ~��3o�ݝa���������q�������e
]!�j�ίb�jA�O"M��(��sC_e��GV�*�;e"��q���<�95p����X-���H��|e	0t�vw#�l�>~���$Q�F��~�>W�aQ��:��>�c�7�>�	��&�T��󗠾~��6l?���(�&�[`(,~{�˒ѩb�Sw}����YQL���S����ڤC2We:^F��m��}v��&��~
#���ݟӉ>�U!����f�'W����jG�]+�f�02;�qEy	��!z.%1���E�|�k1_�}���$b~���K��̠�g�ȅ�#Q�8 �9}�`K=y���O��X��I�� �X �����#�%��#~%���>�äX	���Y�`��71$�6[w_�w�'��<��a�E�|�A>E]�/�88J'�b,�r1%��#���ǵ�&h�Ʈ�W�x؄ċ���B	���+�ruJ�Nf���<C��gV��?#�WXQD	�Z�2�(d?v�HE�e�T:���[���`{��['`Ps۳ʐ�m����dgM�}�)����!��d6&�1x���l檂ƃz=��ʌ�e"�/����D�6��!C�`Z4�R�2a�`&�����J�i#�����ߡ�F̈́|�d�WQ�7�R����������6��fv��a S�4Jr�rG�g����`8��l$��0J|�JUZɹ˅�5��M���k,���t(O�Mq�����BIt��Cj��m������`"�$�|/�,r%{�?��ql�W;�LK�>�a�C�����x5>z�e�~�^3r����W޳�DnjQǋ^�1�L�-}��rbX�Q�L�_�����M�Q�ya�M_��9�+#�A�p�`K�:q�=����4��\��j]i�0g$j���k�)u9�k{p�o>R�4
b�7{@���U�m��A����q�Rz]*}�r�'L��h��ĩ_g����)�U���ץM!L=G�|Y�~���]C�)�~��U\x09j��Q��Y|���>T�Nz��x�����ߎ���}�����y��U�%�]\�<�]�]	:��&�Ur.�������o�/��A��i�,q�U�=�e�������֒3G������~���a�)q9{�R���rS��k֛)���a��������%�������<��&��4 �l5��%^�K��.�8�fLE��6&ř�e+���/��<��|@�B�G��d��Zf�ee&ó=o��>����b1T�k�jk���$sYO9Ji~����vf~�g�;��z�,L���4�3�I�� /R�%,����d�8�(�Yye2��]���#��������~d�]W,>�w���:�=��ց]�	:�O��_/��ʺ�3c��;.��4�Ow?-�ɀ�ʾ�b��e�%�&�JH�[�(I�p�Y�Ѕ��#�uͣ\J����Ru,� �� T!ް.�Ω�d�o"ܮ��<m��ExW荛N��j�C�W+u�qo��>��	!=I��H �.g��;W׺�]S�����̽��jn\.�όo!d���V�v�?sKRl�bˬ���Ű.zhRYȵ3�B�*� +̳}Zm��<��#�|Q��<������'mL�rl�����T����b��!^�@nC��/D�C�س�ih�n9a��p�����8�z�#<����*	�&r���9��^�_�����l�s�xbޯ�A��tw]jA74<� �͵|.�����ӽf~��1C6(ذ���+��s�K9K��A	�a����;�Ҙٜ"Ϳ(&�ə�>6���8U�����8ѯ�&?d���pqţ�����y�ٙ����n��]d_���^�Z������ ��d��x�Hȭ��a�{��:_.��_��3�]{��yvU�V�W��w~0.[u,�����o���ɦ/1w�^�m��ݶ��sF	���bd�-k9a�)oé���z���_���qV#Mj��헶ʾ�SSRn�B1}��4���F*l����ɝ;���EjO��t�����X^m��3�#�ÿ|�Nr�&����^#'��l�]�QJ��������^ؒ���V�Z�l�I0��l3@�Q݌"��^z`V�A�b�}-Rf;8$���Q�D�!Q(H�ζ(�p�)�bh�	�N��H����R�W�tl�a���|�M�n�h�rl�!L��>�:`<�ѱ�DQ��3�]Ai3��Z����x��i ���K�#��qE�{�J�����X�Ռ贙`E귒S�{+�j@y $u�ARr��U!���-����C/�
.G�^6'�ҡa8��ZW'�I�T�>w��
qC^�z���mѷ�j~��f ������2�<�Z҉(u���9��4�4��-�!���2|kIަ@���ڗ,P��t�w�vx��� �td6Ø�����!��9~�ٚ�(���W�<a\�j�r�D#�}-k_�	U|N�S2�P���Lt}Z:�z'^;�yqȊ��o#�!	����4Zh�k�E�27S璆��eѡ9lk4H3�La��ϝ�^���(�C�6e���`��cDI�`���T�!����l/�%�7g ,R�mQ��a�²?;*v[P�Gr�^b���8���h��ߚN,.h=Sڭ�v �l�u�}Tm��?���Ս�e�~��_��\O;-���ࢡD�*�v7x��[ʶ]&��o�ޮ䝒om}�$�6)�6
����Z�p1�b�Ȫ�Zp�R$g?
����jE��1��'8z�kX{w�O���X{櫘�nO#G�-�
I�2��Ĉ�#ll��I��;2�a-[�yn� ����x�*�){�����hQ�we�Աi�1+\�b���1t�k,����=�?�C�'70��x�<r;z��P=�����<��yP�Z����C:*�.�`7�|������ʺ�o���4�7?9>M*9%��9kQ�j�]�F �$��J�~�S�d\��%����\BY���[W5~�p/�5s��a+q��ht �@'�v���v��' *5���cF��J)�>��������	p%tG����+c;�[�K�\L~��W�Z����p�<E$Fhm]��u�]Iii�K��t��E��r]��	��B�	�+��L��*0ыy_6�J;H�|*}�����K�gE[f��7�%�NA�h�WO�(�k����f����)�,}5gs�P٠q���X��*4�e���t@�}�ш�[�$�ӌQ�7Z��K_���#�C \no�'�8A?����Zm^�M�Zτ�����*ޅ4f�t"1)ѩ�:�F{v���ee��_�J��ƬvP%��Gj?�qQ�@��\I�b�^V���n��(��vO��b�9"�����jSM>oL-�'�#%�,��X������Pw��t�S�<�ڋֶH1�G�ss���ϥ�t�X��-Q��E�8v{yݖ����E��e�ó�|	o�|�W-���
�/+̵&*v�.6.�j���D�/�-)�EDRi�=Z��:��\����-J���5bz�EȟV/G`AG�'��H���j�۲��Oŧ�	T��Q�GwJ.~����bC}X��]%PÖ����Dkl�@�^~-�����[��)�ɰO�x�<8�x�9�c��?�|�;ņu)[�~���P[��>" P�S��jb.L*t;i�62O�F���Y���M�1��N���wTp@掩���Q�b�b��o�|3U�t.	yN`F1�#j�X+�<�h߶����d�W�#f�+�цjↂ:�|�9�j��B�����A�<=W�^Xȑkqxݥ�G��F�XD��#�pe�R�'�^+�I
c�ѩ��gG1��$���~�e���oɔ2@S[E	i3�7�H��YzY��F;&,��\yx�7��C5���U �ܳ�)N��[�
&I R�Ë1�Sގ"�|��ZcG��2��h^����e�+��r�Z��!��2�&���N� ��J	��b�I�)�0�}t7�.W��|�G܅<��v?w�]Ԋ�nBJJ��d� ���p5�"*�$��/�����g����~<ɑQ<%��ck�A[iz���5/|��ި�K�3�Bfw��~v��-ջ%=�C�IN
���	c�01E������uz,�+H��@���B!��=��� ^S���L�y���ʎ�X0Ԇ�4q�eڌ �����2�B�X�4v��mX��x�OP�ŇUױO!�&�25vf��O:{�:��#�"�\Jc�7���0�6�$��s�I�0AQz�i����;���AB�f��{�}��JT��XU[O��k.^L3�G?����y����8�m����§v�2�2��V'1CL���V�����AƖ">a(���eW|KI�,�b�8�R�Z�q����&�ĝ���M�g�TJ��".����>=B}��-P���ф|�*�����Pe$��i(>�1����'Z�Mo�S�G������e@z{a����%�lSʚX��M&^8w���L4�et����h��
�����-?��-�件�i�������K�"�CcmG,������aO'�6<��mo��@��X�Hɣ�{@�r���ɨ����xR��V�-�/�"T�[����n�VWq�x#�R�;
�ry�X��$�)���}�:X��G]䔅�L������K��k�%�a�C-.Q��^;�@78TF�����ż�����N�g|�уZ��ϐ=�Xh�3���,0��"���"�]_/uD����+�6�@tI������ꡱz>���N��kƿی39Z�v5��%p�j���
������w`�����*Kc��Ae���p�>M���OIhZ�ʲ<���?��k��1[E���b���.X[�S7$��{S�j���Y1@������V�
�H1R_?�6��f9�Vzk�L��gَ� 3�m�b����u�j9%��jBS�^��S̮io?�̽}<��� ظ΅6��/�ԥu��'+J�x�NG�9����*�+n�3[:5�"#�C�|	�[�B�n`?�B�M�-`�4���^s�����;	��	#�a�V��G���4����j)�Iu��r�s�Am	rE:� ��Μ{�mKbO}�
7/�lJ�NF��يv=��/'�g*|	�p����S�i`(�m��O��b��2�P&ں�Vs.ɇ��w��?.�B��g��-��u��'s4K^��T���.K�u.}h�TC�ޫ��*p��"6t�0e൩��"g� �gOn@��i�""1&_��\X�U|���sL��2� ���7l��M��G��n%@�O���݆`]�'mu�c����%��+Xޔ/ġ��1-Y��%�0�\�0t_�r�2l.�Z�4n�p`�']8�Ԡ� 8:B��+�G���R���i�Yߵ7u��p_�{�{��ǩ]�b���kذ�Ƞaw&�*���;�+�����1/_�Ie�h@h�m��*��F/_����m�̜^�uZ���B�I��M�D��p�n!��yn�Rײ�h��n���2^E����
�z�$9�׿������h�fFI#�yuטn��$�󉭁���-	5�����ɾ����l�*�=��-�W�,�9����7���E3��EL�2�07fL��^�@��O���x=@O���10���i�����]�?qb!�o��ǲ;�(dN�O�ʻ�(�����7=:|!��R_o��v�

p%��D��[0�����������
�D@ ��-���PhS��ix�����c�	�}e�����	h������<�G�^�N�4碾ܔ*wOP�T���\��(�4�q*z�-,ӿ��� p]�8ۤ7cK� h7�lJ�K��o0P���@.�%�6��/�n���H�,���:n��9�����B��l���������(<�*���P�#�l���>$ �bk��y[i�����Jo�*N��l��P��E�Xv�0�TCc�b N��������B��f�^�dH?,��.�"�U�XI�n��5�� k�X��P���'���t�n2/IC������0�y4 Ҩ���p���b�ռ�B���,�|���b%7\J|
�E��c�L���H��~��|�<�����4RJ�o�bu��u���Qf#+iA�m\�C�����؋R��i��N2��ͼ�o	�J��d�J@�^���>��)�NU�W�J���<�n�*��6z<*p�E��7弻���7\���Kj�k`}ܬ�܅�jL݊9����r0�t=j#�ƆUs�}vR!��c@e氛2�hq�����������3!l<׈�r�E3E{h�L���LzX�y]��,��M�>դ�X~�~̑�9U���ћ4^Gf�4	����$��|M��u᪜7�5���Zg�ǻ�Ջ䖘��p��򾨶7���LѦ���q�CKb�H~a��<���^�US2Z�{1��0�vo�F�S�2�V�]��2�*̓gsC�}�JZP
��m�W�'��1Gа�>8���y��hm�����t��_~G\ke7��X����)�&�D��<�Q�JNrdi��m�����;0�>D�`����Qk�{�`_����_t}����e����-E��˺�<�-}�sggD��uҏ��Z����t����<1��榝P�'��� k�����"�y'z��Iz�#C�G���*��	��X�C,�@A�9oXDIJ?
��l�%�S>\��M�ֺBD%���ߓ\Wޑ]�@���ފ�q�"K
�QQ���tc�<�h��ZX�.��MFy��t�^C�.�ᘡ+Ƣ���˚�8���:$�n��G]A81��(����+lx�Ϸ��E{�m˜�T��fQ/[a����;�b�n"r#�>#�^"�h�s̢z4 4��CtZy�\DɌu�%r�jky���:	b_w����Y��'Ce/B�qU%�MڒP���<���J(�C�����Z�<�L߁��t@�W_��ӵ��h\�Z{+�9�޴ ��w�����J�,�%Yu���d��s6]�l�U��x ���+햴��ԃ�+m��W��־��ǉq�RrQQ��O�?}�/�\M�7�-��.�B'l�`�1���B#�!�ϳc�wr�J��A�%���ߓ���q8a�=����>,O���DNa^��E�,��H���o�b7�> ��:Dl���s�3�8�_��vtHK5�%�;�_�/�$q������!�{@�M������s� ��1.d���l��5k����Mv�[����禰�	E�l�.V>_.�6��^�'��e��^!]¬B``�&����h���,�A�f?��[-D�b0U��� �l"6Qiz:=ᥙ�jV�d^B�ؒ�3ృ�r���ءn�r�`��}�m`�.M-x��!��(�__h{z_��j� o���E�.i��H��N)����54t.^�cU�h���".�$u��y���碻��g�n޽1<�wSB��'���á��S�N��C�otĕ(�j� �J*��_4�+g�0�P������ r�i�čPB���3Y ����@dWС����lN����q�8ݙ	��e�<��s�ޣ���$�f��^���A(�:��z>�1nz�e���*J�8�go�>�s����l��@L�f�W��&KZ���Y�%�1�~�����b,��@������)�s)V���#sS{E]��Tl�U��K,�O����֎�O!*V\S�h����Q2�%�'���G���N|�������g�!���'�I�G�����)�'�MhG��������_��K����y�,ȕ�C*�l����E<>t�G\ �ۑ�"5OK����ˈ�n���ՙĕ��m�U�C9���Һ0
e��z����#=]@N�묬�/r�����b*?w�L�p���y��;T�,��p&��@T�D�3u�B�I-p	I~�,���M���#��v��$>] ���dv2�G~���֨��B�_nO*�qH_��/o`��+�ݞ��G��Տg��f�d��>AH�sz�ڋ��DϤ6R�*q�>�����v������ r>��=ɜ&�%?�cV\�t)1� �-/�K6��9��� 'BcmA���6%����?��[�_X�Y^0��P�j�3�5��<���!;���x:�G�J)���#��=~�=m��0��A���=��A�ĸU�1�ou(1�~3fc��V�[g�R/���6=TL��r�s@�^c���S��a��]@=*IL�m���d�-��ҡg��%��=p*J
;���u|���Y�m!gB�v��N]T��x$�����J��֎�IR1� %�u�ل}g��p�1�[Zb �+Т�̇ҩ�H\�Z;����arT^"�)������7�d��*��k�,��2a�i�헴���U��1L����)/���uL�8rh[��S�Ea7��j��z�ⶋ�a����s[]V�E���b�5o��8��	[�ld�<eќ��I9i�Q�3���	��I���ب��ݵ ����iԋ�S M4��]�u3,R�B	U�������Zۑ�:�������oK ���rNYK��--���؄-m�eav��S���8@L2[�\�������&EΨ�%-����г�'M���:}��EQ�5N��v�����>bT�ưl2�$�F�*Kɞ�v��M��$�*���1S���?J6�|�~�,�(y04݉��ۭ�,�UT��*��������)�|'�'���`	~��������c�5�T�`h�W�t�r���J �%%���&2^����� p
�����ۿ�Eo^��@��v^�cb�5 ���v��E���~}�Ð��'���$������� �@�����	Y{ش�i�>�A2�V���GI������7�HS�T'��W�**���J�\ @����rNoa�7>�,�8��qg�u�������VQ���ɫ`�
�@|�북�M$�7����l.*F��.���C2�4{��DG�?|S�N8M.x��)���՛q�hHEFH8"f{l���!��؇	�Ӵ/9�U_E��?�\u��O7rG��F�T7ef��Y���R����R>9.*ԩ��C�T�H�
01�4�<R�-��:��Q�E������4}�*j�4f�d�3��+gW+�'�I��De�}!��QdY����*z �
dh�Ⱦ�{ٶ�>YFC�W�?%e��Kg���5;�s3����������M��kDWU�o�|"�3��3� "çh�^w��M��G�B��&�'jA��ϛS�д�~_������$ �F|(�R�&a�����:Sř�F|^O5Y����x4AJ��a��1��{6�	[�\g�������J���M��~�"����e��[̻?Gd�U���� \����I[�����p��S��*$���՛z��O�:�Y�a˲����ѣ0�#ݢ��b���6hZKd�t�[�/���C&��Ѷ��԰��A�s� D�!�@�6�x1���x{5rV�f�dS�Y�m��x�<F�&9����h�j��WA�K]�!��P}8:d;��;���N9��a���������'�o��X��*
�����<#�Qo״F�%�-��d�wi�#�.���?���dB�&���כ'�XJ����������k�%I���s��=AY� 4���G�>���^�,Z��(�`�|�i��7�&�����]-O55"9c���G�%�n�q�҄_*���a�����~����W�5$l����9���.Hp�3A�l,	hG?>�6�q ]F�sf{d %f��8�xFC��i��7�w
�x�ne�=��"x�ܑ�a~�X��&2쏭}N�S-v��0��
�7nH���o����SOK���A�F+'=p�N1��m�����
���V���"��:��q'�/�1����g���'Q3�J�'��B�i=S����ޕ�.owڐ�d�dL_� R< �~]�F6W��S�{��xUM�;���+j���,$����� �e	�)��^ǒT�F8o�d2E*��ϟ�pIP�:qb�8 X`��p��{��*��	R	.Rx�#+������﯍z�Q�&�%�U��S�� ��#�%�/��۷��
�����g4�t�"�#ϰ��Q��~�e�Һ��i�����7�G`����;�@� Ҋ^�1��z����_���nP?��,�����b�.�(�t!��;T�h�$Js�CR�-�����6����)&�M����[��׮Uȥ����Zuv-NW�5hI�䢼�Q��w�/,t�k��s���P|A�I� Y��[�5FX �<WM�~bGo �W���io�7x)!"cZvp �$�<�_�D��)�^d�`d���x���-����p����n��7ܬr^��!�h�$Pa���Z��(	4I�cL�+b��>��sɶ�-���F�]Ĝ'c'���hL2�(��W�q(�[\[&6R�?�J@�}É��D_#��������,4���2M����8@g8�~j,����d�m�����8'h�M�)�8�/uk��x��d��d_����H����J"(��7�b�]J����{^c�Wc@�_���u↾_�<<����d�����Y�e������"����]Y�S�*����bf��{#�=��8�*�2�m���K��` zk����b�����r�߸��:���0j���m�L�a�ˍIs�u/Q�8={�x�{��6Z/�-�'%���DR6�]_�DW�c��X`#5b���'�p�5pE�E��4�$�R�p_D�-T�{���b��;��RB�jش%�X226˰<�m��erQ�'�����&W�@P��#�u"��D�U(�>;X�֔杀-���Z��)���=��t\��2`z>�Ío ���^���)gqxߘjY��?v���Y�wŠ�WK#�3�	i͢�����n����=�e���X}�`յ��g�P%�51i�������`�����6P����g�@)��Hl��%�c�R�&Ai���Fc��:v�Y��I̍1�>�[�Ҝ��W�Q��5��)���L�Ѽ_�^,�&�7�â.�0���4_n�4�:FpI��:�f@b���m�f{�@_��n�S��x�G��V�*�S��,�uF��l�HO��G�ݍv]w�|��R��YA�B��zr8�	��{� /,��v�m���ON�f�z�_9�j���%�Z���r�2tu��%��"�<XCx��� ��EJ_j$�@�3�x��Zk<�S�.n�Ek.��^�+��&%�qOz����
���6E��i;�J|�%��X]!�̦X�,>Oy��m�*�|S����ZSY(N_I��B����e����\��t� {jU��@0�T�u;���s���(��`�6o�k�Q7,;��F��.�@>()~G��R��2�!1��`&���$IH9:�%0,�������l�����C������,����e�gx*"<?򯏟G��~,��X��0� ǐ&�
���E��"�蟑���	�	�"����b���S$l����V7�i�s� ��WLAov����7�������	����o��������lg�2kY��߻&�.�r�}��a�6�
�ˮ�4��>��W%�z��C,�#X��2�i2y�_��rnHG���.���!��zI ŕK{'���;���?��%��ܫ7���V�7I����%����&ߊO �$@��'��T��8*�v���λ�
�� �c���T[��%�q���P����(wV��J,�۝��ݼ�ќ����";L��d�Oh�&-����纭e�C'�4E���Ա�b�H�6f{�P�V2L9yWPb4P?�|iV�0�W(��7h8͍t%ʨ=w�}��tm>��8��UZЇY$����8�n/�W�J٫5�+7�L��ε}>#>��K2H�>����N
g��S�%�h�� ~z��k7�bpq���k �>m-͈m��=�kѫw43�ga;[��������P���o#&�,�2���M>	Cbq)����<�bS�M�U�:��Ej�.ga� �R�ɢ q�w '�O�.p,�'�^2���TD	g�^I��b���=!�
9JdL����N��9ҊЋ�l\�bJ�1��L��k�S�����\���j�C���
�r��X�2*Q��N�q~P�W%��ٲ�:A�c��K;q�ڼ�a�;俴����|�]~�c����}M��H�0���xk��iR��I{�ٌ�?�yg��o	�o��X��רa���<SR�+Ez��R���G��*�LzK��M*M �Lڕi�je�F�sU�ȑ	f��E��
~�5�A0�]�����}�=���_�\#��â�1%������O3���&��=D��?5���
ԣ9���5~H�)[���x>�:�4�vwK@�X! �	(����;��^�Zx�I��GB��\�����ϴ�g�2��'���,�}V�!���e�m������1/Y�	g���E�r�K�0v��@Pv��
����h�7+�i�Z
L��r{�`l�J^�Gd ��܌��]�<l�/�d�|yz&N�L������*���5Ii��v�M�?�{4|�ZS�t��U�	m�cU��((����v�72�:���0��'QTM��v�6�H_�-XC�ӥ%^�&�3��p�E�:�Tk�_
��R>B����ee�pы	]څ�ԲG	�[������~�A�'k	���tu�L��!�>�GNOP�S���R�(�v^�)�<�B�Ei�v��T�W�'7!V����5��܈��\�$V��\��ۅz%	Y�v�H��Р�t�:2���ql�/ust0s'�0�ɢ�}�;�� �us =~�����ZnOD�zz�BU��hs�VA�w�&�����.ϵMp<�����
��n���ya���͐#K.;��/Vc3�9���q0�e�ܸ��Ӎ �� "�k�J
K���͠��Z')}���7��'Y���pb'�b��-��n��{#o<�������:R�m��c��;��{�A]\/�Jj��g3Dp�����^�\d5-u1{Y�+���D������g,��8�v3
A�Ku�Oo�6���C$��>�^h��!}?�z�[x#Ϥ���g�9�[�%��G/�\��ta�cv݄2�\s(hR~��E���OM��z��+
v�04���\མH��$x�o�xn%vv@�9����Is3��(�R�i�Icqd�S��@mCԾ@RsEx�ҟ~��:�ω8[k;ħG�;11Hx+�$O���|�_��Mt�-����h���Y���L?�!xs��SD�� ��F�i�i����ŻP�S�V^��)zL6���Rd�n�c��[�.�PLE��t�{��n`���d��]�9eƤIr�V����K��2���a}&NY���?�W��W$���J�|�+� c���+L�_�I1��p?�R���6&O��+\�|�{�K�Վ�wr,֊�a���a�����A�u�W�[[؊tJ�F���/?2WV����O$)e��)�]��X��FW�+��
�f�N��7Ư��i���&;j?g�>%�4��U֏\�b?�h4s�t��k�C�&�aQ�w�P1������"ؤ�<8�}�x�jxi�_�����>�J��Y
�>��i�D?4��Tņ��J�)r�iw�P�a��|x��	m�F��1lhp�'D��f/��>�V���`?�~L�n���ܴ@� �����bA�������-p��iF'�Ǿ&�e;�G䄞����e��.*N1��ʻ� �Ed�%/縞 >h2ڱleLAy1�+J�K�i�fSOO�H!�#@���v���ݽHn��~�%&��j@]��@�x���zb� 2����&Wp����Z���V�^�?B��9�$�(-ƃ�Z��x��}�3��ث��4ɰ��T�Y�7�%�(M]-����8X^�P*<ҝ"b��EqϹ�G��{<�5�|�B��|��T�(��t�<v�a�L~��<��k5�hY���V^��6E��}���3�,v�HN�j�p���|�� ɭ�y&Z:�-L�����-#�4o.2���{��m@�8�!�ʹ�8�fls{����uͳn5H}6��X_�`���<������g%a-�������5-9�������;�T,n���]ٔ����S0��<���XO�gͣ��k�o��x�s����D&����h�IK��iZ6�������ڂ��Af������`.�m�h{����ՃR�gH\{�.f�]'���Lg ׌\�\��������h�:ђ`%)���Ԏ�ߢ�	������=Q�(��F�~PQ ݦ�^u���a�L�F���K�����\=r�V�kfyN([���sխ�~X�$E�32éLW 
Z���8���I[ p��LiKKn�+�87�Y��Ӌ���y����u ���W�ʥ(��2�6-%۰��(�H�&�
�U9���|��&�Y��F��No��H�职ٗ���-�P�I�pgH��G�4�D(	Yw���\ g�	�/1H>MB���H�3�v��	�ϥW��Y�~M�$P�B�߆u<�aXg�t8�,�>��B��m� ���e.�MT�?,Z% jS�\�n��6�"��u2_�
Iz��Y𓸰#�P�f���Hoz�l��;��k\�6]c��WY{���z���g����=����B�2�Xa�����rC�Ȇ��q^� ܃�*�d����| ����aH�H+��3o�{r�#�w�8����?9�1�l7�-N�p!�[�U�����뺁�5��br�VKŽG�u��?�$z4��h�yn �y$���#�|�P�����,��4%�D�?��נ8v��;�O��AS���m������󚑸�4��mǔb�gGhZ=�(���"�hK�k�k���l��v�R~�(G4��>`���� s�����5�zQ��7UL�p"�`��%I��ǯ��Z�����|zթ)��f`�z1{�	>��(��MJJN�];^P�}pK� ���"���Ş����l��+Yd2�o�F��I��2���~ՠ6fb�$!�z��#�>@旁X��[�|�G��T�� E
*���tj�{}����t�e��%��8 +�9{g$��ڸZ�!}��N%���[Xg�f镄(�"�}�j7e�5δ=�t�,��P�d�ğ�H1�|c�G�U{D�Ś��Thx�zd̖���[�����
ۂ&vC�TU&�fF/=�.�5���k1�_�����E*�~��2�x�����3 ��V�" 4�.�x
t��nBB�F�ǯ�Y|�6/�~J�9�;�^P�,7[��N��2����[��ցN��� �|B���8BV�~�����.���ȴHHKM��N�nΧ��w��Ӻ̃]J
���pYBn(�"��b|*�*�M��r�T�؋��e�zP=JH��;�-�?r �����m�1b.y���^a�_-��0��$jT�$�N�^�ղX��tG������D���&����̥=��� ����k݃����M����ȿY)�}Q!β�*An:IK0�����E���o]�]�x]Q@ͣd,��D���KH,H(��G�*��c��O�z�׍	?��?�����hA�Eh�| v6��鴈��3$��uM���Num��l��'o�t�����/�rr�G{e-V����g�E񬓲��P����8	����B�A{W������b2w���[`l�N~��#�����P�-�\����������D+��0�JL���WA��G�Zk��@�/����&R�E��Ln�
@$j`bk�vi$���-����^������_�U��K)-9��`lF��F�G�O��~��)��1tp�CG��+�v��G���]Gu�O�����K~�������N!d�����
��3�j�c���OI�+����Q~)U}#Ȩ��</Dkv�KHh5}GE);�j܎����P��'�����9�'�a	��/
�;F�r$zߪ��'c/�tG)�T�x�e�R�VQ��W)m�딧%8�'~m93�S$���H9xU$yV��3�S��[~,�1��N�0�ǊR1g/���7�Z,���#���q	I��J�d��Jύ���wHJ�]����k�X�Ȃ=z`�"^L�&Q)N�|����(�z+��JҖ6dĦ��gA|I�e�# �L���έ�=P����Q�v��Zg����Aݴ��^P�h�cQ�Nr��������ߐ"(�T�(���C��g	�ocT.��3�Gg�mF��*&`�e�������V��Jv���������\FӦ%�UxS�X�W��ĸx7�|�����Va��=|GL�1����q˕2m v���p���B�%	�Y%�� �GŅ������l�3DK�""�&6: 9a�B�'/\����ߝ�*�*-��u]0z�Wt�3���fX�{��.�s��dRu�-jwh��$���'0������H����q&����I�+���5�	�g�=�*�PK)q[|U~§K$��PZ������t��
΂1��tr�>�qm�F��cy�9�펿�A古t����vs9 �6�&��̓�8�,�ա�x�RQ�P���}[�Q�޶���e\����2��$ǥl2hÒ���Wu�:��	 �^&����{w |8�^��&,��4�\���û�o�n#	Y���b�e^~���K�l��՗���ӮGى63D�I���~ź3�Gno��!�� Ҿ�{��HY�?���芭uy|Zs��+!w�����]��]�8+�t�4W����4mx�VZui
c[�;���
�m����K��p��zX�I\�'�̔�zŃof:?5uA/��C<�Br���6P~]��՞��֯4+���P.�Cb �أ����_�*Pc�	"�I��~G���:p@����,}� I��g�<��$J��;#CbqU��,��W'��_�.�x^����=r��n|�7v�g�0���GLb��%����;���=��U3�D+��Z�6a;%R�'ؽb�*���/fc-�i���DC?V\ď��6X��r�y�r���[M�����9��R��*��Ŀ-6t���I�܇)U�t��귻6��=��K�ԗ��X:c�D<}w�]$�H�	��|����v�:%<�Q8��X�/U�;�e�##��D�^~Ȓ��0Z.���n���>��OV�>�-欃'RVRe0�s���k�>)ה�q��r�u��&��u��U��8/j�����f�C��D�z��oSW<{�|�Ń�t��_8V�����j+��_�S(�`������ɻ���|g�����)[Tb2��ωz�Q�+ģ�ah��L�ņ���E�0��b5�hG��c�u�{���=��ݑ�mJR��8�aO��C�9�~s�Y���XP�ҏWf�ֵ'�b�.F��>��\W���j����蜁=�Bm��\���@������!甚����愄�!&���BP�q�݄��M}������wQ�{qQI���>��Y�V�h�l/�z��@��lKM���n�3*Z6��E�U6zș��ӓ����!4���I �}�ȓ�������s?ߩ��6zz5��6��pa[�e�Ϟ8̃b"��ZgSTN���X��d(����ە�6��7gl'|��E)�Q�n>��%�E��īM	��)u!�Ǯ��Ym����3������I�$�#���(�s�j�*��k@�j��\"��V%�)��p]-���ph�8���tw9����@��/�Dr�8mK"�WP�R��Ջ�'z(���x7o�����_�-�'��@�4�y�>8M�![�<&����{�e��nG�F�^�wZ9�:�+��
���P��'�~�v�{��i~�Z3^�NM)fN��8�$WI��XY!�w�Lkյ�)GR���ҶI�T�كr�_�����2��Q$��~;�3~R�o��ɱ���tv�i����Vdۧ�������Zxq.���_�Y�6uf_�2~��	���,��ᢣ��n�((��L���F)qU-�O�e#��A���X5p ��L�<;�d9�\k�|n��k� /��NY��b��:��v�«m�������t�L�04���.2-'a{<L�|I
ծ�3deO���PK������]��/���y�`���B���%P��Y��0i�+ �d:��鯤�ħ���$c����g5�Z��f� !�nEK�S�*�)�g{yPw�����j��������x�bG7���K�FE?�=��ǐ5�RQ����-sIOŴ�O� E�IR�Y��&��NR��ڮ˭�ԗa��ũ�4��~HI�~��o�u���a���i��A��	��%�F������H��vEZ�C���(v��ӊ_,�槛`f)¶4u�C��(W�%PP�� �@J�{?f^;��D;p��	�Сn�l~Ԛ� ��S�nQEU����0�i"v����c���FOty�p1��(�v5Z 3h���S�;m�t����������o"\��=����>[�9?�(����\	$h�iy���E^X�O�0�-�wUњ�%�eo\�nupZVW��F��A��9D2��Z哮��Ycܱe:Lۯ�Q��]�^$�i��s�~�����+@,+`�HZG���H�܏�$�!C������T�o{�s��l
�i��>�AF��D�#�Qon��d�GQ�ʵ9�:+�u�P�M�_�$X(V$=�Z��=Vs.�*�n ����W�x�{
dh�����#k�����*єI�w&h%��H~fe
�!�|{D����'p"?��T���W�p_#&G�;����-�p�4h%OaO�����+��Jq��kԼ���VF1�NJ�1�b�}jG�ZUKzJ��F�;CP�����(�Ub�Lg�0B��u����c�i�^5@"���L9�'���U��)�mw�BTJ�rH!	�7�lA����X���!%c�����-s!�SF��|���֟[����=q�Uw����μ��\�M��{X������.��رm.%әr`��n��<�,�?Vr+�H�rql� ���f�R�ͱ �%-����8�7�{t�J=�1�Y�Wb�3�!L�������h���ܣ]��=�2/�ϣ����Oj�<�	W���Ee�1^xѰ��P=}�B�ך�4�J�����~�[�b c	�ˣ�(kV���TP}�cu�s^~]h��پJ�zr� ��\s_Z�ӣ�'�l�r�]ba��7}ԣ���Onx8��]|��dQ��ߙ�C�J��N$�܌��T搆{9��:q����q��1Z_!'�~s#���$�H:��t��V��y�ۈ�n�=���Ν�,&�\� 8)��%�[}�����N��bB��S�d�~�]&��s�{u��~�O���.J1�7��R�[��=�l�[�Ѓ�	� ��˷V��2��<oཱ�B�H{� ����c�Z�ʯ��uO��՟����=#�	0L��Y/��g��M�J���\��ma3�2����@����XSz�4۳yޘ:�p�ȸ弎�Ȣ���Ϫ�|�͟������A�C�<&�`F��[��������[��>o��s�*��@���ph�&����ex.�%AV��D5?���ox�:�O0�B#�'�'�*�;���u�&�2�$�8�9/n�lE��jY�R���6�H��BI��:�u�����	c=��Pg��ݩ\�QK��j�_�(n�CCsN��R�7.e�2e�k�S�;"� ��Fz�w�J���������or���okQ�~�h�$d�g�}��9��+ʘ>)xa�'��1�%5c)"����Wd�xU[��85͂�/79f�1R:�ز�0݅��G\�1�T����|P��3��jԉQ[9d�f����v��q}������♷[ώ����Bn: Q1b$����Bo'��
7�>#6�9��M�`�qgb�p�����rPt��dw��zz�����8����S��5�ȴ��]Ճo�y��V��*S�A��]�����n�H����!��6ӷO*G"/��j�.F��:����sVY�`(���{¢�!d���HS��\�P�)Y�$x���hx.u�P�"_u9 U6{�.���|������0�;8�T�a���wإ: ��y�����_(����@1�;��,jQR
����~G|��k��Cb�4��xK�4���2t�e�uD�s"[�;NǗ��M0T(=َu�(Z_�G|�����1����`i�#:K�H|�e��}�v�l5�i�����d�D��YsW
	&GH%�ƃ��!ԺAa�g�xh��)�?���A�1�CE[,�c�5���?�^��y���!�P��Qx�Z�F�e!wXtV^+ɡ]���TTXK�ݑ-Q���P:������'#�<���I/z��~A��8��M��$��8�y�*&�����#�����(Y�Av�t"�6&�B���Gþt/�Z�hL�'���Ez��T���Z��ՃNMc��8�2(֞�L"�[�C� V�ɠ��yt��t/�#��|�7��o����m�E��ӕ}pG����7�9�3XZ��g����}��I�;.
�XeL��l���	�bFM>z��bu1&�Av,\�$����䒟h�p���P}��ubxQk�������z�Fɸ�E}�M�s���]VY���[e>�=&�7'L=;��	t�M�2�҈��ԇ4��[��L��L���nbu��`[ ���D���O�e��݇����X�xB�f����~��Ѻ�#���qZX�'�X�C�F}q�:/�_k��+�����ٓ'�rB���f���{�-03=���c��e:����yD�4%T�EYbFt� ��:eB�-+����4PI&t��p^*�,��]�=UV�Mr�X�ݸ'T��9�z�
V�%�7�&��v���`y���"��f��A�_�SmQ97���zKrR��2��i՘���e-I���c�IN�� ��Һ�*)2h�'P��������䯱.ry���G���L�n�C[>�����'ӑ )8����D7�� ���.,AÙKq�{��D2���$<���43\B,�R"��o���CoH6���'R�hʚT�w����㫰qٖ&�yv9-f	l[�"��2���_�y%;U�K���W��S���$��j�R��'���=ؾ�Au	z��H��w����2@�T���6�5&��D����?����^�B��PCc~[�M16�}/��W�l��iM�^����[��G���Q�����Zh����<�z��Ń.7,�k���ᢹ�RN�_Y��^L0�dL�s�
+�-R~¼��_}��f�߾�In���ޥΞ^CH��×_Z�NM��n>�E��Q�3���|ǩ��?I�&�o=�����
6��FQJ��k��+k]�H���5\z��U��W��ǭ��Ĥ�Uwc��н���S1�w U�<Ě�'�S��rzb0ұ���E��憧�E�o�pj!� "��-3;Y�������T��U�����6>�a+��>�xbD�2���������J@��`��iBgk�.�cL��̈́�7J�V�|��7r%K���|��=3�]
:{�)r$Ψ��l�JÛ����Y�(_�N�	��Jq5��Kg���:T��r��Gtә�/bT�-+�����>�<(Pސ�� I`��C"�_������s��l2[�օF��s��$�w#�J�󏈧�>WB���3�T&�=�_�CR���Q�*:>C�lK��s���s��k5九��ֶ�V�^��U�a��5�W[�y���Ol)��'�{:�f�8����6�
((tC�@�u4�`��L�5��iy�`L �A�2�.w��|
�MH��yI �:�K�ӑV�9�4BnY���%}��`UW���&�H�Q>�k}5�W�ᢛ��Pn�0/��V�_.AGL���EZ'��r�㍿�ͯ��
S�^�Tn�1m�ڸ�Qu'���{��y�
o����3���!���E��s(�BO��ߣUjОZ��+�)���'��^��[��^8)$�],=�X�������x 7m��U�UO��G$2#�Lȷ^S]�_�H�����B�̍���1�1;YOǻ]j���s��6�m�6�VX>��_ܼq��"M52z,2��sF)=�gsp�����> yLP�S���L1MCr���s5�n3�n��a|�
̄��~?�Jz@�t8}}X�1��q��ջ>Eጦ�$�Y�~����~�E�?GXE�Ľ�y#�p��C��-h�Q�U~+[��(��q��r3xQFp|�b�m~�A����14p���~3��>X~'Ҩ�u)I�|u7��u�D��"E.��h����B�g�Fք�0^!�����T�����?������Fd�jc�PhLu��@���T�47�.�7���)�\}�'#���^m���	))�~�$�ڇ������*�z�\�.�o.��*ѥX�T�� �f~��B�{٦�ų6e�<Q�M�\�ܕ�Y�pE*�s�n�=S�:V����ʇX{x�CsAv�f7b4�ǟ�8Ɵr�B�E�2��T9u$���OV{�9�T�"S������	����Pv�Q5i�Ep�d����Q�LU�Q��#�0�F�lT~�mfG.������_�n��ݞ�J?A�#�0�%M�����%�kO�]8D���Q�t����E��}[�LTC�M��A)È3G��j�3Yz
M��u�5BH�[E`���C��=�\?I��V6�h}�c���Q@􈫚�.��Z�i��-Y���ٖɴ�O�B�X�gi�kjY7�u�=�ø_!�Z�hD簋�%�6`���gF��8�\��8��Z�g�0�)���]?	�B�`��W/�NWo�tj�rB�Q�!��n�K�r���Bb�wjg�&��Y������Y�id�,��k�܃$�u�=z^�p��ģ�^�Q�Ŭ=�2콹�7ƅtV�-��ꧬ,2l���)I�:�:if����<�Y-=�a�a���]q�*&Ak�ja������h�L�;w:�3ii�'��?mY��	P
���7�{�k�(��Е3~½؛%0���8lGI����7�˔"��񖹬��F�N�9�{�O4��Ⱦ���(=� 7���/�F�w���	��<��C������eiE���2.�E�O������d�M����8�3e� 55�TJ�TsS�:��}y�:#�����Hզ��J�'���ƪC�������8��O��T���O V�7��!gf��KJL ;����&y�7���
�� �/����q:�����7+K�1�6�E U� B16,[�,�fk��<8�MB��R���H�^z2��v�ژ��#���(ыOV�>ٞ锠B��ޔs�~�l,��NY	�},������t멿H	�����b���$*B��&@�$��X8}Ц�ǭ�W�n,���	e�eJ�@��O ��U���!�l�{�mx]^h��M$M�������{��^x��ҧ�;�Yܷ>E�|��>CqhBׅnAwgw,�����)"���S ���Lj�3	ؐY�p���1���J!�n@&���[�\U֛�Y��/��0[��Eg�{Ah����4�!Gk��1x.�� ���4;U�/}�Zy#����m��4��K�_�+%�q B������z�7jo����~��Wp��UT��%���*�J�(\R0Y�y�Ahk�oyV1��|�b����;�n8�
t���u�	�L�]�`�e*�5y�)N6�/�o7��~*��n�a�"#퓿��#�sb&�eٲw?�k�a��0aV�DD�\s�:fH��c���=���û�4�U��>8�~��O��\��Y�� ��|#��Z��,L�>�^�M�z�B	��+:�X{����n�H"`�����"��g��9�̳�o7���>щ�s*1\j9�B����w�)�-��=��J��-I�CcT璖��Z�̀WW!���3ښ	��#�]�����F���	3dp�9��G7g��ZC�l{M���v3/��zӛ55e�tCÙ�v��cO�yB��c(�9[x��b�T�o~w�r����6��܆'������r�_�C\� �?�[|�M���b��d�+�xʷ�?E��E�56�(�]�8-�Ck��������l$	zW[0�I�!���ߌ8��`xcN��2�2_fb# �l��XClY�����۫���UY��0~:�(�M�z~%�h��5�o*�w���%�֌�?G��.)S�B<[L���g�(�n�X�9��je@A�{n�Qz��I�c	G���g�AW�c���oM<�6�i��*W|Or�"��.�?�[��d���C�Y�r��T=��T�4Lc,������ooX���%�[����I*E ����3m�%z~y"�k��;Gt��	�k����߱��i[��y�5�Ys͏?JWNcὐ���0�'�IOܔ����{�}����q���;�0C<d��5+I�Ϋ�4QJ�*�啡��@m��U�X68���̒ք�q���o�]���s̞��5P}���:xrʢѼ�w��OG����� j+���jP��� #���^�x����Q%%B��Q�Qΐ��(�ȵN��gՃ#f�@`�D�V�#��q��_cr�����_DA�SQ�U����|@�'K��������>�R.�0�ߵ8���eR嵜h��6=�����R�Ehۢj�U�2M�.!wn��:�Krj;�Ϋ���Ձ�b�/��Cʾ�K%��j_[V쾐��I:�hj����5�����/���׸ں��q +�H�$^����_o�Qu^���imc�&�r�z�<y�c���O�~�\'BKh[��Q&��&GM�ef�-�U^��1����i�pץNӶ*]����v(}�>����V����\���<>-?�$O�c3��@?���Ș����U�?���6�m݄(;��Y��}���E��`��L�έ�P!��,o��r�c�JXI�ST���&��.mR{��鹪���Vrc�^P��S��J��"�յP�0w���wc�=���zW)���VE���5�Y�;�vT]���~��mfB�ݏ����_�UR���
�+KQ� #�u�-��EtQ��y�W��&b��'��eW9��%Ս8Y��+W�ŊZ\�����L���o34؜��tҹI��7���Ǔ r����Ц���rpN��vy:n�H�XD�M"���=+w��,DP��mS�K�Ԕ�nŶ�_���%��Gl.N�c�����h�6��sj��`'�^��y��3�V&#��P4��'�E?A,��:81!7a��ɟ�����ĳ�ﯾ�:��)���12���M�:J�}K�Ln<����S��_���F��X��1��E��X �'�k���w}D<�T�	T��k��|3k&tW8Б��,Ȇ��A7��Ӟ�}�f\���i�L��AYu�))o�����1��]�O����	w�7��}�i���]`au�VY��<���(cyde�����am��>�	���b�Bn+ܲ�81��Wlo��X^u_�f.�r?������K|�jvX�� �z��!�yJ9�@L�*�4��c�ra��l�]�',��x��	@Ѧ6&L�1l�K��6�.r�X���7^�Iٵ|Ew��5Uv�l3��~�O�ETD�ra" ��(fJ�B�O�NTR��k�15�����!���s��4���?��OcVR�h��,Khu�f�ۨ�H�'���S�p�]���u�`�U��]2-�/��j&D1�ٔ;7���?x.� 1�Y䒅"��:2��r���e.[����^����(k��.�ɟ^ ��$���>D��O���)q����C��CvT�g73�>Z>�@��^�-:R��rb�����ݛ�2�=���r$ѧ���[��N����u�F��N) ���0�.������g�_}��@�7�����()��%�w?d�T@~�I|�/ڭr%r��� ����DC���ËmQ�MM���c��Bn���{y��x��&4�N)S��bt5C/Q�=�L��
�v5����G���m�k���~�o���,�R�c�~���p����?=r�_�2��)(`�0]o<�d6�B�$�U;�J��X�4��Ή�o�����()8;���@,]_"A	�LE�ja\��{A{��-��@��2��|�f�/�{zB������l�͗x��ڄ	��L�W�`~>�X���)��˻q �}� �Ԝyi87�����6�;^�����__Ӛ�uƉ��>	y�ʠ2�X�G��91�U�e�X_�1"��q�{'o��`��|"m�.�3���R�y�Th��SZ�ƌ�'�X��#ҢE#��S�ᖙ�K���o#o��5�͝E@$$$�Ȉ&��I��}�'u+e��=�IW���t��5��O����nA�r���}4��V����b �=gcO܋�Z~ g�8k��A�R�5`r�3�u�6���ī�ٽփ���J)hw����$�5���w�6U��
�}�p8����y'3�tK�!8M���@$+���œ�c7�6�j��i�b�h���M�xE�����D�-�50"Ϫ�d��NL {�B=C@d*��n-���ՆD纎�<��㐾1;@ ��ƽ�|��طao������{fku�L�~��px�Y)���ds�����+�C����&xEB��Y�� �>�S����@ ��RO'O��~�)�d�k�`���&)c���������:H�~�aھ=2'�?�#�ɹ��f�����{>��������K���2�cOT�����B��gB��!G���;_�`�̂s�������cbE��k	~�钸"�B��$6�p�\1�c.�}�������l�u�}��X�X��mL�!�
8�x�vI�Ӭ��3_�%��Ӂ��b@i�$�o����ɣ�6�,�u[-���R���f�2
����9C��6�4%Nu��t��kң��L��w�b����M ��@���%����ЭX�Usl<D��@[�Ā��y0.�����4d:�g3�}Ң�U��!��vk;7r��F� ���0���q�#ܞ�5m��,Ӭȫ:���A��#d�9ts�|埇��{��?m�tB���FAQ�^ع!֝zkNB]�\c����Ȅ+� /�Et(�lş���-�G�1J���,��$�j�a	vƲ�D�>^��;/�3,���ל8����`Q���H �|f�,����q�v�\��K�K? ł�p����F'�����'b�H���NY.�ܛ��~�ڇ� .��`�IDڌ0�C����D&�{=,
�e])�?+F���?��@3ȡ[��̹�PEK-8���2�s8��8HQQ�L��^4$@a(�.�1?������:��u��-qo/u�F>�>���o���J��֋+�Q0��ءGj�zaI׮F0�cre�ݚ}���2���.�bV��0Ws�W@�l]ɉ�L����PC�'����0٣�t>Ai�@$�F��C���.Iߥ�sg��x���I�*,�c��;���W2�~��ߺ���b#V�3޶j�����n�+�>���7��L��ŌP���O�0b�U��u3�u���(�
�-���  �;����/ٙ���$����C�	hF0�1�=�"c/�Zn7Q��p�o�7?�v6s�Z'���v O�x~����GN4�E�I��ř���e��f�p�5���b��e�H�ֻ��qS��9�W=f]���� �H �߫wxD�+N �.�x�n�_QuW=���ގ�h
nV��Pؓd��R�����ڃN5�����ƺ� ��O6��G��=d�)����ԉ�'<�UJL�1��\n<���j�v ۇ����|}��eK�xh@h�E_�>�Z��䋠�҉��,~C�/-z�Z2�򧨮�%[��?�@�8���W:33�����2Y�.�Ֆ�oI&i�#:jR�>�=V�W�.��&�s�y���~#@[���/X�BS�|%�6�$�b�#�����Y�	���ޜ�P��ſAdMDD矨�v��G�4�k�,Q�~ƿL�@�g��P�}ːv��"���b�c�<�<}�{�6����G0�D*��mr ��Ո0݌o�mT��ZW�B�ƪ���O,F�dL۪K�p�=�Ӯ�(�?x�:�e_H���v"ŗ(�^��ypG����{�5�v�BĮ��/ZOmC=��`{�۬�&�����V��$�V���[�>�����-�x6��A�*��;A�@���;����۶��qȉd��K��E��^�L%�FN��f��%�v�(7�
�}�v���&?	�E<U6B}�|�<�x1�}���)�rY�}Ԗ&�Ba�|�����ٞ�	0��$�4o|�iq���������P��~�ٱ��e�[�Ж�y>n��M_�1Bt�������m}i��Y.5m��D�����CaüT��h]r#�T��Жk��d�^���!-$��(��K����<ɾC��r[f�6X>�UY!�{��\k�M����݈�KJ,�o�_���[�d'��B�mm^N�g"ugƾ*̼���B��y�3���/�GE��B_�ez�9R@C�Q.m�L^ʨ40)e1w�jw5'b��E��K�6�~;�� G!R�5̃�Lo�M�z-,XՒb&���Br��֐3� ��0w=���:�\Qnƣ����Xp�{PjG-"ǁ�.��Gw-(���}:�<��_K�z�"+���9gkڝ�����P�����9'^ێ�����Z��8�����5ԡ�@�	�^]�����C�O6���!Q��I-I��ᶺ�rD�&��Y�Oû�s�5������{�P����L��gNPϕo��w�.'�2�V�ΟqG?��d����5�Zx�7���0 mV���0<9=�����h~Z3'y��a��~���\�6[��O��Ug�	#d�zvw܈k)�ϯ�?�H�n�62T���#��:��G@C�g_`sZ�����g�R!�_e�M��r��Y����(����������g���7������l��G�aY�� j��pc���ƻ����&D��<�;���{CG� X���⛕�z_��V�C�=Bz�2�h�Ifc�X��
��풞�9�o�@�("��o�> ���G�c��`��C�4��]������>Cw���l�Gq�i�S�0����72�e��ԗ��}��{d�ʠ���U�
=���/�u㤄�s��2T>2�;�:q1 "c�a=��X��da6g���_d�a

3(k!H�"���������@r�u�.�iݷ��A�W��˙��5���`s ~�eC� �I��5r8�`��n�kP��� ��|�ể�s=*��M�A�-�3��կf�>kS�sy,Z����Z�9�M=�aI^f6�gZ��9����p��t^�џ.>Sh�b�~�����jWa��;gb�Y3����x��ry_�w��~�HUoU��d�$>���K%Tv��9�nXdTKj8��(ސ��o'��ɾ�ʳ�70���\l��G57��6��-��ӿ��t|��U�!bW�2���@'��n�Y����fX�iҿ�jZ�]t=n�����u��S6`;�f��9d�@cR�C�Q�������Ӆ�%x�g�o��C| d��ߖU�*/#��fAW����5����F	:��M-����1��f�K&�a&r=��A>Ѐ�1 ����
�_RE�7
�7�[�u��\_��B��̞-��(��`ӀܧhΖMj�T�P[۾ʢ�_p6���]��qU���-9�<'/(����f���'8�������.w�[ڌ��?o�oG��+�]գ �������HI�r�R�5ll��ڱ,g��8O��Ӿw�RN%¤`�����au�I��b�o��"��\���ƛ�#l��橰�9 8`�;��_q!�#��v�]^d�wd����V�Ƃ�����R���L���Pl5]j�����9Ӂ��D9��K�]@��T�:hfɖ�;��@���7u��"�7�lc�ZV�4ȼ���M�_EM�=�2 �]���2�=�&�y/�!~�ཁ�oъ���Vշ���'�):i���A\���'�'#�<��<CIA�Hڙ�\ɵ��:b�<��fW�b��4���B"vY��0\G;|�-f� �"�d0�Y�}� ����}�V>�ϑm)Zeێ����	�n
�6<R��پ�>p޻�g�&3��}�l�e����IT)´v�O`�M��H�_5�g"H
�ӥ�i+�e1�m^x>�L�H�W�\J�Q=�"�a]��?��B$$1d��suWYl�������ӖQ1����oٵ�A]63Bm���Wx�����'ٻ޲V+��3:X��^c?͊���DKL��dD�pIl��&h:U,���b)P��:�����*AցT�s�ϵ��q����0]��QT�x�2�@%y��mq<u�^o�#u�؛T�o�$�V3�e�:!g�S�c*!���q��h�ݓ�⦲Te�����:�2�w#���P[��p�uV�
���tT�0g�^^"��-]GSP9΁�����1)~�D�p�}����@c��^��sy�v�޼������T�Sk
���M��
�W$�fX�1:;,E�6��i�QB�������a��}jrT��O�U��ʢ���%�W!Y'��E�h�]�a{��RA��"����0C��T�1������U�Y=Lv!ԭ����e���#Ǝ�+j��4F�lr�M;��t.ܸ��Dҽ˩�\v[�:Q���&Ȃ��?�#1sk;�Iл0a�����������,t�M�]��0.�Ef0�<>a���@Dj�& �h�4DMB�̃j��[X���k{�^q/�X,sҗ�7K�ph_���Ķ�)�ٶ���q?8�Ǘƈ���s�'WȴG�{���\Q��4E&檤Bb��|dÖ���d@��p��F8�ꪟ�?-V��V�j���*�Sۛ��v���e��Z?Ix��s��v�%C�ir[�z������w;�lfL1�`�]{C<�˅~%I�Lt�J;�)K%�:�'o�s���w�Ũ����w�0����#�*��.�(���n��W�s{��L�I�ܮI� 2?�R,}%*g���e'`�iݓT-~@��u+��s��\<��6i9k3ڑ� �G����i7��KL�Lw��葊��U�|�}�^�+<��A4�)Mas10'��H"��[��X��G/>G��xt�Bh�L�n:�	����GZ��\���YB����mgF� �a+f槊働V���)�J�<㝊�TC��;��Jp��867)Y�+*�z��F]ܩ��R?���"͹��rz���������ur9(jф�@�N�W��hܼ�	��<�D)oN��I��F�U�KA]/C�\��r�
П�4o�g9�z|�-��H;}C�t����;�m�(ۄ&��VLgV�y�{ ���^�ֵ�&G�{����נ�u��UkӀ6�����ޅ�� �^{��S����-SW&�҆S�>vfp�5�HC5ZM-��OM�蝯��[�8��.C��B+hф����j�=í�����"�k�e�2j��+o|����y·ǮEF��ܦ]9���g>�h�-tE@�U��fͥ��͉fm:g�c�Ȇ��&��9�}�.����Ύ�ܺ$�_1�0q���ɢ0�ik�{�_��q�ذ9�E���A�谸��0;{��{��l}0;&���Oi�_�+Rt�s�F���6�#��"������V��]�����6Aoߘ �uw�G�e�����)IT�^_�Jr#^T����	�V�o#�/P$`��#ؙF���yc���$�w��P�3�Pbt���t���M]��YW�P1�,fGW6�r盂#��&y/�^�C�r!�{n-m��7�x9��)�p���d��B׸i�j�Q�R�2�d�a��� ק�d]ΎwPW�`�練�0�1:[u�։�3��4l�O�
�:�+����������ޱȵ汝)	�@����f$�c�M��R���̗�۔D�W�C���J:���.t�J01�t �͜Y����[�A �'e�k,�Pϛ*h�w��ө�����B{㆏P{�pzkJ��7�@w�k r~%͈ �h`,�(��vd�!R����p�ڸ�^�0�]�.���:d�Hj����H*9��͙s:��d�r�(�D�pn�f���V���7���{PM*�����8�d8C/�[W�[�Q�
����]ދmj�QxcH��PEA�ly�"2X��U%V��ס� ۚj�\�]�4��)��:0x��4=���������w	��
�yq)��'��9Yp P�,�Şm!`G�B���4.���&2N҃����C��"c_T=ʯp���Ԭ�p�۔?(
T���uY~�	I�``�0���������i���ww|0 Y����G�MP�;`ah����>�"ف��8�ڗ�.���K�Ia �~��Ǣٛ ;y��ū���8��.���*!cZ�v;�M�I����4��D�s��T�|��ϼ\ �
]e?4�B��H ��''lu�${z�CӸC9Z$zYک).�b��5��Z�5ذ�5����F�BYM���.�{�cƕԕ�"pb��LQ�f���V���f�۬�F�&xF�e)�:��1!���[�����E-�J���m���/�ٗ]ut��PE�ݏ�E{�+"ƾ���8z/���p{2�^#��x@���7@�V,>�<�>ѹۣ�e��-g��Í�����R��s*��s�~p�c�
|��dM�%X�dWdub�t��\�ME��`�}zT��]�Y��8����������� 7�r�e��ٗm,� �j;s@ΪD�4'>z�z��iQq6��3�9�厛}
[��$Mm��#M�!��k��Qcg�U�Zu�iݾ_űI*�i?wd@
rK�I�;�����c���D�j{��wueH)Js�oZ�	�� \){0@���1=vI_׍H����2� z��Ds&8��e=�;�|�SR��-D��O�?������SQz>���3��K��?�=Ł%� �dL�P�D�`}@���-A�=�,�BuD�o��xu��.���%�l�8���k�ln�n��U������"�|=?o.�H�� >����eN�x�ӯ��?�3[z}ˠ��GU�K��?��矧��*��pd�_�b���[h���m��������L��nS��c��B"�A����[�5���^�cՁ��fR1V�ҿ�+(���%;��s�/��.�\�>�ʔ�� �V�$7��)���3W�C��$9�v�_�H�ߗ P��������<@[�?�(�E���6(�W�q�g+h�3^m��{ҡ��}-��� lޕjk+t��9��%��[D<<��>�.Ԩ�e��Lk}U����� ��I��/�^�Wγ�a���X-l���� Ͼg���:Wb�f�?B���؇`��u�v��%`p�6|��шbs�#��������,�Z���T[a�Q�no�	x��O�V(�Î���dA�r���	��14��>@�bۥ�s֎~Js9��h��h�K��[r�Z�dv��ؐ�{���F�ڸ�	�ģ$Ti�k�1���[�]������$�3�pc#�nl^?�[�\�+t!�o<"ю�>���;":�w<��=��#�jLz��Y,�c`���0�C�����2�F�Q���Ad����vt�����Ȩ^�Y��j�z��r@����$7�}�E��M:�������y)���;���M�%�?�鏅��ƽ������6����������`�׏:���k���������w�S~��}�/~�Nz���ɀ�}��!m�I��t`��}z���=�{�ɰM^�>9��ct'U����,ok7L�m �HI�GS��hkNÝ��t�;��oz�&F���3il o�8T�_�U��y���N9\h���ɒEZ��/�D�������޳Q����lU�j�&�I��3$@��PV&����B3V�~����#�lLԌ
,��BۓS��z>��q��}�9�W��jr�`ǻ�rҬ�=��p��g�����r�ՠ#-2�a����\��mfz�y1���z	�O�\����'RM+�i�)��a��C��x4�A�$�%�����XO+O�,���LΕ|�(��ly:�B�(A���+ξha�6b����(�P��Ț=�<��ş�/(�-i^��Q�E�Խ�j��0/�u�=�+��n�u2�Ζ�Lb�L���h��Bɜ��VM���A�2^�'W�`�����s3��,�),:�d��m9�{���f4j�zuL۞�h���l��q�ȉF@��/���T�*�aE�RZ�j�҄p,�P��RC�>K�;>�R�sz�9�h�tM��c`�5��@���ͅi{�B�R��c��o3���g�-C���IO�J �2M���`��V4!>9ߥC�����ɨ)S��,�DJV%�=��N�6�[�D��k~�Ƅ\y��P���@D �MQ�.�Sfiek�!$�J<�V�flo��}���M�~m��2ٍ�`Yy�.���]�P���/%�erɚ�󍼙�ۼ����-�Iv�,��@2m$Mw�q@q��-%kb�KDn��y`��Ƹ7�Sў�O�8(�]�zO���x��/��!5Vit�-F�S`���1�� 3t�C��ٞ�Ph&E�j�)-y�[ouU���tlJA�[���4���Ge5�Fqؽ�M���@��-'C%XMݩ��I�lKj�* Oku� q�"M�o:��ɺ1���}e�E�5s*�Np�i����S��ސ�����de�N���Y���R���k �I_[`��%�/��S�B�WcG?�ĺ�<FSr�����������w#4w�v��zRBަ*��G���<KOP�ƺ�{+-�&^�K6�Ex��f���C<���H�(^�t[G\}B�P$��GB2&`�,oQ%s��C�#�N��	;�0�k,�&&���G��z���x�+!2��,�a|�i%�C��I"�6ku�x�������l#v*}o�:׶�Ě@�x�Ts�-��MPp�u}+G�(������ݽ��%}|i�Sv��6�YP�!����������[���na��ڞ�N�{{�D-;�*���:���W��ZU
R桳�,j.��䆟A���[&��3����Q��)|ck��5���,`ֵ���p��[���mfO�\�,A��-��cX\oV��+�� ��������R�%�-Vl�n�Jd�+�}r}^S�F_��7�-E{)�^�V'�bËd�U�n�aƻn�"J3mW��*'�<@��K�j����	8 �/�\)V&�7�&��6	��fI}�ɥ�-9��)� ���g�~ܭ{���U�( ꂭ$	�+s�G(��;�CBunT,�Ē�s>�߫h�(���$�j�-Gwx��oE3��蛢J���6tR���(jHy�-���̧�rGE��>'�[�l*�@���B,	ԶXl1�R�1��TV����f���,[l�7������qW������q͎���F�`P�oJ!G���jI�v*�q^�&�8v��Ŗ)b6�\�U���hoV�\�����-��0GÖ �8�T���F|���a���B��Qv��E6��_R"٤	qa�ٵ�f]�|���:)햡dʊF��־�����p��� z)t0��d��ӯDHDՠ$���v�U,@DE�>��K>���>��^_32�Vz �-K�r7v>�,k
;lF�V����:�#m�������j㔍�7j��߷)Ů�꬈ң�x�y�gcF�L�N��r/4 jib��}C�������j���b��w�� ��~�lq�����d>��n��˷j��t+kgg!c����!&���O���yxt�� ���!���؜ta`�=��h&i9.��A���9lli��q����`h3�#'�r�A鳙�����"T�䖨�(o�W�D ���!@����8��ї�.�S��y�c^J��J{�8��y�pd��X��q�9��c���E��Sى��֨)�����P���s�s�G}m��Ohm�{�ɳ�CͶӪ�5M����/���)�'��n�_����:O]�B���~�A�l�Ҡa�J���cO�NU&�7�^l뀳�%�S'�W5���==�z�f��Ӛ�p8�>d� N���p[ �� ]ʷ���@"��X��o�_��˓D�k~YWp�<������� 
Q��C�>
X�1��0a8���`==����-��} ��A�S�P���}��1FH�W
��g=�K��<s�m�@��	�R��X�6��tlk<����W��G�1UgO�7u'��F���y$J�MOݨ�9>I��an!7V��؞�z���[�L�DsK_��u��e@�M����.��s����_�.���^h��ͫ�����g`���#D�����\i6��e���+������~�xU_����X��r����}�ž�4�2m���^�w�2��K�w�墏�۶����4���q�����Q�Z��L��K�Us_� �u3��+�a��1��
)�~i�)D�S#���^�y�Q�=�3@Bx�bM�
�	�+��7]Fn�ŀk��v{����^E4kK��8���ح�$W	tY&&���Wf궿 ��}��6��R� e2»+C�"<��<����L�s����{F���EW~9�e.��������V����A�Xo!Ҋ�+��I�M;�I�_���{����RTu,�j�����p�L��7�In��9�\�U5Ω�,��m�sQ�A�3L>@���f��&D�;�!eΛ��:ש����vl��N'm+��(��ق�D�v4��!l7hfB���+[�7���O�*���x6�����Xm!3]��Fa��\F9 ;X���W=~^�	�b}�N�Zv?~� ���k��4��dE4	GK�}.��Hu��/���h�Lݴf��Bg�x�2i�%��쇓z� a�� �$�Mf]��l�UX�҈�n�%��InT���>]���Jq�i�o�*:�&e]D,����4;�А��O����~�s �Ix,D����f7����Хh��7�����93;�?���>�b�9�ga��g���J��v�ņ���:�6B�'�ϩ�W��R��|�8 ���*��!����B	��]9�X��gN�#�K8��U����J4���#'�M�FQ%E#n��R��.�Iw'���<V�6��w�0F�}����6��%Z�x�s��E�$�@�oq0scL'M�Zy�M) �f�$�C1�R*�I�Y/�(o��XL�;�w�(荋 �2���,�ΐMI!㡣jmhhz��R�h� �͛�(��L�����F�a?k9"_� 
e�H�%��K�g"���G�.�u2	k6G�%�B�@�M���@�$�ϊ%��6�bײy9�����CZ�O%����+����g��sW{S��TA�����^P�����E7��?3��G�)��d�e&zv� E�F��,��I�x�p�������.�*�ၵ/7E8��W���A��`g��$� Ԗ9<��/}��������p"����Y�P� _�4��IM޷�a��۠]����S�t�7G�:�Lچ�x:Ē&I���T~g�T�������(jE�2��re	%��+�@�LQ���a�J3�U��j�k�+�0���M9����Ô7(��>1#������u��e�s(�Y��"��	�D��Tg���r]���}�g�G���c%��Gf)�JD�i�"�~E�-�R�L[�w��k��M�{�6��/��Y�	���Qb�3����0���m�TiTl��X]S��U���N]1��A�e�B4���NC�?�W:=#�a�!1A�#��/�Σ�����A��Up�C8gxŔ��@s�Ӊ&�ͷ�4+�2O�e��_@(�%&b��EZ˳�!֑`o�5թ��4���r�yS'sô�w~w:���hk�qJ�P�XЧ*�bQ ��{TL��X6r���o� ���*��I{��!Rk�9���r�L�YM��!TMH���7*w����E�-�13������wȳxƀt�]���,ek,QZ�E��m� �ܪJo،�h[Z�}U&g��1	��
�JH�~Q���õ!����2�6%�N�E���J�i7��A%P��|p�1ٰi�c�����T�\<w�Ք�*;4�z�{5���2��f��g�ަ�#~L�W�L�AX��p�=�뵞jRr� '�܁��mm��^1b�ZF���{{��n��B�J}X��9��z�(Z�6��zZ�+�qa&<Z%�<o��x >�b5Y��n�c�FJ�ZS-owL���
�U{k*�J?k_	��	"s�I��o�����q�ĉ`h�l�
 L�[u~�+f�e�$�ٰ�0��G�/�Ǻ���Wf踭��~���Yϗ�8m�P�c����\aDD,�*U��0 ga�O�K05qut_�V�G���A���>����,�@/�5���t����}+-W��VP��l�eT=�.�6`��pm٣F�e@��cn���I�OQ���j����T��~A�5����"�$�0J�KQk�}%��B��A� ���;�5e�^d%L�R��7���m"'K:X�)6���rm���H�a[�d�|���g[���0�-rY֡
"���tm;�vy��/���s'��J}�\9�� ��z�8���r k�'��K8��ܨ�	��n�5*K��b��=�"#v�-��[A|gx5	9SHO<��X_���l�����'���"h�6�PQw	ۅI~fp��J%��}��L�}���U�z?��!����)�8>�7�kѾeC�L���a?&'��I����w��iyx'\�1o'��P�Z!^�@��jC�LÞL��Z��;����?��4Q�yw���V�u��ػ��eIH��/F��s��	��|�r0��d(ʞ�I��e����F<*�nx�m�`K_tx7A���)�T�����mi�ak?R�ܰv�zkƺ����5K�l5J�:
L,���Sny�a��}�P�wZH��|ɲ6�Y�Z$�K�G�A���#��3�(���Hs���P4���X��r9
����% }�9ŉLNY��u�����|��x�uC��R�]�Bj��I�Pw�ȋZ�hz!L��6Ed�Zۢ�p�E��> ��$L΃/������09v_��]ބƵ3�L|��V�F��RM8A�5d+-���ܲ�x���S��/���X;eP��Y�� Go<9�W�H�8�PV+��������4�nc)Y<��C@���T��1��ʅ�\l���I^�ym&Xn2�P�_��xi���6��!YF�O)�����c��@�&O��^تr�yV�}�`��hv:+�D{�W�N�n�^vT���&���u?r��OZ� lɥ{I�˵�� �AOl����o]�D8 �����Pk��X��\����U���_;�eF�8:u�9ƹ�������S����P��$���{<�ڝ��_^�W�b�5	WEw�=Sd�5�t��c���T-\�s�O؏R���PwZu����2]M[t2QCհ�������o����QI�TW͞Vf��ǞT�dW�?�I�O�BF@��@��]�Y�Ӑ'��م3`��wП��}�N�+d��g� ���څ;@�ÆHΫ�˰�ccx���p|f1.�"�Vdή\��\b�6:�vvQ��[͋]lkIƾ��Q���2�Un]���V�͑���"a�h,��!�V�3��Ȳ]q�iE�8=�u����א�� ���+<�͔���a��DW�Si�	*�fj�����#.7$�vVuV�k5���[�'۾ ?�n(A��e\h�B�Ū�:�*�;�x,���p+���)G>cd+�u=G���:Q+��a���b�܄a:b���B؜��lѼЯ��8�m��(e�80o���R�=*����.O�or���P�S�`T�I��9r�=d�1�BoM,ҐI���6�(�v9a8����ϥז1���z�iq��>y���d��G�,���(�Yz�u#��f*�l·�3��nW�����R߯MJ�spG?���{�����5Ye�����[kehG(Ʒ_�7���' �vs�N��,�2�-����~b�7;آ��'���8�@���LA�d��v��?>��Sк�,�t�F��^�#���X���y�e`�\s)��CmdSP������[��j`9q�L�*���B���ͨ�jx�Q�;kR��&��-X��	�Zs��p�BuUMEh#��[����t�ɉ���u΁~v3"ʆ���H��2
�ɓ��}��O��ոx�Цp��"A�r�X���^��~)R5����m�$�W�d��� AQ�zg�l���)�Q���>E��;�' �f]���5�{PY��5ţ^��Icl�ϨD���?D�f��^E9~C6��Vؖqo$�e��R��e�����
<�{��%��h�V�y��R��U�!6BƲ�]	���-Q+�l�T�ۑ�3�'3�n��>2�m��4P�b0 �裋��������K�Eu{VϑLA�n#mL��yA����1�g�M�u���"�#�ro\����l��vqs�d=���"��,@�Վ�G�h�Iy^»��ν8�B)��K�M7�8럶�::��x�X���fs��L��]�x�4������l��R,��.9�[� Nb<��Ճ��~�������F�:��U��~k����U2N��m���
@�{Ι�Xv�9=�6?P$���o��"a۹��Z,����u�7����j���j��j{Q�uz�ElV7������x5�%�S
t�B<8��:�<h�V��@ֺ]'1��%`�?{��U`�P@��RN;8�X ��Ƅ4 ���d?�c�a�9�=*�}��bbcpF�(������Or`I�K�r��>K�Z$~S�6-"؎;D�f��<���;��Ъ�$п�Woç`�C�k]l�	��-L��~ނx�)F�,������~����T�"C����Ԟ!�m���A���� :jSQhcn�ɒPN� ���Z�M ��C%�!��P��c���Zq������%���Z8�	e��0���ι��#���c]�#���~��S����Й�<���`�(�G�����W��{<q�##��v��7-8���o"�;s�&�e����]��WmpΪ���Z��{@{u�l���z�u��L���� �HHf#�퓎��+�(��wEOo�D&�H��y��B����͈�V!�g�Ыs�4�+���$�e��]���E���ƹϘ��O ��4DB�r����!��8цb,�^ϫ��4��HX�I�u��ޖ�+�Ь0�J��|�'�ԭ�VN�^1L�u��ѻo%z��=|�2��8�B�ا5��n�3`��oF�oF���v;y �"��P�i_�c��n�s��}�se�C�P��q��9Ѻ*��<�Zt7�����:��kG�3�qg8K1?�c���_�I��[���P��l�e����]ē&�O��_L�7߆�/�O�i�x/M��]g
5f��_��f��R+w�_������5�I	���g}Tn`0-�d�6)\B�XB�`��NX���(2�*?�A9v�� 8=j�)^�}��v !u�>�f�sl�9Zt6r�-b����1��$�^����)��{�z�e{�oiX�� O``N���������;�}��jkAi8�V_����nRH�8`����6�T��2I�
{��l���|��ME�J����{��t��ёB����ڔ�rӏ�1X���RR�� ~;<k��X���D}Q)A)+C����A�s+��V��!�L�kXYAo�����D�?��|�=W�w�(K�5�4��26E����R@ƹ�!}�VʚBm��g�HO,��������X�u=�Yt@G�j���������2�� ���?~v���`Ŕ&�0ad6i�6��7;�>8~����yh�������E/z���܏�Ց�R#D@	P��'��v����ees���ݹ�x�(Q��î��d�0�C1.���"������9n�u?��$���s�X?�mq?Y;lu�_���Aw�ؽ���a��R=4뜸�9I��LE����N8��;lb��C�,W`{[0�T�n|У~@]�L�E��S6�H=����T4د�[N�:�iY*���:M'�s���,�ݻ�*���dg)������],y�e�0������J�*�@Z=_����'l7L�t�?���BS�o�A񛝩�����DN=�ʕ��"|	:��{z��/À��!~�k��>M`*��E��&��eP~�$��]��:LAwe`�:1�nP鴡tr��Q�=x���_X�:*�{	)�G���n�j�����\�OÜ�����-�� �N;3�ĭ�fV�`��_�^/�)�p%���1��I�w,y���,75SN�4�{d#&B��	d��|M|E����Ԟ(�D�2 ꥨt�k�������γ<�[�_�PJ%?g������o��&�$_4��F[�ݕ$���V5N�K�7�vm�I���%"6��'�	`'r����
����U½#K4� ŞG�M����ryCS��,��Ks�0ut1�X��z��+��V"{(�8B�3�a���j��
�Cc��<��D�ԓS�;���E�-�cMi�vu�;���'��	�iR@���]w�˺�N&�gD Rs3���Za�o��|(Ǐ���6��5B�;`_(��վ��a�A
�|� 8���l�2��7�KDNf�Wi��n���dׇ��^^�xy~9��%s<��9�Dh7t��Q�I�K��z����r	�/��w+�hum�S[24��B0d�W�2$k
�� �<[��8�չ=ܖm�TދI���39_���(��T�.=)�"0a���X�Ud�:,�1���QO�`��PI��2M����s�s�2f�V�V��@�"��<�<���[%����y9*��I)k"��5u;f@�#l"�����N�e6>�&����q���]қ�4[�r��0���㑷��wL�E[�uS8�:b5xQ�ك���u��u�q�B�V<7۸ kvc�?6Y�d�~]�=tG��^̟S@:��A�>0@ct��G��/�È���wk4>T$��%��˭����H�u�u�}6�[p
\��7Tբv��Ν:��D�/�6�)��D�VS��jpО����p��X�&|�H��tr���Hְ� @j�8�!m��ݲm��u������� ��WD�"��p��Yc����Rԟ�~�Ϭ�r9Q.YH�����0b����=�w��E��H�;$��x�� ���e�|�����
��6sQ��c�7�
���[tN�7b��9�'6�A�D�C���d.���B�\ӭxv���mN��j�B|���؏�k�.2�!��x��z�q�ʃ��m&��	]¨��=Y7�j`�7>�۞6��v\��I���7�K�Dxc�%=�R{�acK�|�"�S"�紗��%6D����,M/��s-��s��\9N��Ҷ��ȸ�
�i*�<��� ��)+�åGo���B��rDc�y��	�;�Ty�_ޛ�ib�b����[�V��ѧ{\�Q�#^-�ԃ�T�p�bm��`>�7��Ml�E[���lw��:ْw�w�g�� ` $|l).���4l���W�ꡎ�Ҿ�,Aȁ(��-F�.:�(V@,�C�E���{j;�����(&�3D�8բX(��T|'�W�7�*��ɻ3�t�"�U�a�mh��z����pW6�l ���IO�˕3s�����v�:���	)�Q��*��9b�:�����턃_��C��XA�ْQ|��~)ylp␞6њP��w��Bvn����$�h�xpi�Ƭr�j���K������\�1��ԓ�+|5����8��}�d?=I�|/�$�X�4^����@a-���k��!3��+ue�!�#��0�u��;�Z}�͆�$��-×B ��W�Ηr�Y�=MІ��oW�9<��}�+v��$i��2�sE�agF$�d��?Z$]���(M��B�&3��-�>-�������Hxٚ��?�r�U�P#O�J���ea	�`Z�;��n��������^u�/�ë(�ʐ�	��I.v~ؐ�(����ϩ}�\DQ��>c f%��> �[���L<su�[�}~��ԑ����������EXLB@	G�:��}�I�if ű�N!�X,�%ye�C�-�tLL�,��Ԭ���,YlS���d�Mg4�[Wq���c��qUs���ss��n�S!ΰ~�����?�����5� ���U	�2jd0 {�d,yWB6��Z���_����y|�N��q�Q�����0����)�(�Gr�v����w�RI�2��E�X4��ע�)a\@�`]�a�DE%\L(0��nh�顝�o����f�p"AZ�9uB3�-%��g���9N`<�ҏ@xc���q�
�l4�k&NO�k��T��E��+��n�ܙ�S�����b�
����ynԗL����(|�i$a���Ia	����}� �>/����8����Snf���ѡ�LH�t$�d�^.p���hx�f�5˿����V=35���������r��v�w��"���sc�,g*M\�F�w��N�d���2��[�4I��t� g N7"��#�D�DkS�8�'؇��URYN��o�&�]�y�W� d�lm-��ø�3�G(6C��`�n�\�ӗJ��,�9"��I���qp��]#�D;�*c���<J��Րú�v�,��ێΆ���p�:�d�����q1I��s>�X�}���\Z�b����J�Z>�C���h��vceUJ���5�<-�.r��pyB��	ܪ�������/�%*�!�IԊ��A�V=������|���@����3#��K+v8�I��<Ȅ�w�v��eW�NS�K�̩�Hh����$�w@li�[���j�,�w7�²`�WDYy.D�5�z��o�Q5�;���פ%�ph#)�<I\Lh����VG�K���Sh�_�M�x�1�����o�1J �ĉ�C� ���K{^��y��y�lP��6���Rg�K:P!�����@���K�3�4_,���/��|p�'���y�s��o07S"��5:�>a�h��XqI�Q���ƒ�L@�-%tC�:��߽Q������(VgX��k��B�e|D[s�,�ԏ��'8ς��nh�hb=��(����k�5C���	�����C8o�*> ������8���.���m�\o8��*N����VH��e��o�y+�LPb���ѻ��l��@�i��ɥ�C����>�=�D��R_�����I��`�N�
��w{��.�A��*"�����Y$,cB��9�B��t��L���]��pC)�r��[C��9sP���&VQƑ^���	c��^ �p��`�k�p:�WB���E�M��ޫ΋KR�M9�s5��crU6��D����pv�gb
�<i\z�}��J�m����miןH����|���>�;Nu�bʒ��W�*��PZ`�ҒE8Y�P��m��E�F:���g�H��#}=j1J�D�^�=#䖷��KM�т5�qU|������=��� �<�r����s�"���#�{�*|0R�)U jy��N�\�n�($�"f�7�Ȩ+0r��{�k�J$�[4�=�ł#��� tہ�;
tSa%_�*��u��7��>�A��s�����o��(|�i�T
x�� $\|'�Kgǲ����Z��|���4�Ez`B��R�k�]�-�md��3{�K~���	�;����w]���N/�g�
�c�!�D���Vc�;���:WJQ�TL�u����B���ѹ�p�1<�f�<��z2ow.�K-����>�� �\^q��FX>n��n%��S��"�#l��:�Y�F-�)|s�*�Bb��_�a7!п�?�#^Q� SOپVj�Z�Pa53y:���ϑy������}�F��>Թ{�|\��ؙ�BWn�9�@��;��xCh�7쥲x���*������)�M���aڌ0ȴ���H���2S���骏��y�>����.�8�v7�X	Pͱd`޼�a��O9�kF�c��&M\����[�}��N�>D����B���_�ȸ�~�]�h�,A^�ik5���3���F���J��tm���,ObW�1w?�vn1�䚠��3�Xz�.u6	�'{��G��k�p�xC�F��X�hL@����眍����h���h�I�M{�,9P>̳``��Tz�a��|C	
jG�"���ij�H ����K��fQ"[������ԑ�m�N@����M���`~��8@�[)k��d#�tN��%�"H��%�3~���H���m wv"Nr���&:��Or
�������#A�~�Gl���%���b��
P;��
)��y�j�l�/�Y�J\��_�I�������b|���$��u�� d�Rt���M-A	�]�O�G�t6ͳ2m��W;����88z�k�R�K�P+��i����s:�%�h��W�J�8V]tv�5wjg��5�z?#��~��5:�
j��eOY]*E�}<A|��|�m�\h���_9�����j��j�@��ۋ����	\�yta����f�)˭�02w�+~BA}���.��я�p��qs�趾�bQ��nMTHhܠy��h�}FWq@E���-'G��,ʑ�ԙ����n+��3-�F�e,���J	��k����6������u�C�f����j����-"z��	��W�Y���1I�km}������^�WS��~�T=��|9p�o� ܬ`A>S��c�_�F�_gnd�ѝ��Ga�>�{ʄ�%�Dfvz��龾ҍ����ɫc@ɋr��Ks��]��ՠ��p�\8|�l!$�n^�\W��:=��4�1(+��������c���NP�K+�'G&��E=
Y�hX뛐�פֿ����0�\�0G�UV뙘3����k7�m�x�o���G��ōXs����Υ�M��sZ\�[���r�i���H�r��T��i�N/�e��ꁽ����.1GnW����u��!������T��ǚ���l\�O1�`�Ƥ��p�4�.���ubO��]5�\�m�D�`�Vv�]�$޳!
�6�W2��G#y���c�:/���2��Q���Ůt���Q9�6���T]}��u>C��Z*�\6Hm���y���c��*ly'����O��%9~�N&ɕU����
���wߝ�����j�Ē��C��)��޴��E��еV��Ď�w����Wn��`#dEHv��.��� g�'�����E5�p��o�gV?��eB��ú�A�<Sg�s�H���y�ڠ+P�F=9��}�ASԦ�Mb��C�E�\+DL��!��J(�: D��p�K��
��Kc���$�b+�5��J��QN���½~=�P�/�!�.ݞ �ӼAe�*d���F^EmEq�����k�3�N~_�%�K�U��j�m`%]QG�%�%#�b<�Ι��Q�N�/��Y�1�M,v��\�y�i%Qᮌ'G�g�ԣ�e�f",�*����&th�)f�+�T%�QG`�7>q����Bڏ�H�MwHfU;V�]���C��l���F��1R��aC�
A��]��;������&@�X���;G�������2L�Y�E`�!7L-�r�>���� H֐}-�C�i��,w�i����&�(�Y �{]��Q��ģGl�(�ݧ:*'����:��	�m��W�
f��ߤ�� � �݌4��cb��v��)� �(��)k��;H�W.�a-��(>��D!P@a����^��K�EAͧ
�H�Z{���,��h�3� ����Rb-� ��1DPJ���i}�T<�����g��П �-�R��qS;܏�A�-N�)1��_`���K�R�j���;R�5?1)zS���oTAJ�h �`��2Լ�2v)�hf--9#>�g�,���`G�6���K{a��/$���ĿdY��{�����0�%�
s�eK
>Y�(�mc��:����^�ۚ��;�Sdm���_~O׋��і4O���F��ޭb��Ԃ�u�]�o��8�K�� �wD:U*�z�.����,-�I��s�W�5�?1�!�b	���D�
���MZٕ�Ph�$[�$%aef�(1�ti ���O��^h��)Jy<�R	=vN��o�f͜���p��KdLǵTm;vc˺nd'�ӎ�(w�����DF��dr����L����b*�����k��
����Dx�P�2SU m]."2{,]���S`l���@��}�$"��~=�H�#�?�m�c��=V"
6���)���D,6Lߝ�u��rE�Db�J�b �i��tx�D_��m��fD��f���)h�~����f0�/?f�7��_D�?�O�H���㖋D��*%JV@%���pJD�O�*���Z#��a�_�SE���L#�T�s��0���F<��X�� *�/�mO�P*U�j�����(
�,z���e���D?��I�@_��7'6�'`L�ݗ-����w݀A�.�T�G�@�G���َDhK>��Ȗ?�!k^Ov@?�.�������\Y�e��2S��s�?�@[%�cQ�oW����D�"�0���Zge�bk�H4��C�)"BiQ)J�
�����K��e� ��;�b��.���p�|/A3N�ڻ7۪��c��>6͜ݩ��wT��h���-� kK�pਸ਼ qۅ��/,���3�@3sB�i�J�����d��xᾎ�N�˃��9ܼ��E❿aXu��{R���G˂�{�l���,��āΑ�AL#/؊�FF��l�wR0*E?��.��lb���D���z�k�+*��<7ʛ㿾��A`�j1�fm�@�P�{2Ƹ������B�!Z��|�L��2T�@�8+��Ǜ^&��B%�pP���1:��B����x���� �*8U�@�����j�⑸~;�6�Z嬬�w}.R9A�J;X0�,� 갏�_˂n������nt�d�3�K!�>��|�}�Գ���T�~�m���Ll$���7bs���H��X�H#�cY�U%(���Ts��J�y�����e`�z�ox�����i�n_�S5�`L������Y\x�dϱ��&���:�^@�{�y�e���9&�(�P4�H6~"��#�˼�Jt�;����_hē�E]$�@Z�$c�z�$&���ݫ�@0T�0�C!)ΒJ��#f{Q$�o�F������Hd"�!����`
��Eċ�����Rޘ��#�l���\��������2K�1Oi�S���l�<݋	�5��{�*��呌��F��sO���j�����s�G�2��2�-��l�����kKˬ�ԭ��t3�����4���u!�H�����0�t� ��� �BXKPK��!�#Ć_2d��f��r�wX��Pu����^M���k~�4��k����T�)���ݟ�ɥ�"�z
p�g��a㢹'�0$�]ޖ`�)H[$����G�P���Զd=��|��oq������&Ӡ�-��6�'��0P����u������_(�Qd��m��H[+5^u	k	��R]�[���FJ�\��>cXr�{e�����]�5�Uv>ifm���4 l�m̶x���	��<��.�_<;e��q���dy��.� H�o���="ˣ�˩�;�u(/����8�[�U]��L'U��-�Kg2:�[�w�g�w��uB�E���;�$�f�J��[Q9�y�)ֹ���H��f��C4�S4
:�x�zܾH�=w3�t���S�m}׈i��ʪ����Z�����%�v8�<JK��v�X���Cs��9,P�&�7$�R�`�9E�dyTҦE4�ҩ�?�^�@3��)Q���V�"�1�2�e�!�T���G�Ш?����������d$4��}����d��q3h�wZ�ά_�~����"���[r]�X�cJ���"�\�s�M�lT�	Mȼ9���?"ܛ,�n�t�� � �ʟ C+�k��Z�n(+�R,x���nt�$���mo��s]d����W��:{4u�E���6����ڈKo�+p�����;51��_
��~Y(Z*��qm���'F#�s~5O��*ߺ�����Y��]]��ϱ��*�I���O�<M���F�����Uz�D��Q�.�ܑ���V�������������|��Gd�B���0����0_K���Ѯ���l�H8�x�]��w�l�^��K[� �h�E�� �>��)���F�^�% ��C�n}�"��ʓ,�{*�q<X#2�dn�"rX*@���g�X
:�S.(����7� G 봲i���5���ĩ�����f3��申�"�ѹ%�p	x��D_~��ˏeQ}�/[-��s��i�O}z]�}��E���p8=�����S"$@4
�}�& c����>R�r�wz���l��e�0}�Yb,cO��S*8g��[~s=����<)M�Ԫ�5�w��<��n��-���4bv]���g���~���J��w��b��&:��X%뽄q?Z7?Z���U/1����-�D��2a	���~y����]�!ȓsC~�0i�C4���[���fr�z=���	hC��������j�ܔ�I� �|�)�/	�S�.Ot���M+T�^�ri��Q�A
iBe
��L���w�A���)���"h�vL�D'�6a���3�6�S	*�d�`�\-'�"�̼ݥupzk܇|i��۵]��>��F�BYK|'ŝ����Pq-r��Wޑ��v�QK¸��d�Qv�m�i��(���x�q�6B���z��<�1�[��s�{ަ��ӂ�B���|M�-����R`�La��6i�~�}:%N�3��h��2À��~�Oa���G4�MP�8�{�Vl�9X��b\"�*?���˘���h�ǉ���h��'�&l4���Yy�4{�N4���<�C�241{�@��aBrz���x��<O�0s/�M���d���¨��H�ɢd��nm�H�j�]��?j�l�=��0��-��.���} �?��	��>a{NK]Rv#����FJ�ƕ,M�#m�;�+(�[�@#�!?�������uͳ�}ȧ��n��xK�}$N ��c��~��Ĳ���'1E��G�+��N��ݴ&�$�+�@�&����_���;\��C���F)��LX�5�a��.5V#�}�%F�xl��З�М��ǥ��qm���y�,�fͩ�{�z��o�)�w�8�
�
����:��5�%��Bl��x;��Zy?�u*�i5��9\D{0�R-�[\�h�
�ᕈRF\�9��ė=�W�UF�J��.k�o�Y�Wx!��68?7�%�[��t����s�9f�Z����m�?ݔ�`��ld.X���;F>F��	"�u����.�̾�6���Zr�P��+o8�#���o=�$�O_��������-U�p�}h�*�+���Q�8���+�Q�pQ��C�`�/Q��1���A�e��.n�m̽��2�=;�˅t�'^׊��H�O��*�Q+���n@LK�����FX���Ђ�4�5f��谑����lBSMZ�t	�}��µ�*O��;m\�t�֥̟D� �- ��y8�nm��=܍� �!������vx��K���Ylz��g4� ���P�0[ �Õ\=
&�U���^eΏ��� �V8CF���Ĝr�־ ����QiREgxݴ�mv�&�-j�X/h��y�Ӊ&�`�?�&�S3��X,M��j75vS�>ҫ��ss�U�����.�ɔ�y}��<4����2	�&�[PÇ@A�s\_��o���l,�
�QO��!���5:�{M� r,�G-�Nݸp��3�9��ڏ������;?c��C�i),�[vΰߪ�	�|�����\ M�2�}9/�2,�+���ZC�qK� e��3/q,c�M������H}ۃ2b�@���D&d�R��54�����.�X�6��P�r��͸��z�B#�N^�9rsZ��H�w�K�8x��-�FE��i�:ק_M�Q��B69<�V��g>��?�~�A�`m�f��T�W��M���48�������}8h�H����S��L���c�_"�BmdE��|����Q뗗M)�_����ZF^�^�'�gA�p�M�E�Yr�����GU�P}d����:�"�@r�'��:�����������C�������i�X�ѓ��BG��@���^9��7���f1�7
>N��0�1������ Z�Ξ:���~4[pi��'ű20�����?-��qvHT�)W%}.H�� ]!��L,9��5�WK�;\+Gl�>���h�w	��Q��7f"-�g�1SV���B���6;$ݠe��,����l��%!�,�I��^��$���B�7�2�J�\��L��Y�<�ZG`��HF�bq7�aa=��;)��v ��6�;\Ț!���W�&�F�̀&TK�5�����Cd�ݥ��Y���w�3~�d�ܚ��y����^��ʎ���ܪ���j[����ex0$�~�刞�O��Բ�����x��"�;Ww�W��{��&?�Xҳ|��rn#�?�z���./�������r'9�/�t$��d�(�^�&���m�P��2�~l�����`%� ���ǑB��|	���<kܶV����,�d!�=��tC:�zd�v6�n�pU۬dEr�B�N=�D����w��&�6b��U�ѡ5���Z��@[�@�,���Ԗ�
1�B�!!���P�������e�j~Pe�|�ˆ��L(��J���ךϧF{im�תa��p-*�JCO�����q�����T���?Q���Kg�X�E�Χ��(�9\����Z����_��3�ѽc�EFz����L]����$����S�"D4A���j�����(q��C�.q.������[;�}�G��[���-q�[��M;]�FX��p�t�c����5�H�c�-��6rκNXXO����_�߫#� �e��*�d���&̶~��M� ���n%+ߑ�L�T�z"�y'{�P��p08xR���nub������ "���O��R�lq�+`+���@I�t��~In_�|��{���_�Vج�Dj��	^�,����! �:2`��V�Q��Y���mNnW<�f��c�_9���ޝ�I��*�5�m��e^�*O!��ג����c�$hArj0����A?��V�C�fM9ŏX�Z��yE�{v�4���7��^�cZ�o������=|7B^�Fw5��q7�����v�`��Q�4������w���*.�qbJ:��,b��a��A� ^�uT�J�8�Z+�qF9�� � R;�M[�c�Ĳ2�:�#������@��q	�⢵�(�~���XN/�Fg��ǣj��ybm?=�dRՆ�hoߓ6�nx_�,��i��s��m��< �(��<�M��.a�k; �U8��!RCM���L@�e�!�:C��fa��C��	��S�����D
 �(�!J��,PŐQ{w,�l!/n2 �N)󆇦�Jwc���}�|�ә����V� �� ���lLQU;��Y�rc���%���&����������3�[/�k�A�!-����2a�qLI|X���$����i�w:S�(^8T�+y������򕌣���K���b���'b��� �՗&!�����*+����X�
R.��0�����n��Z��zo^r�����}�a	�?���_ճb�8C�,4��&�͍e�g�Q��&t(}jݗ3pU����Tm��<�j���O���tXr�����͠R��%܄�C���f��a�I��8wEbmΚc��U��N���d�s��xǻ���Zq����
����߽�$�ZqR� u-^wbS��n��������6�d4�L��ZM�Z�ݐ��I�͝Y�._�F�Pj�FxS$�����A�tVX|岤�g�������m�F�����|Ph[A�L* Sn���3g���\���+�,$������<p��C�W�yE��C`�L=wya�p�+{��Mi^�0���p�ЬX��LB
�� �̽yJ:��m�+�B�*+N�A*����z�
q�}#M��+O��-�(�1r�/&(�O�IJ�}�c ?°���sl����k�q|Y�9��Sbe��~��Cg�?����%  ��+O���
�f#�������A��ڣ仚xLf*1� ׁ�م����P�P���3��zb(A�'��nW�`��s��`��떹Z������V�B����Rt{���hNji{�@lZ�C�븲�B`3����e�����ہ
w�:�SO|�u��>�_@�tK�JN�HWEy�MO���a�׮�N�b.ijW��ꑝC�,qU�������:)&���pA�W���\�Y����o+���	)?3��G� x'o������?�X�Q�S"#�=�R/@<���B#A�����8�)�� �/.- ���S������)Y��ۭ>��GoE��Bt���ƹ��D{��$#�^���q(Q���w�����+�������]ve+/fb�uM����x��~Z�� �03�ЧI�Ψ��=W���&�삶�;�	 4:�R�\K: >3�6J�%rӰ�����#]-e�Y-h��Q+Da�`�t���<��K6s�w��ua�߉r|zo�$�^��#�Z�5P�g3�ꄂ�]l���Q��:�Z䢖%�~>�er�W����N����!b�/�4Vj�`�[,�:�F�>�P�vF�:��MrƩn��'|��(VH���ۗˬ�U�ؑ�r��Ȉ�����v2n���֨�M�� �J���(k�2�]�LTk�B���fKR�KN����k��#"�l�m�rtt�8V��>��A��͕*�w�νh���{�$Nn�V>�I����n��@u�e��OG��4�9����/15��ę)ݙ5ܯ�ِ̾B>3�M&.Ղ����l��&��$,W� {��8�w�8/ڄ�k�?	R`�{̙�蕬XMQIx8�5w��<q�@&(����D�C���?^c�p�" �p���:�|7��<�o�ɓN8�O�ӏ�^��UQ%�c�>�XSB}F^(t@���S�w���(�XU��Z����I�ĿD��KFB�ԫ�"��?���(tCuG�>F����ݸX���^&0b$�Q{>�1�R#�� *�v�ж�~����,"��J�]� ��\�H;�p]YJ�s��n-9�]����?�M�}���tb
%)乾cR�J]$U2�	^9mz��u�X��"�z�(}���D�5zT}�i$�����7��v��H.3R��CN�>$�嚴v��Ig�SP�)O���Q���k9�n;���C+�h�y��H�h��i�m��T���.M�*#(=f�ҧmV�V�Z��#*�2�#�ҥ���3�	>��/�V��k{�Z�ꠣ	]�r�)��JW�f���,�\��M "��-Ɠ�Sc���#�*��U�#�ח��A`D��؟(��R��=�Z����U����c��Ś�Xb��i�`ʻ�QI��f�9�=�q�{�c��Z����jP�i�y���]5_Ĉ���"��t8�k�z�mp���� "&��K��5� ���������P��N�������nP��Rg,3��~倻�[.����/+��k6���k�:�g/^�N�$ec�q���@�-�%�=�rBn�9�&Y�kS��OR�y��"dӁ�*��������,Lr�<i Q�����}��^�N�� &����g�ׂ���dh��#�m)=\k�5=�&b+]�>�"�R���p(���\Nj�Pz�[��^]��'��W.Xjp��4��D&/$}?���@Y[�*$k;ɱ{��1-�oy�]U;9���*
�����~�Rm�ޑ/W:"���gi��^�������s�%R��:6���ȑ r_�G��:�}jx����,K٫���X炙L�C��� &����^��FO���H6R�"�}wp�K{ʚ� �m��վ$ex��J�ԕq��w~Y�M/��vϚ��Ȁ��$+�=���qG�6+���@�
!�f�����5o�(y�2�'=y��w�i��#/��Y:�L-�g:�p��'Z�����/7B�O+^r���h�9`�����D�a'bt�`s3.�H�\4������V�U���$ F&"��F�Q�Ip�ā�����Ba�5�B�1�B��Q�v�åT/`ï^v ���,�tW����Ynu@x��G���b�2�PŰ3WHֶ�%�*#Y�X�wL��Z�����	��`ߩ��!'�fH���.M��`�M*�a���`*���J��h��:�S�7��*JV�bh�'~�Q�E�~E�0��Fކd�yҔ_;5�
]Z��Ě�p:U�=��������3x�7{w��p�b^�1|ͩy�b1#��)���;���5@�T��� ���E�f,!^"�9t���?x|���;m�U��n^�Y�E�i������b%y�$��Ռ�ts� ��J���Q�ޠ�l}Hɋ�W�n+������������Z�p�8����j��ý�j!{Hw�%���Z�"�M��KL�`�$Hxyi�VXw2a=����_o�	"]WdN�G4���mI���y���6	W�i���t8:	�<y�FT���e�| qQYn���U�����a���M*7B�6y��L�:�җ7�t�ɶ���i�7ȍ���!���f$:a�2r����|$\'5��_�5�L�����ж(F�]�w�Oˬ�#�ѯ9ލLg��\&~d[�jgZ�������Na՘�`~�k����G��m��������ߍ52��O�f׌�QσA�G'JS簅���к���w��`,Ҕ��&5	���W&he�{�C|}̈́׸(�� (�5���0�ag8����ʍ�!��0c�CR$1�20f Zb�߈|�K�a�̄	%��|=�"g�����;���aUM�'��j�~^�׹R�[ ň��K2�!�
���ٜm5]�Ε*��uW8���s���+V:KlP�V7{E)���4���M�Y����WP�>�-[�����&]�����<��AL�"��,b~�� ����_����iOmd���ַ$I�d<�}y�6���f�K�L���Q!ZT���%�i�f���%瓍����щv�GY7W��J�\�q5��-`,��xiZ&4������ʇOC�L��╨x�6�o�Ӟ_��NO6%�Q�0���Jn�NYZ2�I�Ĉ�ϖK��pu���+wQ��i��z�ϊh�l���[dC�5�[j	��v^�P���<����bG�ڹ �{X�3�s>���e��!C(�It��d8�jUؕ�0-��Ȟ�g+*�)�/�je!i� δKdƚ]'��oͳ�t�JR������{�s��p�R��5�=��u��Z��������7�܃R0�	Q�'M�ߡ�h'���
�L�Y�o�R��^ ����&o��iv����cW^��ӌ��ּ X���a��[�&8[�iJ�u��b��vsv�}�����|��;z:�Q���@����~[DD���֡��4���>�Z���Gt'쏑�Na��C���L)Z���;!b�?�eAޢ�,�@ (f���F8�"�Sǋ�l�-m�d�%H��Z���e$h`j�t��7\�r&�#�e���,� �b��� ����ƹ��Ŗ���,���wyZ����y����N̮x ���F.u�S�7�s� ,?������f���U>ү�?�� w��t�z����a��a9o�_�fE�]��=��F�&3|^?�c�'?[̄#�2v'�39.��ͽ�671xHd�v&��Ү�8-@��c�$M�H+75���Wl�9X��he_�^��+
|;��%�QۏFp�:�3�h�(���z��dˎI�S#<�n����Ɩ_)1�E�?���fb�k0%�俄���U1�X団c�m�(\�H4����eǚ�L4?!X]�NĘ"b_�U#�1�M&r���y�
��y��O*�ŏ�D16�G{y=��]���4��������#Fe��3��0�w�b�"ZOyA��ו��-�@�o͚�@��]��ǟ������6��o:��?��~>ڪ/��FFy*j
K�!܁��_�	@;�9�����$Yc�AH���K0co6=�u}��� 2��Q�������=P�.:qu�W�#Y�4���7�'sv���[V�	��m�ɓ$B�GR�߄�'!������������@	*���x1F���`�b�r�����X�@��]�-�a=iO+)J���5q���:�08v����l���U�X�=ո�]�naQ*�Urs�;d-oW$���~��U�U�e\�ҏn#�>K��<�w4��u�LXɢ��N��1��_�&��;;Ս^y���9��/�X�xR���=��	@Puˇ����t��23�?�h�ՙ���Z}��`ѕ��]x�,�<��|$�y�7��|t�jX��m��$ͧQ޶���%�d�N�������h����őw_ϖ�ࡤP�DE�/e̺� �P�9]��B\"Kg�Ns�sd�����T&��*a���o�����W9AO�C}㹾���Ya��N�n���҄�ȃU�UR����S����o��3sd�뒦��O���� >M* �����*�D���S�=Q,Q��k�C�߷� ��D�x�!�Z�"�㻊��y�.�Ĩ�g'4���l�g��4e��W_���a ���&��j�)���/�^�_F5�����F0�6�z�N�@���?y�}[��%<ۿ�փ�s�E�-�ҵEc���d ������s{E�u-��*٣��DZ��b�S���O��Y儑j7����n1]�a��!Q�X�}S@ѡ�6�ҧ�ˉ��S6�U �΍Ssĉʍ,>�e�\GzæA���4F��23��L�e��`d�4#g(Hԯ�����8��Q����*ef�-��p��*�J8�sv�C� (u��z�g?�;�1��w�M��#��ɳH,Q�R���龺O��Ul�,��Mu��!M~xE�KO<aʱ��LlO��VØ�FQz�7����^�>v�CN
%'����H~+��Ǔ�?��i���=�(���7�������x��hC��C��ҥ6N���v~���8��-$2���O�OT���+-{�Gs߅b���d5[[�����sY�Y�xM\}��=�:�~�ٯ3>(��6R=u:��x��%�J�SY��`�� 񥇗��ZŸ}��<ΘN�|�Ӽ��5�����ޮa՘����� ܏��gk�� ��o�X���n������3A�uzR�������K�Or�</��Z<Y���
?y
�9���<z�p�F��w5�QmЧ����.F��D��]k'�����smȶ����l���^�����ޠ;�U�< cy���W��b��FZ/�Xo��G��u!�\�y�	�3�`�Mj�]�r��B��v�EZ�!0-�{�)ݞд���� ?��[�P.��:����<��	���˓B�m�^C�#4z�m�3��ӥ�O�OG[�ݔ�ʺVZx~�����t���ebӇ�z��?�������M�*jc϶���X?gʬ41��a�@k��\S�g�uЉJ	U)X��y#�zՅ�����BG0&�����e}4���2�Ji\ lt"����F�&�5�T�f��ȑ�o����Q���Gi�
�E�lLMf�;�gK'A��o��̮G}w	�o��Q��@`4��q��B̵Т�r ��ML؞I�F��m[!̈́����/�3�R+r��2��N,�<�?��Ǌ/�t��Eb=ΐ{A��d�-��6����nU>�9a��2=��/�&��n6Z�Uyw�urF	�����Y�'��`��Pz���4B�9W��_7��<��in0�����)���F�}�MD�L�:�z�}_a�IU��";�ZAZ�	#�$�a-I���� ��፣Ϟ�
<��P����k�٫�ܰG�s�gv�U�)'j 3��vqS�z�-��^���2����I����Rn�q�,����E2�]NK<�+8�cj���k�M����'ҫ���_kW���x U�n	���!��S^��j�)����Ӌ �O4�~�M�'�с���i�P\7�ʆL/8rJ��LK�t0)���v^�h���M�i�"L(�:
!Sb�͒h�{�׍,�SU-�N_�b�G�8��J��j��,Є|X�d�N)��=�(y��d0�g�~v����t����MB?p
F u�@�/�Jm�`�1�:�	@FL�h�)��e��k�X��[�$f�'e�!�n#�P�SQp��Xw�m�sɺ��j�ٝoX�v��������K��0J;���v��p
�R�Hw8z�����z�m,Uu�Z�4�A��QZ��D*[��Z�fl6�eZ#�Q�w8WXN:��6rb!�#����TM��m�o���=��(�-c����a@=�Fū4�4R�[��/�ye\��ԓ/BU�F�8��^g��;�U��Vk͝�2�*�zhv�*@Z�`F�Ɋ�񒰍�K�&����K�igǋ���q�t�+���]�e�^�A{|�LRFV�
����X�E���@���M�VŜG?���<�(�6���D;��]��С3�Y4��1�n߸8( �Bc���r����[���A�C �GzS
�l)�\��+5CCl�{����α���(:����Z�|)Z �Y��!�c`���#a��r��ď�,T�o�z�h�v�S��Wp(ǥ�^A��Nwe��� e>��r������r|���|	�^o�9]� [U��[0w�&ܙ�~�' �eQ%� LeШŮ��6~�6��$>�}	�nµ}M����R�d6@Fݼ<7� <��X<�҃�J��Q���Tr�P�U�v[
�����_#�����)-�{b(;K�K�kn�u+#TT�m����+�\v�dA��¸��7� �]��M�-�nio|M��Ai@ޡ�����9��6ir8����Efj�R_\i��Q����&��H-w*�@���>9��A����XFkb�m��M.�i7~S�R������	C�3M�yY��k�S���:kq�{%4�8�v���#��6N��w9����)�:�c:�����V�v�E�<�0A<༆����P���琳�f�^_�0,��J��������P �	JB�E������Z6�IC�����EG��� &H� �~,�%�D
�PKA�M���սB�uP<����۵�`����l� J����M[h�(`��]��-��#�I��N�F3�aJ����wg��L�|>��!�D�>C75x*�c��2Z���+6�t.�E�+�3+�|����W.���x��V�?��_�QgM��9 x���rY�1K�%�P*�G�r�Vi��hOi+͗w���&GY�N֑>ѕ�Ɔ�fO�F��
�-�4���q�@B��Nm,0y�TFj?4�u���E�/���\���I'pu�ԍP�������H攉�|',|&aM�1����ZY����Y���W�M�˽�����V+2��no+�[�,=*���������5�=eҎ(��H�v �N� Ȼ�/k�����l228��~%>!>��P�y��g��ι�
�JS�o|ѐ��Y�Y�<����vU�P.�=��(_tW���
�F_+}e��+D�dR�EE� iX��f�)�l�`9���hNk�Q�%���5y��1j.&���Q67@�L���@�b���l/��dH(�&��:yV�����3H�P7RC$~	)T�՟�A�P	�86�5J�"AaU����D�+�VA���/^�wH�R�v�B�>��쩭��)�=Q���s�r
�_�-�9/&����=��&З���4kz轙�ڑ�9�����S[���ZeF�����v�3����tĂ�S��Wb;��ɐ��R";pgk�WDZ�X�W@*���=C,��&����N�[f����+U���0,c�n[uR��p����&@OW,��{շ�`�>K~�"�l����@ީ���S�Rlr�-��iɎ|(�k�G9UdO�e�8��F\�>o��B�	Q+�Gi��(%�|���-�����]��T�c���-��A��h@�K��C��W�����k")�lN#�@E�������~)���%�16I�}#]پ����m����5C���ٗ���h0ttO�`�?��~��E�i6j7l�O�.C���ž0�a;��J�&ԋ1��v]J0V��4�������p��J�f��L߱���G4[<u�|4Q���pzþ����p�g��(a��O-�B9����λo_�0	��%q�G����vR�h6�#��{'��#�e���;�Τ��&�ɥ$-C�'4��x��g7���n~g�`�1�hR ���k�Y	W)]�3����;k%������a�	[p;���׫Ci���ee{s7�k�8���Mٟ�p�d·6lA�^Ȗk���Z@f�p�.}86�����'�f�|��2���b�ّ���~oux�NY��>X���;�l�Q�`���*b��4U4a�S�m������"ꨄ��р)�Ó�t=�/���|��)N��]�폍9wFz%�c
A�<��r �"�� N�RklFJK�p鄦�u�r�?݊��`^�ƚB&g#��|�e1ٵ'|���Z@_z��}_/�!�J�IOi5�炲�=�5�lŨ9�[L�Ϋ���]���#s {�����q6�98�y*g�p�E�xzPuT����^�u�o�W�G�Fal��e��eB}ȹ��ケ��6�\[��1���Vz�3�F�q�Nf�����,��2�R�,)���>C*�)$�T�rly��r�1�Ѡ���^�4���|k�]k���ր:@�ɵ	��u�~}�{��p�r�w��cZ>:VC�;���ӵ��� *?�vKTM��-�/���.P�E�ڹ�5����;k�9y�b1���W�gN�D�f�d�d�a�������Y�Ymt<���R\��i��a��L�'���M䁙�K��[)KQ��@���� z�@��G�t�P_A���I��թ��1�����z�2�`2v�zgo�/7�'���Fo��pǇ��P��0�X{��^6M��4��Gr�E��_J<�fũ�3?*Y��E�p�
�� ��7Q��i���dP�������hN+�`�=���r}�����d�!��$ h(�u��`�b@/���ܴN��j�+��ߌ���B�9��Vq�~���X�=%��j�%:S�$<�E�y�=ČnI�c#s�@HH0Kr�yu]�D���}��U����Qn�Z`���	��+>��A�����h��>�� �L	��N����P?@q�0cֳ��[�ٶ��O(.tD��m�;��������z�����4��t8�:r�˫b7}9?ȱ�C�8��yy�?�&֣Q�W��������g�i�"oPJ�M~G�-���o0���d��s���������v�#���p'��I)�75���.���d�tT�T��j=oB�4��c��%w���p�l�2�Y�ܱOG�sr�pZ�UrM�����ۋH��d[SJ��#��i��=6�0%̇�q+��?�?�$.m�����f�{F�s���|?*G�9�ݏ��]�����	64F��5��q�&lp-n����@�6��	Ӝf�z��^�;��a}=d*�'�2��>���P�bД��~Bˏo��'��U1P�q�7��"w��Q��gpx���>�	�XC�9��B �eW+H���F[��(K��~l�/��e����H}��<ZY�-��+(�(8o��X5:�jK&��H���_l��Ɠ؈@�~ �9W�c~�6%w<c�5�"��ܚ������Ő�@�v�2�v��*g7���ILF܋p����F�& ��,��=YƯ�g�(�V��0�_#��(�(�ٻ��q� v��}��-�؝Ҳ���`Z�>���l�$�yK�;K,��9���9ps�#j�����dn���_�T����,=�v����ޢ[N��`���Y�ۏ�(�F��8u�Q�u��� �%@�	���E�d�#���|Rh��&:��3�ʈ����.��g�b	ݒ.c:I�o�|�ME���6�a�f3����/�����8��k��{sa&�k0SI�u��u���&�tX�ݐ����t6���+/q�F��xZ/�8��P����>�w[=�����-���J@x#�+�Y !)��N��S�N���,�
ܓN�\|�Rsg'�ٰ2F2?B��j����~}`�:� YK�XC?�mZ�z�oL������N_��O��ָ���8�8N�����?�hq���%Q�a6�e �����moc	�b,(�<-<R�=x�Gԭ��,4���~(�ץʪRM�5!���%���)�j�7!�*�]�AQ�[p�������qc������M�s�nנ��N}��.n�P��Kv�G[/+����U�~J}��L���Ky(Om�r��Į
�x�D>���@����N��g�y�D����t��bn�t�AP����bZ�~����5�`y�"�;��N���g)|�2*�
3/��{�c�W���
@��ח�t|}�(���i&�pGY���Ў�C��8L����|�����^��0k��}t���:��q] S4��`zork�`u��I>K|��Dɂ��8M�0�Fej�lc.�x���T�6�ې��WפI?.��*�N�T�v�)�Lr�>�#�%�Iz�W�r	5HL#�e���.���I��Pa�Im2t|��N���F�u�6�j�S�O�h�`�0F�&����$d�Z���;�����(�������{���A�p��^�	(F��WI�e줹�V[r�"�HJ�Z,Gn��v�m�R�	,*&��<���� Z����5���P�O#14]@�0(fj�p㍐{:c� �tcʮ�u�j���"a��Z�~/�W��{�C�����N�,�^���)�^�W�i��t�e]L����V=M�Ɖ�[b;������_��S���tY�/�rg����Yc-�("r<�V�5aK�q�N�H�/MVT�҂�f>���L�Z�{[5�R�ye�=(�s�y@Qf���1�Yi7�n��V��UlT2����le4큚	"4�r�]
wD���D��j��.Fu����f`Oh����	�Z���[���0������1M�$ÁY-<�ն�č�J����%|ᾨ�?`��x������q�),�*�b�%=�C$��H��GU@��1�x�AM��(?I*Y�v��S9]��`�(&����T�)F���PU�D�W�tq������������n�8�Z���+�ԁ���$�(+ք]�^	hm���d�36+S���B�ݾ`5�ܱ׏n�]�x�{4���>�nC�6�=�����?Ŝ| #IZѽt�9`&��L�ɰz�g�*&��P^
O-���e����w��K�Ȼ��A�;8fu���}���|-G��rM�ӄ��[���x6a���"�~��6����x&�#���[�H�D��U{�s�x�*Fi�N�z*��R��-*��e6-TЮ�Z��J���(�����A��-�(��#G )(�����ޏ���G�������)��u#�Y�n��(�2]�k�T�N�MZ�t�D>���!��g6\��\�!G��|�K�w���B`�|`�In#���X���:�}�;���4~ĸ�{o�M����V�o���%53%w�'j�nMW�	�2V�0n�����/"�+4����R7,��{�N��u���1;	۟�.A23�Vα!wf= ���-����H�#���[:{O��}�m�vO�6��p஀ X<4�CԄAg�F�<h|�����E��$��PO�4J�Cj�ЁL+��ڱ3o�v�<�o#f���t�IRx~�zh���	����e'[k�_ը-��lί�Z�@�j�EL��Flh%!	 &6}����P�%�WŁO�W�8$�6�s|>JL���>qqL�����kƯS6Vd�=�R�����Z��E3� �>e�����\�����ȧ��KPAd�T�t���M�5�ȸ�\%@b�wX���;��r��6Z�ݡ�:Rױ��>ԎN�Cv�7)��̋�m�+��DZ�(�>^����Z�� U���p�,��?��b2yDd���5,jP�R� !&����e��T��n��1r��>T��\3�I�"�Cke�>���rr�f*�c��O\^sQ=�#@$� �17�y@�9���))	�������嵭)c#��t��%� ѩ���.	^�X%˓;n�r���W�� �}���!��kr8%���ߐ)���!������D��+�yE�փ}\ˆ�g��N��x`��#�n��Vh�7�Ǔ��݈�h�Z����#ћLUR��U���������^��٢x�@Js��,��_M�������z�c�hE�ZX��sѿJ�B��Y8�ٸ�y�=A��c%�in�2�������f�̯- ��@�Pq�ݸ�9��4�r�=��K��vϛ�j'S��p��7{��w+��,���Ua@ĭ�,/�/�2'+�WI���gnn�lc7��XNI�8'��4��Ǣ��hd��ͅ�k���gk�����%[�a##B��kb�Z={G&T�Q�߉���t'.7��C�z�z@����P���j<�r��`���Gsf|�����f
�
�l�i�N�a�ZϋŗpNm�=��x��X�Pϛ-�L@nY9�d���r}�n�9�9�����%R#��A�	�^�?h����9�g�{i��%q
�e�?l����')'M�T�ʏ�s��̅�U�&1�F�ޖB7m4>�D~N�fOhw���=�ff�G�ܶlQP�?��P"������u��T������S��	"d:C���(A���g}�|�$�����w��Wr܄�
�}oH��������@�{�e��A�8��M�X�ȱ�����@sp5yې>�������k~6���M��}��aڳ�+�[�o�8ȷ=�n�d�`���ev��Jv��MN����ŘbB��c9�,��W0�R�]ꊤ��?�g��iZ�;��e��q�+4ؙs��Oz�k&���Fm�!]%����"�
6�F�C��
��ߚ�j�\Q���7�'9�G��|�[u�M����fj�N�Aʑ�5�J3Trk>�j�,��0�tƹ��l/���T&V����@��1����	1Ĝ�(G�Ľ�H�m�<�i��@y��d�o!v�-ȱuy4�v�pD����9X��	����y��B\R�Lo��L�������5��� g�񖾰�a �܅���{G��wD��$�Qd�6����r�͜N|k�
 ���n,Y��c���x����t�\;O�w� �cKm��T��"-?�U�l��}��L���u���5�w�n8��;��K��%��ش�K3�  �������%��_)�L��4n��@��ב���H5U���p�Q搿޻ �%����m�[�Ѡp]3Z�>I�%q�DE-�G��M�Z���}�w��+�!ty5�?�H��鯯�!��>�Y0�yQ
�����G�H���z��R-�/���KcB���=�Y��;C�5� ɥ"���br��>w�aX�'s ӽA��Q�:��j��T�ǜ�z���Gh�G�� ����}�7-k8���Lv���OM$��Q�� f��ls��T�fk��҇}����3TN�=������<�;�j`��$Z�nOC�>-�?D�>q��X��ĕ�ZJ��	�Kc�w�w|sK�]�|Deok�T���Si��$u�jt)��C�=v��m'��;٫�+s���-�Pf��7�H�O7��r������7sx�߼�b�R���l������h΃<�6&J&L>w�b��������m�V����t��5�L��M|)�ۺ}�Qo�˩����=�!~��!�ҭ���hf�ł�<~��>ߋi�V������bT&)�i%1j|�Ϩ����{Q&��b���Ci[�'b��s�W��nAB{X�y6��ۦ��R���e΂�9]���Q�K<v��#Dޖ�XА�G�?��������YHi�8>F�v��b8`�H�%�� ]C�O��,г���>9E��R)�w��9%%e�t�j�=5^�D%���v�M���=ڔW�*5��#��)���-��7D�3���0��z6�h���2�xMsW�*��'���v���_%���d#F��IАP�2ҿn�*-9���#�D��C'˶څÒN��Hn����M=$�QYy���P�h�&{a�)W]/If�L�OF�ۤ�;k9�_��{K��ڐ�V_CP��C����ߢ�Y w&�xFu���5��&L��	=-%a�Ǘ���E瀎B��oӺ���ˮy��ruYy*M�܀�`�!�β0)�=h��x�"H:����h�8o~�n71�mj_��	��78.�a�u������z�9�m	�k�&�h�{�w����]�C���[��f6�Rʨ�s��(%}��� �N�O��Op��օdI�c�mq�Ϫ��&����k&�YjAq� ���2�t� s����ڰO���$п['�N�ҰK�(l���j�t�d�c�J���Noޕ,��7G"FqXK�iC�|XS�t��]����;O��}ɲI�#P��]i_�.En�{j�B�'�ϵ�w�D�FSÔr�3͚�ֈ���'i	˘��N|=TÙĳ3�%��^����ױ��4_{b��ד)���ba�/(>�|�'@&.�x�^;0׷�}U�J�Xt��ƈ%��Lv՟�A� �|đ$�L��;��>"���f8ACޥ10�ߧT��4�zs�Qr+&��{���Y�ҼJ�� Y&d2�fi��S�Z �v}E���m���W�2JKN2/�F�363�3�C�1����Bx�����aս1���~\^�恭�LM�`c���!g�3��V����E)�؊64�q�f^8���M˛�hn���#h�����V������j��cdWA�p)*��X٠�aͷ��Yho���\2}��Y�f�Kү��=�0���3�6����8�.H3��Y��G1����>�w�`�����!`� /���K�:����������[��z�8lMT_�����=��)<���y<Kŉ���蓺}�@�F�jz����(�G}ڗZ�4���q�F:�y��L�Ҭ�v��ǁ7�u�[��o�����/#��67�ZK�%�m�Fqp����g�+��t��:	�N$~G��/h��~�R�%�;���W�z,)��VP�H�rG�p��ő$c���E�`ld=���n�N.R�l�������љ�Ch�y�Eu�~{�R�'��_���ը���� �{tA�a��QA����[��+�TA����M6�a/3V�֒��2�����>���tyh��e6�w�B���|%}�������m�F"<f�k���*t�ױ'v���LŠM�+����S��Od�D��S���Q�z��a`j�����d`8�w���`��<�Y4w ��Q�|����L��u��p�N�86�Aa$���ɚ3��\Fޗ�{}5:���m�9xkCq~p��� �j�q�8���uG��U7V����Rj��Z�<�E�wc����-�ʐi�n9�����?v[�?�`x�m�B�bZw�y�ENX���O�M�䥼���K����KGX��|�eߐ���ci�������r�Fjo�勓���h>�I�/{��I�iE��&��-���I���b�I3�	�5���	�`�� U�
�'��B�$�����x�N�y9N�4	�������ѹ:�$��W2B6�Y;��6iU{�Mz����P17��O_��[��j�4�{��J���'t��|<��f'X�#|J�, �~�,t�n�l�Q\a���g���6ƾl>:#7?�:�
�<]�Usd���}���痈���o@G����$`>�G��xBF���=�����I,�b�6)�2�<��Γ�D����:�ƌ�+�G=�����΢����N�������Xc���2+.�%"8�����Z]��Gg�a��a2P����0����ueV�Ma�%e2�T�{�(Y�uI �;��y;�vh���]��*L{��<1k�1J��aLg*l����HV�F��y^uk��6OE�vc�d����G�.�EϷ��!z��8^�W��ֲ!�A!����Xe�?�O��c(2h����Q�w��#,�փ���Z��d�$���_��#<��S,�1�&T�Q��P�BCD��/��b��Ϊ��{sX��h��u(��U��&Z�c��@�fP_��d�w<���ckj�y*�Nk1YJg��|��<ˠa��h�W#�T?b�����i���mKv>|&O��StV�]���1Ǵ������j~r�J�~�tR���S���h�f�&�^섕��?)������7/��0��1�8W����3E�9�����S6K�n�`���l��Rm�T3��c� ������g�n����������w䥫96t�&�Q&&2��Q�\f�l�MK-�f�%���hʘ�2B܌'�k�!X�l��=����a�R{~ZK`�KҸ]o�Ͱ��d8�j>v��,�N��*�-ϩ�oS�N�.O�Y%��S�y�H[����ۙ�u���ST�]e��������6���/��������(e�i�31�<Õ�~���bG!=��n,��l���2���<����S�EK� 3l�(,����z�N6��5	���r��]���~@h׵&�@�b��0�� �Zhsv��;�f`�����ei�=��|�.X�R�L	�D���0X����TF[Ŭ�g���x����;u�������<�H6�T����ɭ#�|b�2laF�����^�3/�τ?��zB^���P��1I<u�\u��������+~�pS��t�v�V�n�� �#V����c�Q��珽��VV\&5!^/���Ʊ��u���G��c\�%�OK�g�AL�xk�je
�wq3�
��GֳW�:�3x؂{�7U.k�^����7^@xA�=�MIl!�z��'?�1Ÿ����q�gJ!�_b�4d�f��*�|3l��Td�֌�&�i�3P���1_?
|��A��[L�p�`��͛օSХ�(&���Gk��.� �V�3��Vo�W=���$%�Q���`?�A̦妺��aNN�\���p,�k��QP����@�����Q=�Q�� ^u������z��v8��r�c�jK�8W7I'[0�!��L�G&��T^��nN��a#/	�� ���֋윰ɳ	�uc��)�WO\�M�����R�$��珀C!WpbZ'Zt%^��L�I�`o��&�I�-�H�)v�;zږ$\ �eR�p�����3�(��pUj0i�`2�M��u�z��k��3@�w�����`j]l�]v�� zyȤ>��mgDɉ����}d��{�{��F�Vo�����0�e�P*��)�R��������}�8B5���B�`D��m	��o37��}��%;�`�DL�h��Zf	�D��=��o��sۥ(�*���xEQWs`
3(X�����W��4�&m����=���g�N���N���9 �7��D�� �ZG����C�3�\��R� ����p�C�k�x�]ʤ7�mi1�JO��yg���Sw�6�`�#��DT����l����ݩP�j�<6͝F���i/�� �����Z)����.����C9�S��g'���y��AJQ�Q������`���Yk k!6��]��� ��&_�2�S���� ɷz���l{�6��P�lQM��@}�i�<:�-�8�e�!����?Wy���H�̔�8L����������EuA�
��y]e*��ٞ�?������^!�&��"�$�u�[�o���[#����}����Hm!���>�4�?��EY*R	S^�*޿ǻ�T��	���y��v�����؝�ӘY<��r�s�!����Yb<sWt�ʭ��D4��
��J��Kh�ݕ��U�ܩ�"e�����7��qR�X���BLd ���3΅�o�~.��G�z���_"�:D�(`0���CdY��N4�r���u��(�M��MSR�G�[�]��%�%��n������U��k��9�%����S<6D�Typ:�k
k�c�c3p�㵥���%����v�5���ǫ=�����n��<j8�N�i���`��u������`��"{P��T�6`u�I�����Ѡ[���{�Q��s��.Nt(J8Y�L�d��p\���h�"S���GɄb��)k�MReT���wj`~���X{C� o��A�%�b�G�\��3޼�<1oMy��@$L-�[4�ߍh����@�ЏQ�!����X 8�1�W;;�&���_Z����;�n_��=q��#�й��+�+)*���Jv)�e�ԭ*l6{���-M�K�/�^�6dݚf�y�YKFW��������p�2�P�k��|�"4v~�F���pY��}8����xV�l ���? B{�]��(D����ߖ�F���R�t鐥#����|��i?Jڸ׋HE0ʛ�h�V�n�U���e��Y���zJ5�<��@J�̮n�蜙��E�X��3�	�E53�76�<>��m�P���1�5s����B��X������tł�_ނ��RA��#+�sܔS�Q���-�Nv��Q�Q��:�!p�B)�z���?2�r����L�1I��qZ3�Һ��k+gq�h�j�~��p�ɕ�����	j������Ř���"�