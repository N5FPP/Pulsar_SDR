��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1h,�mwG�� ��q�
dh������n�5ӫ�2
�e?4�K�����ps�/)k޼��������a?SrL-j7%�"�1�z忄Q���͗��2��B; �/^R[����wd��\���
A3W���w2�;�uhs�SE�%�i�6H� �P�6��v挻g��Z2
�*UO?���d0�0B5(5��������\�AԻ�#�B�!������i�R��B�jm1��q�M,�6�
s�b�ւ�_���Ԥl'Âl�/Դr�v�6��Ro���Ϸ|�5�<��?t�XgK��J z����/���v��ɈGe!eW�0��h��Y?�W&���fZ򚯥����������J��SdQ��x�@e)C��ȩ�W/�QQ�^�q�c;Q|z��	���p(�g�
-�����Ն��忎�'�a�!88��#� �/�R"!� 5{kq�h�t�עU���>FI���s����!�*���Fn�U�>��*9�e�-�uc?]�7��wr-%^�ũ��s�/v��Ӑ����H��)�M
Ĥ�4�������01笍�K|�/�b]�y�B���	
�����s�|Tw��:���z��1Y㆘-�������|�]������h(�>c8����eq��C�!����ܒ�UE},�#gV�Dz����"�� "�c�M�bS��J�YG��Hx�I�kԥ���-���?v�r\���Rx�&1_>+Vq��<��Ҋ��#���4�nZ.BVi���q`i�� �j\RO.lo���92�`��*K���~Z
4;�3��h+��; ֈ֦Z�����p��w:D��b��PiUb�v��Y�m=u�R`z���]H6�0Y�4��=�T�HD�F�ou�tDI��s�����.��6�9�Y�g�&���6�u�J�+,9}v"vS��q\6о�(������4�'a��!_v>��"����t��F35����T���z�+��̪���Zz@�*X<0ɢ��_)�L�o[��B�E���!GL�9}��AF�������.O�U(\�ߡ��ʬn]�.l_z�k[:,�x����q���S7	~�j �(RvK<�Ƽ��凫����5���kjlY?���xp���D��)kT�at&�yxEE���Z��8���qk9�زT�mDg{�Dl�2uؿ���P��.9�g���m�Y}�4D/��ls��	{_i�gƤ�[s�*.�j�}���ᑧE�D�y�p��7����O��yN" ��>���v>_�j�f��?~�����`� ]�~<vok{�쫟G$isT,��7X��o�K�g����^y��&��v:d�T5�M$*�s��&�KEo�Z��ꆷ��R�N'�,�f�^u����43i�a#`mn��	�s�*�y!�҄��/x�/�`IK��</��PHm�<\���!S��˞9���=nX=�}�3�0F�$*\�/g5/X?g���1P��oG��sYq{+�ak�w+�1=�F��aZí?�ԗ��,�D�]�FL���U��obN��*�� S펥I�֜DR X�]_S���	��auڗ��[����U��"oJ2"l�>Α��.]:��	�>�kNJ$�����y��Ѫ�ė��^�Q&*&�~Mʫ�T���J>��'58wk,R��?��H��d!��#_�p��U7ȑ���Qn��f����e0p;��;���^�R���]�W����G���_�/��8���'�b�kh`/�YG����a?q�f%�q�n(Êp`�.����WA����	���r-��?*gv����ے�:$���W��wӆ�\��	��"iL`�u@�ǿ��|��vt+�����zK	�	���A#�9�ڄ過��"�Y�<�j�^�8�:�.|����ˏ?�������l�u}�E�)
����/���(�n툣Y�#�MGȈ	�����R��y�֪�����c�{X�%��cRd�+���/�NJ��%ͽ��*��+7n�`��I��y,����O0�K�XL����*b���I&roc
��"=�v6w�1���w{Ha�7�*:��-�)�Px|�:�A-�kSo}���jH���p��[;5SM�`�j��	N۽҆6,,�!�C�$�է4�4Muq� �e�o���gLv���',�,�� ;*#��O�֊M�yx������>K�e����@��@��.�v�����`���UC�e�[�('�n$J�غdʝ�훅�|��ڊ`�A��H)�`�~�=��	F��3����1�FL���{��;�g�h|��� �!����@���[B�Ț�P-��������B��UN�3k�&O��h��?��/� �ݝ�?��櫽j�'���f����Ӡ9%Z-�O�dnv�;���������F7�z��]�*��r�x���wޑn��Qq(�*o���S��|&Ȇ�)�!D��rM�ʴ���o2� �Bѻ�tP��:�|-LXe��o���C�c;��E
z�Z��&�4�B��x�շQ�s����z�XT)�������L��"��f�ԟ�h@��3��JH����nT�����J�u՞ϣo�]|*��� '�6Љ�mJ_A;ةu	�� SrN.��@b���r�zl�t�6�M�c�����.C���&2)|W ĩ�iDw�ki�^å��L$c�[j�y�T�	��K��m�r�DQ����?�]�4��i�������K��bo����J�S@ܺ/y�l<Ш
.6v���P�=��)���X��aࠊ�\���^���t���	{7��v�� �J�� �
�h����B1�˹4��s�⛺4��/&]��8?4�oVsո[c��v�~	�q�@��I�Ɔ-gM`J�9%�(	�6��n�F���Gyu-\�	а������~Jz��n�ɠ����5KRo:ʰy�񺕈�z$��@���GO�?O���r虥%K��ZE{O?ؚ����RC���D�P�����F�6x��XQ�}��/P!'�������H�n:�B��8���/b����8kw3���n*��@QG�����f�Ϲ����
 �M��q��Dgh]�ItW����|b'��;��#��x�>!d�E��~_&FY��_��8�q�h,�$o��G}�=m�(�(�a�V1:��Q�|:��ܚá0�����\F��2W���Kf�2<�v������癇=�4T��U�Đ��]#�/��y�}��7El���_E���.v5s�,�k��3��"u�MwX�GO��3���8���Y���-��]m@ֹ0�.�>h6Y��^����~��/E���"ȚG¸m�a�r�����U?�`�$��P͔��Ӱ�DK�̚%%Pt��2
K��d���W���(o:�B��iˇ���l���rE�+W�~0
@��E�YEY�z��x���$p�L�T>l_�zs��p�UHK̨��D|�&kN��Q���'+��@]/w�P4�ܯxz��>�~@T�Ti��Wv�=��=����ȏ)G;v|��P$���QBx�ә#�B�>?]:�齭.ʇCd(�����Wc?����M}%������J]��,��.=���J����*��mk�ke�J�#H�L���5TP�y?t���2��z@z��yJ��e��^�O��'m�)�M�R;u�>�����:��(��Gd;lC(�q�X9���LH����(¤��vsc���tm���9�
WKeˁ�����vԱ�X_�E�xw0��W��������ƻF:�k�k�m�b��7t��^*'���h�+�N=��].Hd˶�ުq��8X� ��1G�Zڤ��`�"i��L���6�y��w�L�������2WD_��?5F����I993���!�3y���\P#y$�,�7Bȉ��K'�qҧ�w0sp���f���bTk6���S���2r�c��FUIBa�
�R\@+�)��~�8�6 �cx�Q+&� �s�����˷13�Ah*?������H!	�$�$�~ހk|�#�t
ܢ�՟��^x����%�� B���)���Z?�p!֧���.��N��p6�N�O/WxN�*w_�k�dNT%y��Ϸ��_�hwA;O�_��ɀP��(��B�|��oO��
m?$�
XX�)�t�$$]42�?��א���y�(K7s�bC��DX�zTU)�'9�_E�8u*�}�mu�<����eY�R{�B<�i���xA��Ҷ}�����*ouI�������F���X���nd:OZ���Fg����bl�]M�.P�I�`L���
+|���N�t�-:B;�Lvۏl��/�n�؉�V�L�ş���="�K$��@���q�pg~{��cX]�Π���[��~�WI7�
��1���H��@��X��%�%|��,���F�)��L�,@ǻ�����˒!p�
�g�v@uF!֘�P�n�=n�^��W�[�2����
}k��D��]�jI� M�`0��Ūx�DE�駎�k����_�2D[+<l��	m��3'q���j\-�{�m����jF�ǽ�]�y�or]������}`J��,v�7�
њ,^3ޟc�A]�Pɫ���{w�� ���ź�Jw�'�*�r������LӮGq}�RAM�S����*���*'-b{�<)��
VibMPs���\��Y��������T'���^(J�2()9=G|Tjs�逅������SHTh��&(+ P�M��##��ؤ�G���̢���C�_F��5�_��ak�g~��N���,0=ԦE�*�4P�![h��s�A-�f�	x�����v�H�v%<�B�����PL�_�r��d����~HZ���:�sI�J��+�T}g��<aNh����>y���/g�lhD<q�p��ܵL�����'#Y���\"���0w���6����ǩt�E��ð@sR�W�,hIn��@�xY��7:>�������=�������cE�y�N�C��_��4d|�Z��j��L���x&��RI��y��	��W 6��.|JoM�VM(�F���J���<s�Tm�� ���O��@�y�UA0����ɩg<��*��Q�w^s�8���R��h��	qL~d�
0�m��Cs&�5���V����fY_UXd�Pz*�HKx�6��[�E�.2|s�ڄAe�h�S0R4�����J4@��Fj�y! ��A��j��������T�Z3�U�$M+�w�S���]�V���t��+��w��ǘ,J�-�"Xzn�Y֜�ȸ
 /�L����P��\N��0f����V`_[�_O�ށZ�v����2����b��L
�r�SE%��zZ�Q��*4Ydd��H����jR��N���me��������l�"C�iR���O�]��jYBչQ���K���Fh�Mf�(�B�;�!M"�ֽ'�2��S'z\�nN���% �#R�T��G^o@Nuѻ��� ޹��սo��tA�q7W��4;��~F�Li��J��+�+׹{d?���3hM�;"���<u���`�",���.��,���٤�����>���,������O�8|C£�O�(0� ��Փ�K�1'x4��Ք��E(LRx�m���UА���0{�C�p�R{��^ihj����\�9 ȱ@O�2���p7O��t�#\�Ɨԇ̲��l!� �C�������L̹#�ɶ�#<�s�s�AD�w{Z�ϓ�x�-�C���R���p2f�]�$�c���1=��W�rDP�������\KW��9��ଁ�tF,C�'���C�u�cE(xV��ŭ�"1��L+�%KSڼj45y:��<����?s��%��bE����D�����C�/��H�}����ͳe�>hhN0������z'$�T�O�.��;�R�mc��їdX����?}i0{1�3�l���b����˻�8q�YNb�'�����=>�Ǽjd�_��+v�Q��u1��Z����Z�кj�
�߄Fr��D���zX�!�'J}�zV鶾}���(4��Z�@��d�ˍ�����	�E	�z�o����-�|#�'�|��t݀���WO��¬��wIN�(4NYEyJX$\��L��ޠ9��%����$K̠l_�JI�e�o�c
�\l���!�o����WJ���ƀY�����r�����1%~�����5"�PK�jl�N�����N�5���g�$��O�>��lB�����Xn���DKI)j�#%�9B��\qq١�89q%�k�k�d��)��D�c�8�W3@�k
9��&W!�w Mh'�������[�m�����Y�Fۓ:� '�:2��&,�4'���3�&����V�?�G򸯾�Ȁ�TK���������C�\G]�
�z�V�pU��fH�C{�xH�z�l�����Yt�5��{��Ո�]I��8��N �\VH���w�ܔ"'j��@�&y���Z+"EI�ٙ�q�Y��9H~6�3nka�����K��loD=�[0Q#ˏ�Q���[R
��̈�;:	hE�{*�d�=~C��<J�(iO��=�!]ڽ����'���p�+�Q��h�p�H 3�z�F@6����i��]HH_���r@�rQ�&��H����(��+hR_%[3Bs�@f^�{eYo��p���tY �w��2m'�<���'DĘy7��~Tu���5I5�ȴ��˴H$L�_�p��g�z»fl��Xq�^�:	����-�ŏ4m�J�p�5��L�-�((���|��-��nCU,�(�o~�� ��Ҿ�23�	�[ۺ?�	[|�RA�g!5��Hb �eP�-:PuEܷ2�қ,/6:"Ѯ愥_�����f��ƺb�5t ���)\��/w~ݢ����W����U�<RT �ہ2�N[�� ���[�k3�������_�����w�R�,-�s9_�Z\#O� q�>�i�;N���ˊ̿Bp�]96�VB��k0���[�tl�ㄣ'��	��>fW�ݚc`
3�T�[3�΅Ҵ��r�����>Z�K�hO3Dk��d�j�#�>���#�c �n.Ѹ ���"���v2�uRS6;W�~��÷��}���A2��W��]޽��*�8C��q� ��k&ּ`���(|��K���\u���R�8����td�q��?9�YO\e<.�a{ ;l��P4�s.���8ˡ��h<��|����n�ނ�fgyl��34�g���M:���A�����a�n��#���229K�6��=�(�%��v��5��%�	h3V���7& ��'�Z��R�ۆ���)�H%��u@��)�<k��0���W��p�h�o,,���P�l� 	V��$�i�E���O�ԙg�t�s��ǯ�XSG���Y�ޒ�թC�ڽږ>c����5|�hQ[�0�?�0�T��l��hX��O�a��rߢ����׉󯽛�������+}]�1NP�_��d�^NC�1���'��!��ܻ�9ZF:$M@�v‏E�I�lN/�
#;_�P��s���{$f@���'2�,��AE��5hG8��hhW�j���'��X=א!��Ϋ�еC'7�e�������"_ӷ'b��ʑf̃��(2�Ehq4Kw�e	��#Kt��mo��`	�� ���Dn�(���]��*x �M��d;h��Z���b��f􇳴��qd:�n ��i"Q�@Q-��q�=��������)�H�v�(M�'�j��o�4�V��_7��s�}��#'No�Y&�_�LX��^�>�vX9@��{�6�\�rӐg�� ID,�jZP&]����rr�Mg���%�v��47|�FL�I�g��Q|�f �y�_U���~�Ca}kwzu���!��ㄩ���.)E����@(���$��ߵF�"�NY�WwsL6�d���!
����j��oz�Zc���y��hX�|Zӣ�$���2��Z���5M_r%S-8xY�c�Z�4�j�[qg�3KVU��j!]�����v*�G��$�i0�/,[u�H���'���G�d?�X�T�a?QV>f