��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY����B|�9ӬgY���;���^-����Ax��Q�Bf]� �r9n���%Х�<|�D�i ??K����q*��Iz�ZčgՒ�(�v�2@�=���q��9d�[587���E/��6w-s���7�ޛ�g�4�;�����tE�b�/&V��#�LŻ��S�i��d���>ϕ3v����lw��Q�[���.'�6��f>H��� ���$�]�8�(���7	ԦZ��4_�G�W�����;���`�_�A�N�i Ul�dI(��]��)/���Y�(��KA��X�-��]��"wxR\���:�\|�md9�Y�l����@0�>��M�n2�fԍ�����i-��*�JЖ�����M'��{����ŝ���V#g�V����ϕx7��h��A������|�����6�x���Gx	C�Q�Wإ�$�ޮXA��f9[.X"���W����4g�a��V�L�[��z>��f�NQh�rxPB��O\%��
(�q�cXvUY�p"�1��w�^@�p��K��K��H�K�T����5T4��`{|Vr�<����X���c���}�#!�sw�V1�RF*?>�4��� �s/�w�Iȩ�>izmR�K�+�(IxX�>)�q�7K{��'��L�����0Pl+H#�2Ć��T�-���G=-�27��E?I;V�V���x �\�h\g���M��Ɲ��d-'�x�--�?A����>���_i7v&P)������p��J��8mkh������h���! �G�J-��r�c��@��y��{g�C@q!�ʬ��n\Q*�倾�0�G�	�ȀMɷ�l�32�[ӾE����ȯ����,����rK�z��,��?���ߵA��׾���~�ǭhD����j4���<<���u��Ϸq�q������tbeYV�K��QT��ۀB�{�����A�<�� Ի+�e��s7a_!��.݄l���� @77�U��B�M�M�吤����C_T�n����81�}�?���}rgzfG鴕TE���q�{7��U$~��0�����r-��[�����Yʹ�st�x�k[��sy��x�x��Lu���Q�E��f=l5�+_���)m��J����8]Ń�������-u�L�	t�gq�i�'�k�UIJ��Ī�$�e�x���|�v����9��Ŧ�k��C>�l��N�3�e"���?^���!�,��Đ�hz�/K�~���Y�䇀iR*8{����@��z3�1���!Cf�!F��p�+">Ja>W�]��\M)��:�0�?�([�6�����2!y;��@�e�34H��=���L�>E��(����Ԁ��������6D<���;t�!����h�ś�`�*�����󵊤��ݕ��4�Z+���5��Uˉs�K�"j)��-s�70��Ά漥�"!}la� ��4s|S`u�]��c/b좂s[N��ܦ�g������v	�u��7�(��B�b���m lZ�j�P�~�>(QL�6����UͽQ���"����ʻ�hf��x��5s�;4�<k�#Y�NU��"hY��C��8�X�(�ǖ�I�b],��08�z��О5V	���H����T20<����� �ʧM�� �@A�w���)�X���ي�����e��Њ�!4��؃���P ��rz������R�s�ne��1�������� ~�QZ^�'n	�����ǿ��h��Я�wt$�/=�l���W*ou9i�Y����α0�<&2M�\��N�@�?���셍�+Qt��,K���]��0�g�vA�5=��nyDҾ�%���Z
�g���cT�P=k�@ku_�X) B+Uc�o���*D#��]�jq_����풧��Q'�#L��h_ N��w���16���P����y�n͓�c)�S�^���-{
e
^8F��?�H׈vzR���Xm3���T�WJ9�v|��ѽ��%�^j%	�H�a�����}3,����'���\����k��^n�4�̘f`ɧ�(�@�nK�j�D=��K3�� �hVڀ���q>��;!�~TMb���z?�w-�H���� �4d�gV.?�F�6�A(�7�@�C�"��B��fa�/7�"�_�n��7��&5��_0����~׉�e��T;����w~2���;��*��0�=�Ő;���U�Q�#^�h��T�6��|�r�'��R�[�^��������}X*�J�]�D� `�A��7�%��(����1y��1?���[^|O������$�Y����X��� �1��Zl�� �<FX$�O��}�z{B�ۚQ�A[��j�2#*�!��T�2���
ʟw=�x&��i�}��i�����d��o�֋;����.S�6%�67�0� k�߁=�}Z�y���,�dx�(x0��?9UcNz�>�4� 6�HF��;T۽��yHiB����l�_0��x�z�q���jU[����~q��
J��G=�й��u��x���x�z1�M�Zq(�����*oT{a鄋��i�=��%�S�%F].��l�w`1�$%��zOE�77 ��#�T*� �@�������9�XFF���7�Z�ۃ�m>A�Kb�=��oXxWECP��i�es��r8��jPz��� �4�c5�͎s9F\�ll�uy��='rd�y�Z@� �j���Q ��+����ڇ�8��+��I��At����OB�t�d
h�49#����~��X���f�&�.�7�l�}Jl@�hZTFm���s�D]�B�q|�?�j��� 6��2�b�-�ߴ�|s[�H�[�	}
~�gZW��t)#gL*�����1�)ck�$i�,�!B�,7�8�K��n<,�HY�Ш.�X�P�޿��"0]���G�/�d��-ϯ��+�2e�X0*q��+G�9Q�Yv^`��2gMJq`w�`ۥ���� D���7Y&e�}�&��u������b�6�w�)$I�ڲ�]d=�,��q֣B���ݿ�
2�;�z+�fʥ����o)+��={h�7@���`:�*Y6�A{T��Y���ٰ~����mf�O����3u�W�����U�+��#�ŢrC2�9����t�	H�ԤY�%��ۙ��e ͢�A`��S3�~����[�;ʴ�����Y�!4����@��U]�m���l�l]�围dk��O��eaS+yL ~�S'X����3W�lU�Bc� ���Ly:\���Z����n�A�j,��V	�!��W�\y�cT����J�i��N��rF�	F�~�A?陙^(�g%faQ�5Kb��u��e�7�b��T<�~6�X.��� ̽K�ذ���F�7G�{��F}��(�@}Ϛ<�Xm�_�l���}�7	�����&�r�B'^�˱�E_ʣ�O���)A��ϼv$/��rZ-*L���\��5���q�|��3M��&0i�gx\SCӁ�ڧ1د�,�eY¢^�v5�J�:N��~�Y��:���C�J� Q��6�@2�Yck�drd%����x�B-��@S�%�X1�+	��H��5:b�UK�-�����Z�iL+�� @���K�5�||�y�"*D�V���*(��D��B;5��S�3��d����+�h�p���|Y�̄u,��j�[�:�u^WTs���w{��4�sK���Q�c���e��4����N�f�&�z�}������h!y/M���p�����?[�S�O��m�[�k�cT�J��sHV�K�������6��-�������U�D�͔�����x���h����R,��{�d��"kf�wp��?=&e~����t�^��p�*qܜmU'w焴�f������С���k��i�J@}[� 5u��@lz$O<uͤ#��јm�!�K�
{�Z	�W�ֵрƼ�����tUL?0�DI�?��3�:Ծ �������!�7�CH�H GX�R�7�;�h-_E���Sd@\����c��08�3��l���m�y��q�Z���i��O�Z��^}��@a��(�ߙC���'�jloNz#��~m�x.�����!it��"����N?M����&���*D��e{Y3�)>!eg��W;�q��Zxxw0A�
E!�1� ��2!.�
t�>I��\����mc�*vֽ9�5�$N��S���sHG�W�¢��&�C��@w���著[��r�f�Z���������r�ا��)Њc�_d+��O٬�~<�7#^ǀ��yf�E��r��Ot��ėMh=������NWU�*��|\:w2�Yt�3!{��;�p[%\���;p�?�q��5��Ah(|��[�g�Ԫ<���p�F^�������Ʉ�����F؈��9(;'�bPP��[r�ޢc9��B�͇]�ll��˳T��������qm�6CKHg���l1ȵ���x�)�`�zd�g��E�'���s%���Ks���OR�]l��eaI���x����'d4��R�݅�ٟ��5��3Z��E\���_o�<�|�2`�o�N�8��D����pD7�eZ�>�	�C�{h�
�A�t�����@nZ"B�(���},�=�'i!�Uپ(���V�ԡ�bF������� #�%�5�b��D��68s�B�\��s��)�V#�,Bg����K�7:��P@����p�_Yc6�gu������r"�����<�a���aAb/�������f�PCT'{�mY(Ȩ�Ƚ��I��:�o����ja�t�k��>��E�u�T��6��m���>��M6�R���>K~�������2C��k{������mR�&E�Q$U��<�2��,hW¿��ֹCՉQ�<���q�0�Q���&.���p�Ε�@�ty�^'Ռ8�{�}������Nu5�C}�-w5�0~w@�WJR�h��:Bţ%+$Ꚉ��R���&7M:.��/Cר&7-�9�����J����� �,��SB��p��m7��R̪��0���{�w<�٢s\�	㶗