��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY�ً�r"�(t��~�6w�Ύ�(	��Z���y���h�ad�2�K��o�N��	$J�d��}��e���<?����w7<�6����:���<������і/��d-��h�m��bS���]�K�SÖ�?�Ӄ7��d���b5a�X����P���{��%�u[��B�M�D��K�T�?a1xB��<�yX�#����&��#ٟ,W�I�P�r��Є)n`v�Բ��������'�3�y��u�C��?줗K�e�u�::���ݨ��d�#Y��P(��7�O |?��icM�;�� ����N�i�<�Vi����T_B7�������a�����o\���D�^�\p����v��e��I=���vZ��҂{��{�7Zq�Q�{H��qP\�+K���v�%�8���ty��ׁk�j�Ti�������
������X���]�Z���A��?W��H�ilV1��_��a����i7���l��SE^�Y����`�R��Eϩ�u����P�{nԒ��H&�X���ɐ�,�3_;^=E$!���OG�ϯF$�I֒.�G�D�(K��Y��^����2���xD>��N�l�f�yC�nU�<�����57��K5��6���J�)(Zj\�O��͈3u{�g��}0�3qW��z��ci�	f� T���^N]��B��j�Ɖ�8EG}�_Q��
���8�FWv��K�E�%���G�~f�����t{��.�
���a�a�%�Xɹ�)N/�e��Ŵ�D�3bbڹt\�%�B�$[�1�3&�ƩSrn�9�iK�2�L�9��r�n�ɕ�b&�S��ލ33 ��|쒶�����&p �H�8�Rc9P��}�/��;�V8�i��aqOM�C�1!�����RVwY&�P�^��&U�((z
�8���Wj�=�q���\_01�:�+�NX�ڕ`��{q����5t�H����k�v��<(��4��+c�s�\٧����Ʈ��,�ag9m����ɻ䐇Qw��>�^+��oRt���g�H䭊��o�h�����7w�u�)�f��WV��<R	T(�g ��<�J
V��1G�1T��q�D�,���x�8,�Y�C���^j�S��+	��Y�GR��ף�Q�z�'g4y`�~�(�G���	;#�3��T$ґ��Q���Kl<��c�2�.ӌ�8
#�н|9@`�Z�Z�o79�8ۧ�|CQ�s:���Ϫ-q���W�)� ���'}(۬��Z<�؁iV�0D�� ���V���g��kA7����VՉ�x�:_�oWN�H�������|�dZ���c9�,�����P�G� [,A�E^�y*�.~�Yk41Л���'ڌތ�@N��hc<�P��12m,��߀�D[����R1H�ݵ�W+|�`�q�Me	��ڑ!�sFs2ׇ.�?�1�O�
j٨��׋��<>���)ڜh.4DlvjNQQ�h���~���@��������=�tx��~o�˓���w�QW�D-aґ��[j�n�<C\��������]���ʻ�� q=�Tmm)%�i��|�D�>�r�.�_�r�Ķ.2�W�Rco^��b�Ǧ�\#۹�|�q�	x��.ǝH��2N���4��4��V��
~7���:����b";k��^���-�<Ҕ�YV������皥����w<
NC��U�Mh� O�4Í����T�~0�.���b�'�������P׹U�nxՐ#@���zs��n��t��*c�Dm��pQ�y��`ӳHze�\bJ����c�o��G��V�80�-����\#kt&+���W�d������0�D$��-!��@�5�nP@��%��ܬm�Gsr���[�
�{K5�yw�hMD��[�0���ۘ���-'����0�/~_)+���r;'��� �S\��gS=2w"P��h�/b������KtwE����� ~�aE(ℳ�)S��bڄ�^%=�n3#z�ᐳv����۞nt� ����[�,��K�>0��͙��?>����V(~����Z����,�"�#�*�h$��oRB!�#����7���c�;"��
$]B
�{I�nl!�.j�z`h���Q�����S'���-�7�
�l6���w��p��Rf�cE�x[?5N7�m��q~��6�1��1}��ȯ[sSX�h�ky�]Lg�
����f�N1yO�����W�zi�o����F�ݒ����!��w�I��Ct�W�;Z8hf�C�A�s��q:�$�%�I;N��eM��{߯�{�ED���Z<G�.��o����]�x7�v�����s@��+��9	����T�>4;֥���D���w`�j!#�:�$���?:��A:���xm�^t1-��M��o�Dzd�+�ُ��ۡ�c�b����J:+�����FC�J��nDg���\"U�R~0az4����Q��Y*Vl�f}J��꩘�}pӁ���t#���l��$�3F	4��Á�^�S/���	58�AbU��i�p������d��$u�Jz�0�&�.-#-����V�JC ��jd��F�u�������Vy�}�y�y:tT��sh�������2�+X��N��V�zh�������1+�<���\��uٟX�5�ԹL�^��T6��KG��D)�q��"+c��8w*I��g	Y�*+"���션�9v�/�؇VgV�k��s4R' �s�A�s*��\g��׎�{�
� q��E1.݀��꼽��Mf8yk�,v�z��,:Ť�W��I��-/@v�@��mc�شsէ͈a��£,�M7F� �3�W��/H*k�֦���]����n�`�0JSt���'��6��8Ձ=����)���x%�lƉޅ\�X�C_Y� ���z�}>Z'M�cg/���?���ƈ��\fH�y����~dV,�6?>MC4�K|͑��l�=��E��LZ�@N�FQ�->^���>6�ũz�\�B��}����K�ѻ�Q���L�gaw�����	�/]�8�,ȄEں�XG(�<�qTS���`6�����9�*O���F�3��A��9^�H#�OwyK�T�._o��?�O#tF�i�����t�v%�j8�� ��0��H��y7�^��a��w�d��ґӏD���dh䲟�Z4�V cN���v4i����N��~}n�q1�1��A�#��s<&���s��<lo������ ����LH�B�z/9NN�m˯�1�E���.J�F���q�"�49��Ҙ����!���-�!����;|mW��f����2_'a�j	���S{��+r�MW��r�P$a9��?:��vw����ƞ'ϗC�P��RU��{�d��(��S��G(��ڤ=��o��=�cP��@*q�B��C��ha^��{5I�`�%�������-�TE7���9���� ���bG5�$�~α�t�E�7[��-�~T�Z��ٺ��a��C{$:�oQn|@�ݵCR��� �64�yE��q��F��Y�*�Y�!��`Ī�6�t�|w(F͂	կ�E��YϘ�����a�~���c
� �,Qw�c�)�Wf���ī�m�,bz<�(�_��
��M�Ǝ��0/ J���˴��aNY���Z��
�f"��.V鑓7�s��"�if$^Z�ڴe������ۤԪ�'�nu�m7�$��7�����|�B_ �0�[t���i��9�)I�����
jT�Nf����CS[<���H�.M�+5��o�Q�!]D��q����u����m�~�4K	%P��N����+2�Έx�hf�u��r;N�+ {����F��u�9	��� P���,������l�b!.��O)b��,��� �F@�y��~�����W�++���A�>�`d��7y��Ok��1��kFM����t�z\���T�,�$��쯆��\���%f���ghu����KUۗ��8�:�-g��a����U���5�Z���f�p�H��kG�G%�>���bA��Q̣:��:���PX�EXiZ��7I k��*'9��q�P�ث�,�����,�T8<xrd�?�'.�Q�Wf�7�	)����d�m�Ԡ��:��`�ʸ��_�3+�y�~��z�:Pp�g��0 �u�0C�[���z�"[cz�A\Kù��6�/بVK���U0e7{u����t"9?�Y�E�>x��U���m<��M�u`/����32�`�3�p��sO��O�ӫiW_�#�t�7�7o�[���../��{�I� �Ϸ�����d�6Sdj�0�k�@�5yRA�b}�����D� F��5���
/��]YF�P蒍��mϑ��m|�}�i�ul��_�Ks,
�˼H�ߨ�Yl�3p�����}���B`S-C��NT��>�l�bC)�=���К�(}<���"�6�poQ�M�^�C���˿Q�������·O�<���ern�^��⣺+�e$���t�`�q1�<��b��ʖ��<���7���!�!5�LUUux*��	~�|3	y�c�וJ��w�Kyf�OX��/%B�FE4&��I��g�\�@G�Q�Ծ�ŶLDDJ�fL��*�J��Vp"��Ϸ�*4�xd�U���э9�KHqa��N�G2�<�F�\պ1�-���Pf!|��h��F��3@�"�����
��sr�;��i����1��!
��̧��UZ����{9h�*#8��N|m�v�ģ�E�8	��i^H�I�,s�PT�eW���g���B�;�A�*o��<�D-1J�_��C�Q��K�sY��ׄ�TZ��&J_���oF�æ^����`^fJ�aBW����,�Уv�"7uc�i\(81H�}�AI�����ph�]�`��E罻�1IK��г�j[�;�����X"����Q`*ݤ��j�iLѥ��*ᄟöP�VM/�ma�p2��G���*֊7��;�-Z�p����Y� 1�N��������B�{v6�H�=�W�{ͳ��C�����/�)���p,!M���D�8���� �4?��^i��qM����Bɵ�0���1dk���#��G�D<}�X:��4�~0�8��g�1�����m^ثm�`�{5��79<[�=���NSI��,7$���ނ<�}둵��iF�@B"`2-�P�~�.�� n�������u��̙�xi��s9��Ѱ�6\�W�"��3<�ӧ�+������̱�e%����
>��;�Z���k�@'=A�H�n��� ��(�Yi�"�.4�}g��rb4�%�u�0O�F�*�BFY��͝��R�,�����(p�u�����������kb���-4�Q�9��'���
�RLP�xy�O 7�e���%�s�0#�"86��uu��7�G/i�ב"2G��u���s�#[=���l��q�3���j�;��I��s�\���<��T2j)��1f��J�qwN�2�3��.�~�t(�	gT�B�(f����%g�8��S�a(���q}"G`�������hjV��ԯ��y�(�V���H�R����I�����p���Dy�t+U�C�r�s!��8�����"ɉ��ک�L"��Uf� h�C�r�0>gs-1_"��!��@��Hb����w��"��ju!�g�fn��ba�%� �c!#��j�+s�?L���ڳ?_'�7Ne��㗉�l����H�/\���{�&Ѡۜdf�!/df���g�<�~��jˢ����V�1�N������d4>=��*��(�^;����C7���ힸ�ŧ�|/�<N�p�t��9��$�;�G��<6�׭{�zP�x;rU�2*(a<!ΉJ`qwv'�d� g���B�.���}L��:�O��m��G_�
���PL3(k�(���T��yg?�`�$?\Fu�����LXd|>�X�S��p�U;n��ӏ"g�$���w��m�qo ��;:�����F_W�4?X$��������q����}�+���Z��P��p�5����@� :�[K���euW��r�X�8�`TN��e�]��㓚���0��9�۶޴av��ܢt흉x�EtN�1�r�Xo1Cg��c��(|��,��(&.���[���E��6��m��_T��P��l��
��yY��9��'(�� Lqw�G%��I�'¾���'�/(W@�46|"�X+'v �p�W��j�ۺy':�.x��|���0���i�����Yٵ��X_��c�2�s�����{�(b��(@[�-$�fݽ�9@��.^۝��.�����7��8�^���R:艭��ӸH!��4�i��S���(s�C����(���W����\==tw�+l�W$5���������݁�A$~e��D�n4�T\�w�2ɿ�j��JS��gOF��ʞ,�����2�?l����t�曫Di����o�/���p��C�~��d�1z���~Bzh���g d�6�հ'0׀'�����\�2��	�{�RE�'\�v}N�{Nd���<�Q��}�"����T_/�o*��_	�r��hkQȣ�kʚ�o�S�8����
/J?��F�Qx�J��51�C<��U��u�	éG�H�XH<��8B�#�+�6���*����h����n���,~��?���L�h��3�+��Msw��ϝ��Z�.�����������Ynǣ|>r;��ll��'|�j9�u�T�9�$�Ձ���8ˇ!�ܥOK�W]�d�,>�����o׌��\��aA�<�U���H�f�@�l�-MEA��D�%���b����|���q'6�������w�ΑQ��>#� �uqd�ڿ�� Z�ed\B�|���lBS Z�h$��B����M �(:�!(�{~S�%d�������<�h�m=��~_q懃�f���]F؆ќ
"`����7@�������5���R,�R���1��ȫt�2�: �>Q<��s����@z��FL���q�-�ufwBq�iBg�"�ͻP�J�M��W���#j��T�(b�'�Ja�O<\�"\�ί���?���C/����DO	p������t⻿�Ne�Gzĵl�����	�Sp�p/牉�K[8��.v�R��ű*[^����t�6����Ӣt�E�/z��+��{�[�w�YH0vv�=>��bS��%?d�f=+C�}Zf'��)����I3Ң�2Oj�Y���!����Gt6��`�k�J�0fu���;(j�[U �7	+I-��V�u�?"Ǩt�\�qn@�R8Ú�x|W_r���dg���ד�@�ߊ�m��0+,r��!1,�O٬f%�����e����7�
�]���*e���;#S�|����m�>�(L���R�b��(W�N���63�%5��LmwX�If���� m��n���4�`_V�_���E�\���}K�PsM�[U����VZ SVf7�	�[��T9�N�J_PAe�ixR�6R����[?eYi�����������lٞ���N�@>)=9�������9�]�������������t��+F�b���!��s�0�.�����C˰E��D̝&��X���H�����	�@�����O�&��L���{����H&�4P3�8,J����d���sj�-���w'jT�P��N*ԁ\��(����pe<��ܺ�Zj�����"�&O�ڷ�������5E8�፛�d�RED��q
����X|_7�b���������z� +=���2H$Co��-��V�<�>�
.��$>�Ve�|�S"���+m��e���J���Ժ�|�"R�;�؇��Q�~�t�$�*NL�ny>�+}���<��9�����x7�����k��Y��q���_:�ٹD����@�����#��Y*�8��Q���0�q1i����}��:�}�~>�-���>�X�Of�mu��/����5��Xj�'�!ۺ�d�n�O�s_�x{µ�1�lҋ&�!�t!��Vf���p\~���# ���+W��io��a����e��'��K)��^�ދ���$	^�S�p���a9�e"Zߓ�';��ο��)�r��)wW�/\z�0��B�el�@'�)�wN��,\����	�W��S��󌩓d��ÅM��u��
X�(��>�6�E�1Ԃn�8��DY�U�H>R�N��E�N���o.lF�l���I��*���$ �˅s�Æ�I�'��C�2����@R�����ۘ�VKp�m;AU���z6����Ԃ��C�ѣa��PH���Cg4��=2��²���G��~��W�\�c,�zݒ?{'t[z�q��n�������F�/#��5&*�b�c��4����g�V�{I�˄ԥ{�s
��֜mɋ��D��TƤ�l�giR��h=��9`.l�)�1��YU��Ékb��t���|�#���p��;�ૻ3��/���!���=w7�Po���,�i��<��]�v�U�yY�?��[q�C���
D�\�pᓝ7�j���5QH���i��ZT�]���V�`ǀlk}�(�(�Q�\_�v�� ��ġ�F��J}0��ZT��]�53tg֨��?&�뛓�F��)�&ء�q�%��!A�<ثa�C�ު)y��qW�{��.����O*��7V����7�l����Qm4���w��T� ����%�n2ge����4����W��ۭ��GAk
��E	�D�zJی}��P��5tl,f�/5H�a��R��g]h8V����=
�d�����>�e��.�m� 88��{���$���OO��Z�X�����S���������n"�[S�kl��gtmW��V9��Ca���ܽs�7$�����|ڌ�/�0�Nj?�vJ�W�WmA|>��������l�D�-�\�f�7�&�}���K����ϵK�"ȚD@��둢��o��p������P���z<���CԌ�;)�8������e�S�BDp��� ��7:�DH6ת$�o�6���ݪD6�7r�'E�O�i�֟p.��S��J�m_��*l�c�zW��ڽج�Fwʔ,�ن9ϓ����y�Z���Y=��=���g�.��/[���*sٲ ��"/:���8B����s?�)z�Z-s~�����J'-;�Mt�u0� �v�m�J䤉q�dY'<��d���8�B���Zj131#'朣���؜(Ab4�V�����yѿ�T�� �	���2��
(�����*^��͙��C�����K�������"�WML���/�@�Y}��S�<�vX
�o�7��Z�ׅ����F)�~���&�_Z��#���!\��	�̦ �{T�<���,��ީ�*w��h��Bܣ|u��q+�E�'�0.}�n.����0k�)S���K
�`=�E�	-^���!� ��ǐ����5݅Wc���1p6���ɾz�e"��;��'�?��	�{AP1�|W�oI;b�?9��ي�XJ��q��>��q�L���(�v%_���1���J
�R�v�)+�gc.�dK�G�D/4����$��N��J�Dm8�Dx�R��=֒ԉ#��U{�L}�����G&B���@J��{��C7�'��5GQ�ھđZ���	�Sxk�2&zK���^D�t���O�� ov�j��y���I��eg�Ƙ���{4zz�s��2�_9w�3a�����GIC�3�:W*���l�q��Аp>�+Y�*���fi�����)��'���5#N����4�"�y�V�1�a�?2���N�jAtS?��`���x���BoJ��Vax|麑"��C4O��X��NI,&�,.��D/��N��H�j�7f������9��^��olQ{�X��El�A,Ѵ��r�8m��ˑ�ye��"����I�©. r�X	3��b{�t���J��i�e�4��{~�z<�ن)�'c=��qm��A��*�lP��<�'�E+U�B��a��j�Y�Q1O�2�3�>S�C�Oa�
��io��.�A�ĥ�l����Fm�o��'�r��1Q#�ܚ����ty�0Y.�����AA�p�ہ�X{P�/���r0�y�c���, �'M��#:x�4��8�)Rn.v�p�O�9���9���
K��/�H	����$DZ����f�թ/��&��K��﹃��J �y��ܡu���(�"; �lA� ���0��A��"/��O)U�;�n��%{3>>P��lJ;;O�H('���q=j�?yqt�/I���X����	P����j ����#w��_l�v��#����
p������K�,�Oġbf�m���"?>[j�CZ�,vI���*7/��f�	r�1P�օ��GC��1+h�$é�r;7i��o���J�<�.���r������;������sڷ�]�*�|7�7�+7��)*+N��'�N?|�	�V���VX����q%)7���b���\�j>N_mR�f�2���Fl�6Ǯ� !�y���dV�G{����g�B?*u�����r���Ad�-�Qv��t�� p씡v2n�f#U�pJ���B�- �D�E���q�̀G�iΉ���P�yv	J��u>���F�+�bzaa�O��E+ޕ��3K�=	v��H;��H�n���|��p%�?��;2��;�^m��
�h-��w�!B7����JO|��L��sHR\�B�F"K7iL��94��O�z*:�n���HI_O j�S:�� 4#�<���@�	�o�:{����;��({�KP�����,B�A�,l�m/Q��R(?<���]<(1m��|�yq(��z�<���z�ۯX��W�N"��r��� ���s��w���tU=餑AM΅���v��:��i['"���Q�s��qדk!�(s.#O4;u&�CpS�F���QI���K[u�7��O�q�дA�y�*_'��胫9�'��Β�Q�A�!��j�\v��9ӓ��� �t/�&�6}}|A<��kݦd�)K�-����0��RA	~��:�L�	��7� t��\9�����˄�ڊR0����U)�[(ۋ��ۏm�B(�5���}�ϝ�L��(w����WAQ�x��:��	L}��_(g��>m������8C(����E+O )ǭ�~0�J��ǟ
ɱ/�yZ��g����f���CAH���1P��t��^ �!Ht��wBs�V�� �E�ԙ��'�L��	�VP�neM0+��nE���Y���HG^5��'ѻMJ`�K�u��r!:}�����24
��E:���Р!����ȟfI4f��6vI@m��RX��Y���Ɍ�U͜v*$D���Zr���M�=.hIw����sM�[���"J�cR�#7-��%2S�J���˱a��wj�>|r��DSĮd��p]O�몢M�^!�J�Bxa�U��� B>�f�~��1�o� V�~9�市��G�[
��m&BH9�Ž�F�~�J���E��c��٤J�i��tq��#d�%͏_	�y3��㧷����l�<�y����E�|�X0����Fa<��:�����t2�lu��ҵ#�4 ���\p����~� ���7���+?��᥊��e�D�+�_gI�'�Ӟ�[~��/�Iu��ݟ�wJϒ'�l�V'��&����2�ѸI����-V%!)�<j���?h��t6o�/��R�� d�� ���^%/1H��ӗ��(k��S?���R*��㭧�ȸꝑ���Ϫ:�U�D�#�#*�9������%�v�.{�uu�m�i2�	�{@=o۟�!�S�� �,)i��6�����uM����7����)����~��v5�����(1���<���\\�K$��#H��ⲸݥZ��wu��|2��9��}�[��6��.
�9ʼ�Z�en���Gg�ˤ �J|I�qWWh��"	�	�����fx�Y�|��>Ȩ �Bt\nT���p��Zc�L��l��<F�p'8�c�_�a�"��q���<����xc��؅1;ğ۟�d�
,*��b�Z0�C�A�z$+���������Fx#2��?�Qݪ�ཱུ��ڞP=�sY����um�ݨ�8���� x����Q6G���\IJ� ���$$����.��\��}��d�#z��X�vi��-�BY�wً1
]5�y�%��L�j��M��R�w�����?�l�8�1�┟=�A����$���q���`p?��oR$���%݁�eNp�&n6�����!���+�2fk��K/x�9�e�J+�\_�l���ڮ{�|�E[���ъ���[��H�N���a<���^�ڨa���"�������1]Fu�$|��]�nP�p��	�%$���oxy[-�7�j�KuFƔ����o�1>����HqC�U�Ȗ���8x�^��j���DFv{ΓJ���5�ixK��B��_�O������մ3!ZE(����ҙ0.��Z�2):�������A��PN��/�U��|q�4�3ΗȂ�#0��M%��TJkL����ɇ����9]�*k� L��I3-_�y4,R�]�)_��c|�)���Y�`v��eh4�f�8co�T�t�)���Na���HYQLng�����
d�Q��	�6��7�W�a�Ix�'Q��拥��<��>��;�Xܥ���xv�������SD0 �𬜢 0_��$~%�P<�k$��x�8m��gI����F��P} �6ΞV��4LL� �.m�+����p����V�'z�����f*�$�$`4vEj'g5�ԟ3�X�90�>J[P�CDs�J�#�	xβ+���V hI$�3���V#�'Hچ�O���9�_fɂA�'Z��k�Т![��{��5�ZV��G}�#Z}���c�\>��Пp����u�٤m|L.�I�͋L� &P�3�� ��jA��9Jwo�S���R�@E�[%uKy��6v���_�u�{i��T?e�mZBS4����PcR+�mi��8����9�{-a~C�v�[���S3J?u%�k�)r�yG�����mjZ��j1TJ��k�:(�v�K7�;Kiu�:"��yS�J�an����읣��@ ����S@�.�� ��
%S/,�$r�.chI�XZX�����
���m�?��F9������r�M�<����c���&4��p�-����g6X���V���B_6���!�9� �H���J��gLu�y�[�Ü��e�Ay>��u��y$�w�V�w!9��F����M�˫B�u��)=u�Ų1:n�X��^C��^���Ҝ��"A8�3](�! �\���W��@ЊPU��e������i5�"�,�u�[KW}St��O��%�1(_ioe�L�b�bT��L������$��W����Y�X �_�P�'���V����QZ���X2�r�L�!��Z8}���<%�J߇¢�i�0h|�OC�������Ϡ����u��ʀK9���2��!�,���Y�T����
�-�%#{��&���H{�� �yY��?�^?T�<0������*&�r����'�W����g�/#ǉ�����u�|Ci�$�%�
Y���oC� �ˤ^�3@�+���
�@�m,��nYC��}_E�h,ؤ?�+��3��p�5:���os�`�=N��g�s�ĝ��!��!�9ѝ����!�����.
t}������7�3�I듕���N�faF
|Xl�õ_�n�J�ye���3�0Yq7�Q6L���n�G��o����n��Si�Q��M/7 RZ6h�f�����\-��w�������M���J=$�4�b�@5�.���C���>B��@�5T���)}���)��D���-���ü|�^�$/ɴֆ'ꭵS�)�
0�T��I�lk!;d��U����o)OR�AI��Y�{��;�)�}��B��B��)=28(%�P�ɓ����ab��l�T��?�n\j\�K�Vh�I�������[\�(�&��⾀�A��z���A�w�Ɗ���RV�����8�"+Q���e��W�?\��WK*��j���w�}�%�#ȫI'+mV1��Nv�0@��l�9 Z�L�)Cs�C{��l��H�k�w��2���Ϣ�Wgw+!��od�n�Ofj�;}��?�W,IC��S��Y��hD�-ƪO�}����M�=�d�۴7Y��@�����X��9���3k4���7�D��{pONB�� fnQl[��BZ{����K_���Ѡ��=�Vt.��'��Fj=�"0�2���u������m�)&2aę�]<)�(�"q���:bu-��@����U��Y��L�Ι�kL�!U]���{r��{n��MZ��3_���-�N�l����yDm0u2�#0]�ֿ�<�����U�<�9p,��+�d� L�YK �`�$�ʮ��e_@�J��-�_�NYmO ���_JtU!��m� Ur��Ħ���I�k���I�M�ry���$��=B�� �?������= [���\<�UH���4����?B��⳺�A�/�P9�S��J�Fv��L��l��7mC��PF֙'MJ=�+3]&`\̟j�FJ��x~)���2�Ԫm�]���
�F��w|�U���~xj��+<�}��c=r��"����
K�{���|g�ԩ�z*r�G2�WS��LLY�4���������t�Cp�\����Y���
=��1�"�O�o/A�7�����!4���ppS�����M2�?����X��jxP����!>�n�-]8������F�h�6�Tz~�0�<X�\}#9��F6�K�9��uT��И�"�ż޿�AeK^$��OO.����@�u�x�I5�}�1^{�՝)`�ц��aΝ�l�9�(L�̈́r\���m�(������R��Lbz�F����M����w��������x�����ZӽC����1� zݡ�_�ߔ��|n���~P�����t�{B��.�2�RҲo�kh�N=�18�}�ߜ'�w2o��ɐ[]am8�Q 3��V��	��STb��N�X�,��a��I�����)Ɇ!����"D�:|~�yNƝs��FOP��,���Z����:�g�;�ƕdp�+�&��WOC:���������bh�>n�O��4fw���]��7�w{��cD�1��pW蒯S���a2�DDE�?��j���M�W��f^q"�K����}��N�*)���HƆ\} ؟w����^P���Uh�n�%!9�N�D�_�s�}�g� ��?Qk�ю�N��LY���@l�ў�V���6�O#���k�S��� �p��q�5d�ם�O4�ih=�X��c �z/�]��D����d�P�Z��u���f������h�Z<��%���������_����JY%� zY��>�F��$qrm�6�#)IH�a�����Xi�Egz��.>�R� �ө�����]��N��7����<"�fC�\�2�㇕w"��v��L��t�W�9�/�����ש�~y[g#m�x�"k�H�@�x(�oO7(\]�U�hE���K߄��S�M5
��\�S���
���7D����9�%�K��mp�<;��ދ���f%
ܮI\A�֊�ˍ�[�Z���@�$�lٓZ�|�l@�N<���$F��8��1/6\^�y%?����0�<�VG��r2�>ƹ����d�E�Z^�{������ �$�0k��7~"\l��E���-L,Ry��}���S+�a(<m����w�ک�A�*3��A�{I��hӓ���]�F@�Z\]�[�g2	�f��0�K�ʡmS8,�H>���Pc¯�T�!��v�(�� ��}��� *�&��)���j�wR-��)>���W�Mƶ֭wt���^.�Q���@�yi������YN�?[�xm0@9��V+u�+��қ������ �`J�sZ|K���a�y��읬�kBt��"6�(7��`6�{n��{��{���$���U����2��щ�;k�j��Pԕ&,��`_ ����N���/��o!��7��z�J�5�{NYi�#��Mkg�ݚ�]	��w�j���XQ�i;A�}��Y+n�M*
�R�)˙3�� ��Y�k��!����������j̊D֦�<�o��}�:Tk�r�򴙔;���ܱ'9��i��+��)���H���kgʈ�O%�˶�6m]��}��4�Ђ��g�j�U��&�o�>8h��B�M!���v����	Q�Aΐ�*V�#"�]T}�YB�o�=�>Ō���$c*��V�xގvb︢�ʤ���X��� �?���"5��V���*����&��� D:j8:�͜�?	���@A�_\h�>\���N��R����Bm��Ib��S�{ #"��d,P~��H��{i��?3]�0n���<�v�Rp@\y�秓D`Loh��Aw�Ś�O�E���p�1DB�vl�*+�Ǹj_Hv�%J�0���6]�/je���*l���q��L����Q�R3�q��N�@�G`�!�7���i�Is��D�0�,��#���\8��L����t!�y��7��
V��֧�5u5�y������gl�� B���1�2�84�|�{�낮c��Y+�7��-H�4'���/)?p��00�;r+ ?�q���S�j�q��+���T��c�t��C?��:P���aN�PŤ�k�d�M��+zW]@+��P��Im�)bZ�s�J�_�"+N��v̪�����l6��R�G�G��[����oHڋ'�[s�D��|B�rt���c��k�"���i�n~���'�c��;n"���D��}�W �Z�M���ԕ�p�!���!��Fh��_[��g���R������3�f%�3P���)8�������Ha�d,1��װ��������G�M�>�J��6��&��:<�bV���U0�am�_��F�����g�",���0h�3�/�}7
w򍸸݃�+�@�yhWQ֭Pj���P���5�3�+nk�!�>�4}�A��dʊ`��ֶ�#�ߣ�ܲS�V�D4�W�	��0�pizn<��AL�Ϻ��e�H���;��9а�F
���:����:�c6���c��wf���"��8�dU+Q����5�σ�pa��[���Ҭ���O��)%T�'lZ�&-�a�$%{�#��5�����n�?���m���-,��g4���Þ�r���AO������΍�#�Rx���]!��M��Z�-��^��)��w䋫�$7*��:��I���G�,/w/!��3̵�p���@|��C'<�Q2�Oj�
�Mj���vk�Vw��j�|�����9Z���ek��(���u�͊^�{�#���
@�p��}|�ą��O`�%��퀜�g;$���$�����9�p��J}snҙ���7L�3m�®�m������i��,0����j%����[��1;'�������b��CQU�m�t���7	B=�+��n~���e�cS�jZ��84��.�	<�n����'o{��hK��>�}�m�B��k^�e�����d>t��3�~ұ	��%q!����۾Ih���䵪Ƅ��E�>����[��bwc��\�QCv�w �A�2#F�!��뿑��$�/M��U\ҥ��6:�òfc8ߪ!�^2��m���1�ޤ�<���u"�\�F�����w����'��9N^��<]�x�)k������������t����6��)u�l$"��x�Q��}.S�	�N���e��gW����5���&K_}r�7�O�Э�5>U�O���\}�R�|�ҍW��,pN�^i�������Ch�ѫW����"���8G/E����
���@����7�*PHsi��/�е�$�Ȑ�L�k����΋ɥ2�e�(��^gj�ڙ�S>�m�r=s���
�c���z�L4w������s˷˗�<X�(j�]�����V�?V�&V�X��|��DAO��O� ���L᪐�e|�F���$�u-O�uƶjE31�f�崨It7��p����]�_
db
�p�<��9O](�ޗ�9�)��G<Q��q��&멠H#�}7�#��j�	+8��/%����=���7~Y�A�7E(�H�1T��ֆ�}Au4u��;���';��#�3Pwv����υ�+�<��Mqm����PWYX��a�:�j�oZ�x<
@n����t�Z%ѤՍ����!�'jpm�Ù)/�x�߰4�2���ޘ�p��G,��G�t�R?Q�������D݄�����d�%W��$��s�����Hp�,����j̪���!���K���A��y��-�
�6�=�N�YM�T��.��rB��䨿�}�xT������+[`��8���x�×�P��P��l����5�_��/����A�Y:�����B�u��o�֥t/��w�����[���Y����Z'��������J$]�{uh�/i�Є��8=h�ښu��j~��R�R���[���[��M�	�-%������UA��ә��/�N�5|���>��i>}c��[g��%5ei&*FN|N)�\#t'n��0r�wT�S����TSS>Ќ,g� (ș6g�T��������K~�e��N/IG�3n@Nt��/T�2~�s#���s����%��9��&n,H�ižM�����$�'�˫����p������~=D!�^��F��:Z�/�+������?��:�I�1��`����t�^)�nAh��ު�P�%,��$�VE�z=�[h����������h��f3PϦ;7�wY��"%�m�M:�A�v�����q�����3��lt�����$F-diC��G��բ�&�~����ڸ��[eLf�_u���Tؠ��q�L\�༚+�H���	�S���E��\E{2HĊ��C9��r���=������i�}��OO��0^��e��<֜��[�F�~'�1z��[� N�9��xP.�1c�L��0uFxfϽh��Bv&N�Jw9#T���%�zϸp��|��1@%h6L����fq9n�Z�y߸�SD���rS ��Ɩ݆�S
��Out3�#1��MB~����b�聚��vI�X�Q��[_�d�gz����|�(K��Ұz�6���] �Byv��� x���J���ư����΄���]ڨ��E)��μ[	�����X���3��t�WD��N�6�PQl-��S}��M�Tf�ߴ~t#��I^�g�5��ߗ�>o��X�km�LA=7�>e���5ɲxU�u��5���~ߠ�7 ���̐�����a|��X�������C�5���y`�R}oa7'hkLb������Y��Ѻ_)�����Ь�`�,_���a�qT)�_(/Ft�^�l��j7���e���X�޳� ��f�*q��}�VS�:1���D�K��5VX��z� ���}�V}�ZG�@���%�� �^]� aNbٗ5�Bwxrm�h��	,�;����a�|��i^��^>#��[���؄seV���x�����X����ދ��^�B��[j��7�%��	��h�Acp�6�9�T)5ے�;Q=��{��3�y���QP�\{��U����wb��[D�ND�����9��q�b����u'�>�z�&�M�	�s_�4{���}r[=)��/�����d�L(���8y^]{�v�W˖Pf����q���A*��ɳ��S�7��x���ZT���~�`��]�W!l�VHp)�%�/"�sɋC�;,	$��4�V+?s���7;4ٸ]�}S-W�^oy�M�(E2>���^��XCd��dn���Q}I��0�M:�X'`�7?��c�=�B�j�P��+�]��'0k�ޡ��5�K3�KO
�֚	�%��&�\���!�y��{��7g�̯�_%W�'Yz3�����V���ܮ=�+�4�1~�Ľ��Wld4׏�Bu����v2j=C쀷[^p���C�+��z#
M�x�;��1[nLP����˪a��+�8	��k)*������ɡ�Rc(�w�)$�'C'M�?m���9��;lf�Ȉ�G�T>��r�P��c�{�x�R�
$���9h���S4�G$�����B�`դ?�d���%}�}~;P��X7=��@Д yw޾���� ��'�N���j������}�x�:�c��p���bѱ�K��,*|0��()>���#���	��}��W�i�� ��ӁK�N8,7$0��>$�hT�vN� �z����!���m'�ݸ���O���!zu-r�!�+��gӫ�WG�iS�����/�V�'R�Uԫ5f$�t}[�s:'I���6���5���m"P�-7�)��׮�����:"Խ�5_�^�6xՀ2~��&v��j�K�������Q��-w��ZB�yú��kX��j�u�7�;��'���}��e�p���na�]8��DV�̈r[������t����Q���PQ<t����4%��ֲ�-9�Ԇ�kDP:�_�U�:A����h�ﶯ�E���s�%;L�zJ���c�a�=2}A�>�yZ�4aÓ�La�|�:�-<���H���)tB�K]8�m���E����k2����yz�Vx����g�uxu��J3n=߳I>�*nM���V^����y<m���y��˽4��p"�V5B��p�m F�_��Y�����c25k�_��Cy��~��b}�*��T��pvOu�ȫg��R뒵�-�5�S�J��2kZ-O)��x�H�É���^�o\��+q�{���H�&����r��qݷW� !�7�k���/���?�6�<���ݙ>�&���[�@��cܪ�9��7^���Qa����t��6��ԑ�R���l�Đ*P	 D�Ŧ@�^���F�2�Cw���k�C����xz�I��O�Wy������NS7F>Ş&���Zd񖆷�]�R�%l�b�]�r��A�}�_����������_W���G�<�Z���w3�6�0Q;�'��Y��s뚔	_a^�tH� ;�!O�"�L�m���Σ� .0jh�+vH���|�O�O�ip�H�9��ߺ�(��M�p��o�s�������&���n��L��o-H7<��Ӭ59`���n���g^�3�n*+��p�����Ņ/�EX��QfHm�h�Y#��HSw�)�xA�F����	�:$�4����+r�+'3���К!"S���e+�_�HH��_�pZ�����);,g�r6�D�d]4��_�	���
��Q�{yٍ�s/�o���	V�_�0@i�氩�'D������o�1��Z}{?�7��6|�9-�j����i�i��;�D��I}D�ݕ&�=̡�g�}J�4O���7��nW=�����ph�H���@
5�uCQ[�^R�'%Qi��}�v���/>
��ˉ����?�����v�\�I7U,���_��J@������4�P9�t%��v�]E�� C�@@��Ѥ��B�.�')%v r7&{���t� ��C*By����N
��V����N�� �
�ya�qV��1������� {��&`���v��^=b)�9�j1"ޜ������hDn��2���� kb��� \�2��D	�� Ú�yR���#� ����H�+��/VS�ֆ��s.1S����s	`F�7��=���}<��Km� 7 a%4&m�eh�����l�Q[�b�>$�7�t��?E�䂧-�j�w�Z�:��ƺ�����5=t���\����s�))v��\ˉӐD�{�l�5r4��u��_�X�>IqW	��S´P"B�g��Z0 �V�)z��
��e�v=*E���3�#NDߑ�8�yD�ļzD��9�s/7q����D=���Z�'"Z�\ r�����<��_k���`R�D�B���K�w^�1(��Ɗ�	�ޅ��T����hT�Nu�i�Y��) ���<�a�\���>�E�Y�S>Xʵ�o���9�N~��ɭTzzBK�׾�ML9�0�A|���&_\�8�dw3a Iz_w@���N$ߕn�Z\Rz�4����d�-��4ƑSm��6C.R|/�(�7Dٮ�tS�)�.P<��r�4���)bQB�ѹDa"A��m}33h�a�g���#������"�6p0���#<���У/`����6�L��6e�����#�����"є2�K��tS�c������R�����cbFz	a∯������R��h�g�&Q���G'���<����}YuR�M��,��v��>�-�f S�?��2��Ɣ��^�_� ��׉�����Ӿ��D$�����P��d��I�[�>�� ����pv�fO#<U���F�%��+�1���y9Mk�޳i�鑷�����.��l��5BW�,JV�-c�%�`)���c�  ���,#hVͲIJ@Λ�\��)D�;�m���}V��3J*��R}�gn�n��.3l0��:��}�lȬr�]�w,S��Y���71G3�	����9�u�ue�͐Q��9�s��__��Aoڪ�hW�m����k����DBC)�
e��{�D�**��<��Dcw�V��qۜQ0�<~4VAb���h�#vB������$�������IR��-d��Z�iv�Y#�� /ĤP�Вe�,�2�)鹋F����KRh���3 s��u|�J�`S�jA=�
���ϙ
�2.���;0j<��m�P�����T���+�����GSj`��J� ��eB��U=8;d]�=�?�%x䗘��ߞ
��l��H������Y"��-������&��죧hf�w^W�������MMLۨvA�?_� ��u�`����[4�����0����~�^WH�>�cRG��Z>���.��c�p�lKz�T�_��1�}��g��Mk���Zb��-�d׏�8u�sC�T��.:�Г\t~兰�����]�:�^?6q�m���2s�?i}�Pߪ]E0ٓ����E���Ԁ9�W����;3��D�_��6x�ˋg$��l��	�>����MO	s ���n��T��_�ʼ�<��V1�m�]b]�eOj�
�����Ҕ}k�s���t�6���k n�%�ס?����Z�*��s���d��j�n�͘L�4�,���؎���AR�oJ��f������EW�Ǹ_�[�@KWB���t��W�ȡ)L�8+�14K�:��/����:�)��g��(�k^�|Ƚ���T��Ϥ���B}J x�˻�	����%���|(����ɶi��7��a>� ʣ^��r��ݼ��6�_?�io(����Ҥ��3娑}�f�S�i��zw�{�5�`���!�Ҿ0�/Yx�0Ĩ���
�7R@��%��C0�d3�9EsE�O@+�1*���CoZ���W���7k���K�ֆŋ���SV�/M3�
Q!�~J���/Gr�����9�cgD�k�qgK����9�-�T��W�sD�A^�v�}�у4�����M9���jϸ�_M�������~����=�k�myҹ��p�f"V�i��z�)�s]�@�z��2	}=���֖
<�0�Na� 2T�"���������G�%�/'E�L��ًE\��HN�)v�_�&r��F�M�
xhqCWs�u,���}g8��8u�!�b�J�k�����ʬ���~���wE���KR���m����}����
��9�6���*H���؋H_�,p^����{�"a�(aRnO�E^����^��O���ĵ�^���*$���xs֘�<,ny�r��D!Nц1��b{����Y	c�ʍ"~I�����t������w�3:s�9l�z��Z��)]3�ܘ��*�-��L������y�%��KF�M9���RS�]qn�/��ӰyV�\ր��M����d������g\�b�w'��'��QZT��%ѧ� �^�k>5���!Tn�/�"	���x8!�I�����(kl�3��qr9��ahv��R��� �dٌէ홓�����P��501�Z勌��l��\�t�Ϋ��K�dB+������0�:�,gc|um_�1�sK� �Ӊ2�n����̒�G�"։�od'��t���o�2p���\jC�6K� ��.e�%� B�=�Q��ً "2��I�i�������H�}Ϫ����I]oO��D�ޛ:Q�Gs�[����4�~��QXz=`��R�GA�� Cɖ���F�	���8��
�G�#e�c#��T��,�(i�����O<�V���$c*�P�D�>hPK���@<�吠��8��Hl&ι���Q3T3	62�!)-���l���F4���5[{g@�61g�9�=��ӣ}��F�?�����������|�ڛ�w)O_$ ��pQ�ә�LskT��c����N K
2�۰���)s���g�GÂ5�.%��s>�aR��UjOx�O�[
��o�3MGdwNY#�ZV�ï���fu�F�]���O�ϊ葐m:>�5�W灩d�:�����͠�\]�Z_��%۵�c��0��x�H��zPgȬ!���7R�j�w���C��3� >�9�5�Ϳ���Lg����Mb������8�#�f��kx�,;��v�o� ,n��BKࣛq�	�2���0#��=������
� �e��L�V^͟+@ ��ʉ�t"�=��|[��hr_ሓ�xpQ����m*���@��Ho�y��������r����f�/`A����;J=�Wj=�go�d~�Z�*1�^~�]&Cn��6.��BY �l ��!����kuAc��x�
�n�H�@>�4��^r�,.��ͺBtEH!�E�4k#�C�]��Vp4�O�P~�8(�.��M�����/R:�J����h���{���9(��+�I�1�J�/v��W��݀��R�{�(�̡F����
�b�{��Xt#�|�$�2��д�?��
#�-K�g�*�J#u�ѯ�zH'{~|��<|��t� ����G�FISI�Q��
�[/���PA� ��G�"��d\�Sk'E���؁d��kb�hS��+_8���4ě�+���ܷ�꬝��ұ��ݞ�P'�)[�cS;'P��ʊ�c(�RI+"#�R�_����ِ�P�ˇ�`��F-�UQ�y�nK�ɮ�Z��W6;R�4�L��h��-�䆗b���g��s^���!�GXH�+�);��rHCv�LV�ȇ��%�͕��U��&����T����`�����)�6��m;bd����<_��\�Pms�/V���B$�2���0}Lآ$7v*,V�q�~���PO��y����e|n4���MJ�%�%����B/nD6��W�SR~P$���D��6�z�۠{M����X}z�w�O�Yy�%`�Dá��+��Ze�#�1�ҞX�@�'��!�&��🰹�.M��y�)л�s����`���vΆ]�������z�Rj�e�e�]رK680c�>XVH�V��I��|Y$TN��*�V�� ��~%o%� J��S"C~`G(֜�C��f�a�;�j��e��7[7�<?"��Y��B}��Se�����oFuU��w�L9-�1�<ޫr�@�RQq�\�԰/�Gyt�DSĭ
򇈗��)�R=���ΓF��²�܆)���q.�o�9�2��^�l�P��zҠ'&1X�ӺͰ��s��9�M}�]�)~�Ö�@cg����/�گ1W��bR16?��饏B��^$�o��;�T�Ǣu�?Q�/�~?�7�$��d_�"#b�%���Wv;�@�;+A�kM�Et����@�E��$b�"y`z��� V���Ȼ o�G����-O��d�l�@���%�N�ĩulc�\$��*7�+d�m��!�G]x��5��ZNU}]�u��a����M�IO���tz�Ε<�OJ6�FO���(A� &䛏�Xf�z��"�z��� ��m��3�8Ɛ�9��D�v5���*�)yJ�o�.��DN9F]P�d�f/��&H�i�ŀ 1oJ����8��(���(��Ne�7��o��YҒ_3S��
�6ɵ�o��\�#+��QS�?��v�'�>	����!��k���>	0��܁�E��G�{�5]� ʱ�*��:�<�v��)�h�{�&���JqSeI���as��.��ݔn���b�����J��
��D�gD{KH 7��z�e�T6��?�в������m�vO)��E�-�p�����"��1Q�����_l��W{cQ΢�O,ߺ�Zn�����~��������P���:��W��d��S\��5LL�ό���͜�k�	]�Q��M�����/v/�vdy����Ĺ,�1j����r$1����#u8h닄��o9�$�T\��&3�.[��W�5tWe������AR/�2��t�M�b�U{M�Tv�G��_��<0D'�l���6)Vo�O���$��b�>m
N`��y��̨N��Z�&$�p:'ec�ϤH�%UIⶻ0�YH��I��^��ݢ�Ly㥛�NS�M��o:�<��0 8���R�r��?v鹶@�0Fy{�I�SW�4_wH6Ft��=t�3�λrW@��;cȠ<&@E3��k!��ó%��v)����D�Wwv�)+�$�ЋLqb�nuF���eK 	�����O'Ƒ=V%��}��MK5YL��We�J}����=��R�6^r�Ij���#X��m��|4V�V���Vn7�ډУR!QT��y?�EA�I�]����lS�5����>���K�pU,�u�SB��8���s��l�<���5��5
�?����ɝ�^��tLڗeMW�,M��e��M�R�ک��B_)�Zr~v�l��m�7�&@��]�S�P�}����s[/D�Q|m�1����5Qs�_Ot�G_� �v�����cqҲ��v��XP�]��r+\.�.�*+��0A��,$��͑Vr�R"������,��,؁�D�ձ� ���0���)����e���.�G��Q=lZ�¿����Xk�J��[݄�o��W_M/X��i�y�A�mv�R�_�e��~�x5���.+���I8��3��%���ci
���t�԰\����H��*�d�	l���aK%AŜz_�{ML�n�-�-��̽L�������Vm_M����-QBO-�����)�Υ�I�I�?��E�m���cG(��]�9듧j��������	�6F�y��x���#�E�x����WI�DEi�H�g.%r��W�7f3U���x��!w��^ ���S�tk�����*d��p)�Ԍ����(�h�A�]Q����s�Oh9�P�J�Ai�X�(�<�?~#s"�ȼ��]˹��]~�}1�5�����3���l��^�-4ϒ/[���g���n%Dw���`� d"I��L�
�v�e��r_bV(!8#���;�
i�Hq�������-�Q	OVHc��p�`:�Tm�$n.M�_f���		͈�_���+X��'�T)6B�Fp$�ҾvY��5T�T��A����͸�@K#�.:Uj��?��P����m��=֪�;u�pB��;�'%�v�)�t�X���痵�����tI��R��32��I���&�J«����G�G��?=���f��Y9��x4<�%���B�)�Z�^���ϫ����H�r��R��/W�p4�G֖J
^��lA��xusȣ�`�=㚵����BC�	�8\ �T��}ӈV�˷����3�A����3�iX���lw���f��m^G��R?4�>���6��- �l�<0� -�ϴ���5C�dQ߄�{�d�Eqyv���K7�B�7O�k�w��@�4#K�� �/��}�ͣ��rӐ	�~d9n/�.�%7j���U��!��۔�������wt���ǿ"i��C1�@�n?)*K��He�_hM/#���Zߙ�V�X����K�� `W��Eq�ж��+���(����' ��Wq����B�^e'�&Rm0�HP���o�%���μC����v����b�J�ec�=��8T*������~��ڹ�6,.�la<OQ�9��<v��g++��I�*�N��z{n���G�b���=\�p��,~g�������	�b��pDn3��2���6%y֍?��2ݖ�)��E�ݡ�D**4(?/�1��\���r�o�sCЪ!: ����I���d_�wf��{a9V�d��z�q6���AJ��_zL��:0�	���3��g;�m�u�I�mhtCqI�u�d[D����C��%;<9�U|0Z��mC�#)������t�Ά��L%q�V�>�<�y�8�v���OHpU����P+�O�7[���C|��;�>ݧ��4�@�>�%2��B#o�)b��(�+���o�迄2f��6�w���nX*~���9�jZ���g��ˀ0��S�^1��#��E��ܭ<Bj�N5�e�;�|����b��@y�S{A���]�WN�P��]�ßj�r�:�Rܧ��z���֥�YP��v��% ���gUm���On 8� ]��zrH����F�����q��%/e%IsA0���ޮ��=x�Z�(AZ�� �8�t�jF`���K+�f#R)Qv�W{����n+%m�I�M��2��R��s8)o'1	�|n��"��"e1����+(G��KCq|��C�І������_e�I@����)���AmW×�d��
���-���ި �eC�4>�=7?���<���wx9���rT����Q�N��Z
zdo�탷�=Z��K���f@Uf�BB��(Xa�v�洊��������0�e�~�6���t�����G��)�"�>�g����G��m�ɓ���ݮ �H_�����o&�B>[)4{\��~��t��'�p�և��~m:��%��A�Ǎ��,d�Ƀ��f���^�暴�U��eg���Sz��}5M6�B���a�����H�����\<0�͔�st�]�\�����L{sӂ��6Ǟt2;~v�l�f�	�{�|�|���d&
���%�y񐎂o	1ٌ�~.~b�T����5�7vW	��A��Vɯ=bտc�;8�����)c#ν&V�f{2���ŷs�t�v��Xm�[���{�(�#�X����!,Ϣ����Vi|HHH���3�^GG�R(T`��k\��-����ԭܽ'���}�(��<(u��A��V��Ǡj������zqF#�<���R���,�8�c�}C19�k��Xj�ӛ\�%�Ʌ�)F��,���f���QCÁ8�SjU������5��bL[���ˈï�G���-����RV��ʜ��)��� >B�h��/>V������I�dʨ��4�V�XGVz��5��$�X_�Ay�B�hH�-Jdֲ	iEHrxg9왛+�G�V��zڒ�ɞ!´=T[��� :O?�����-x> `�� %�HAOvYȻl����O��mE ��܎$�)�X�L��]��>�2'�-�'������vJ^�Ѡ4Q0�����l5N���`V�@�����2�E �t�$\R�d��:�h@Kd�B$�?�!'&��N;��Ss���h��}:��F6х���ڥ��<�=�a�ˍ�?��89�(�SZ��n�e<�@D��DR���C���?�}	�([7b0Q��q*>kVA�j�9)0�%�ѳ�RMnW�ՙ���i�
g3��S�Lj������ǵQ�	 S���5��G��ޙX.�����C;���^��V�(KV�I�h���&�. ��j栛������Z4�h��RV1}�Q��������2����	�W�W!���lq�RS	cOAR�w�����U�o&z�B���	�1=��#�D�R
&��[�a,ٓRxBl8h(D�,�Ue����Śx����(1���B��&ߋǱ��L�V% �����S�Z Rf��b2Xb�H��*W�.�8�2���սl$}\��e�˟`
����8tK<g�G4P/����]-�?d�@�2�����n��@z/���ٕN�јt��\�]1���[]=a�\�8O�v X��^|����pm ��-*Թ�+q��9���8��툄�qγ.��Zz��%� JLf֌���;x���t{%���U�]�s�ts[�K �m�3C���c��}\X�e�jn�qLK�>�\=�Ȧ&�(��Ȱ�M�7y���~��Ū��8���e��u9����c}�g||��T�3��v����NR�y�V���:��K3�]��XSY�W�O���I�����	�z����o�,k�ĪO��9�,��j/dqR���׵0c��4���6�7��ҕ�K�=�% ��3����ۨ�C(H�A���?H��pB a߱�p$�q�2xC���FX�b�IB�­9p�:���#m��8�e�S��(ka����j����s,��:�����K�I��&�	�Ҿ�4�)�
�Ԅ�r@<7YD_kB�Vp��Ͻ`��V�q9��dw�<�m\��8$ ����/l�b�iL���u�\&`�y�Ơx���	�w=$u�0'��֨�!�Od��NKzy���x��d�w?*!����7,���0-u�Q��&�"��V�_�����0D��R��gW�����$�=���n8��u���ٚ�ߴye��p$��2���|'@[�o�]Ym���R;l�Λ)*�_6wٗ����ܩP�1��_e����oB3�$FA{���u��W�g�����\A+~~5h
�����(�BX��v\�bt{����Li:���W��ev��x�"��\��4��j��Q5q 6�fC�#ê��ϳ.��ăzSv8&���l�m�w�C���IZ�}���"IU�i܈b��=d�U��:�b���oOHJ���$����h!J���? T8'?TzJ���ߊ+avZ�O��I�%�d���R�k�����<��;�ܖ����Q��b:��&t�I�U���+����SEe27�E~
�}2�fC;(�����Ḟ��{��$�<���R:'�!���O�����re�?��J�۟C!��Gk��:ɛ6$���, �6D���eT�3���e#���]>�51ʛo�>d�x-:+b'�%漿aཬ�7'� !���/���xM7�>�3�H�FlKQ$�@,�\�udoZ%�|�繳���G��Ɇ�،F4�ƃ �� G���(yY�HS��Jq�gxg���Z� {3��1Ke���Φ��
�6�`����5�)6�0[�צ>���~�r��u��p��(\�/��sv'��d5�D]�Jeζ�<-�F�zGT�.:��'p�}�T�"�Xp��g��jm��ؼ�?�:�JE>�������t�Cd�V�A-��v�t����6�|���� �Oe�J�Q�O%ƀ��#��e��)D���NZf2X��]V���Qe�R�i����tBX9�q�O��&,8>��ƹ��
+Rm{,�����t�C�|Y��@9৉t��@ip�ae�6'�(��8&�M��X�l����V|w�n$�ڻ\�#1��<$oa�� �, � ÊZ�65�!� ��cj3�{�kX�-|�\c��41	LVG��~�:°����ƿ��K�Dy�	��B��p$*���R���`�y(���3�-���b9��h���S�X)_5�
�6���*�@n�z%dEx�	����<)�'j���(�HL�2��-@hN'D5�:~�1����S. (y�0��Wr[�<@j	.�(<��;��;%�1����wP>�$t	��˥�uM��=��J�=M�mE��C^�pA�}¤,�ud�;������ϕ���)d� �cX��T������߅����=>���P��,�#���}�L��9zI1L|:n�Sg��r�F���$U\F�;��{r|}tW(B8��>tH�;|ZZ�� /�~�1��L 	>W��%���[���C�4��Tol@J��yo�=��*F���e~̇����R5E��4�c�RH���Z70�Q���XH��Y��zK��D��'�۽��8AgG�@fV����Ɛ`u�*#��3�ߎ`D�JҢ�cO�S����r�;��V�l��R	x\�ik#K�DJ���v�e�䥴��Lj �a���$�%�1��e�ߑ2{�_��5J��SX�2��yk�\>�|ޗ�["���J�ZZSC�b��p��(��$-��{��_<)o��u1wۋ�� L@SՁr᲻�W��E�#z%>}c�� ���>RC���D���Ҧ���&��h�)+	>:V�'�y�
��''ri�A{���:��}�5���o����W�E]ea�rN��$�,�'YG���QC��%� �f,�Ց��9�&e�,@"�(2��-��izVu&�Ps��7�G��Xі���j0���K'���]�Y��<��[qGD�����ʋ�Usjј\}�r��q��p�&=��^�#�9#+��1���[4d��M>+��� l20�O���p�Ɂ�����"^c0�� jP�:[�q-w�����ZE���(��Lݎ��6.I�Q;UO�C�&�3w�CT��R�8[;N��\R����u턨Sy7���g��o���7f����(�kF����ſ��d"�'����q��;W�2���JE�j���"kf65mof�I�m&�c��Ow�������M3����x�1�=��u�$��xL�<oc�a��S�d��t���K�ӕ�����{a�z)�7#�l+��:��-ć�Ӱj �A��pKށo4�*�Л�� ��;y9ò�h=-8�Y�kI;�l	�|��HՂI9�[A����͏s��S�Q�Qs(q�zi��i�Vc�<{�_���� �����'��TC���vg�dowF-wޯL�W@1���yp]|�-�(u�'{�`��+��8��WN-ii�o�ljI�d�P�8h?b�Hƨ�>ڥq�.X)�9��RNO�I�9W�٦�l��բ3SM8��:a�(�ԘҀjz&���:����^{��"���b;z�#�pѡ�=1m He{�y�M��!�@}60:-i~�_�5_f�ͬ�����h�����:jVn���\	n�?�F�N�!�ԡ����d�N3/��;4(��^at�ŋ=�{#��˾��m|�����{�U��,i�@�աzL<�
�������sX5�X��-֟�&ax���;��"6�� D�ʪ�97����\'Z���81�������4}���[��bƽ'A�O`5�հ���d���������s�1}	5�R�s��LI�@��>k�&},�lF�?S��fV|����*�,[���+E{���'�����s�� 2��$���@`�k��MJ�#�K�_�2(�3-\�-Ҥ���x��e��4z�+�� ���N(���-2z4l��O�º�*�J��g2p��X��0��lYb�9� �ӌ���-�ŖvG�l�YC�#�(M�s}[����3���(��Ag
U�!�
����������*�ܪ/ �p��Iq�Ku\�.��1�v��,k������Y��q�0�"W���s��(���`¶h��č+��!y��)�LQ��2}+��( Z��'	����Ǥ�$�`�iF�L��?E"'�?K�ьfܡ�����Iv4^��D�w��L�3a5���&!�{C��U����f]
��/M��,Z^���,�'7~)��{��%��䃏�|��R��p��y�)�O��������e*��ѵ=t.��zfȍ�Y?�sDr�0��\��+{i�:zk�|w*�-�d�*��>���g�+�MW$x�B�aRTRl�K������#I�d��#<��f331H��.��\i�x[YYBU�oq� I�EnT���8�?}'tOT�0ҧ'�z�U���s]�j�s3�MO/J��l�߶��c{M�5d �VQ�SN	�qY΍2f��M$�u�o��q-�C�8=w�Z�m�*Gc�·��&�g�!��R�"N�������vDavS4"���iUL�*������� �Բ�_o�������"`�q#N���=�6���MB�v���ο��B�������n1�`i����~'�j���N�ϲqDS�i�G��om��2v�`��c�|�}�c�͉�De�mCL)�g�{��J��o%v�ċ��?����W{e��<��H|�z��������4���+ʖl�����Y���7��7��}���s��?]�b�?�"��s���|���bS�S�@���1ۓH�)�3ke��_�̪����:�֤'8>�F��O�6,��\|\V4�P� � <ww�@)� "�S���
OF"���6�<�q9��d���K(�J��m!G���=/}U�b� ��|������������j3G(�����=\�	صpq��7p�=hޫ��uyi��_�`����W>�E�2b�]YY�O�oi��N��Ƀ���!$A�|l�R"��$�۵�R$X�M)�%(��?�D>S!�!��`%uỏ!
	b�86.;s�@��I� Ij��r�������Gr�M1���y�*hj��n��1k]�bKH�Nw'΃/B�1C�]�̶wP�U��ך �/���L�<����+v��}F�����%�-@(|T�6���j�¤���b�M\�oc�R�L�H��o!*wE�՟M�!��k	LV���0Xo ��I�jY##f	�˖��+�P��.-M� �jM�^cN�����#k4�"1kq�� �;p�n�U�b���o>�6�r����<
�{�h�u����>;%�ذ��B��l��Mu@*��9xVG��^y��Cm��[축���'c��GD�v�S�`R|S�[d���وǴ�?*�6EK���|)����"��M�H!n|���|i��`����I���Ӿ�JԦ4D4��5&�zd5�>�|E輟"��c���"�IJm��Ui�ֲ�Ѳs��+�X�?��]�N��w��p&�eU:���/��Y�a�sl9�3X�3�B�dH�5bEUR��d�l�pk����:p���;kG�H����3�L$:�� �_��4��wlX��R��iEl�4,$�����]��ڵ:���^z_�����o��d���8������^��GLq��H���sQ�������L�}+�JkRK��V���<�,��z)*�Gb��zH��@��p����Uۮҥ����g��Z[�D�g����w|���eQ�iw����&���r�'y�D~��r���p$쎠���f.ԎD��`eH��?l��e>��/���>Q��l�	�^
�X�?�=�%/�D�&�n7�Ft�vB�?VwQݫ6u!4�>�����!����^�W\'�Al���o�~A�p���=)�ja�g�9fӑ4(�4@�D>���0�Y�d-�{�굡��e������P3�N�A����u�:��S�|I�KU��$KrS��I?�G�S�℔pp��-��׫TG�P�5^{pR��݃yf[�q/�U	s����?jaș6bD_Pyy���<��/kQ�X�!�t�P,Z�"�a gsfp8!Ӿk�����UC�@s 6(�䂂�v��g����"�v�.4��6De�D����I �i>��˻��X�+؃41؝����n��ps�B��v ��s���k$�l�R<�"��2��ڟ(����Ր?��]�E���V����r��} M����%�6dq�N;z��Z�M���c/Ԯ���k�&�0��x�	����?Z����2����M�>wi(�5D�n�������|�����1�`��?�)<%j�娆����lS&��e�bJ �tZ���'X�����I���~6+VG�Y��!����$�8�|�[��4L�*k��QB�~)s��>X3$��ϖ2������[-f$H��8�?AY���Žz{�u^1�؄;��U�H���qø!���t�t�B��mT*b�ChT���	;�`	�$0}/�:���5�=�U�S�g��,���n��!��r`c�*�Y2��K��:ж���X��� �rF��
TBbbZ��-�f�,�epP#bU�K��bO���?����#2�����ߥB����4
�L�JM�;t?R6�{�Q����@Ut�`D����;�\�R)���y>��"o⏘^GaD۶�\G�E�=j����Vfh��+��&P�F�{ػ�>.o[U�&���Uu�)c3�R�$
�Z�l���̱�[H'e�|� � *��-d���5���N��&���i)B\���jj(��l��~�.1�/2Toa����~/>���ό�  A�a�D|��#M��U��U^se��<�'� .\�����[5���6(��?Q�:���r��㭬��z���uSRn�+v����ٰZB�),还�_��+�V�fE�(��T�X��\1�vt���nCJ�ty�)�YMy����O��}��N��>o"1�3�
�0Ǐ�!����	Q5O���0c��$��cC�c���sL��x����'9\��#
��b#P�V^Y��A�X�����Z�`Eg�"[=:�M<+�#?����p�^�=�`���:\�[jXѣx�X�4��R6m��-��%�:�sEZ�}�(�(�D'�;eѮa�X�$ϟ�ĐSso&[y>j b���tY���=L[��, H��Z1�(��^lQQ��j~�Bf�z���ƻ�:��VC�Y��;/׎�h�/~d��7#��R���N.0' Y��V5��s�ZPl��uS����]�N�In�#�7��/\��H�6cV5Za����|N,lzVP�^�;�z1f<<=�S78�^�
-�?��3R�C;/�4�k� ��G��wHo�N�R6c��c�-A�@=�GY����F�~Ħ���@a����O�$9ȓ��J�C(3�W*`��%2Y��x_�G�Tl}��ɐ��E��^��˨V��Ȱa�9�B�U����'T����]�+�/�%�(y�cu1a���0
3m�V���`~2:��N��S���o�Yz��&���"�ȗ
��7*�'�Q��{
%o���	�G���ԥ��@X.����� �9mǘ儵{���`Q ��=A����u��ǖ��aoQ˾�~�לn���α�qjp���n�D��:�9�����3J�pX��_[)�kiL�.G��\&p�'�͌��Yx�<����6��|�&y }x�ɨY�e�0�<K�T����[ݼž�a�ml:,�pҍI_{k�I��#�6�P����a