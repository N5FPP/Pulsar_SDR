��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��e�ik3�������w$����g|��J^]�v�^�^�Ժ��|PV�����_jM�;�:�~�u�e�p{y��Jh m6Y��/��N��X!�4$��>�kZ��%hy:x����}Ƶ4�+;.X�����&5�)>,���\95���tlLc
���\��`��l��l�v�	I)�Q��-@��F�?��y|l �3�v�\D]�!}�C�@\?�>����ps2���x0tp"�	�*�]?�A�� `璏ÀfD��h:#�hE-�"al���3���������w��E�~JN;p�m9�qǭcddJ=�g��7�[ME�eeNڲT+�z�ݷt��h���s����B���'��b�I��	��z�#�d������a�yS%jX�q�z^"�F8) �Y�T�(w
�/E'����2�Q��C��R�z����7t;�)o����':J���7e�nV��|��#�����Š̰4�HaS|� O8	�Hy��Yr�Z����������T'v��MiF&n�rj2��/��sq&C3tfֺG�PA�C��!�Y ��#HSf��F 7hz�q.N@��1�S�0*MA�D����a�3'!�}G����1U��J�_�v	��-B�OrN�͹<'Ͷ�]�b�J��Hy�}�ι$�D� '5�����ڷ��Nn�Gr��j-�W%șiE{{�Mt���[��������c���ᔣ���]p C�1������)i5�/lok��OaG�MϊD���ןt�V�L����l� ��v�?�Љ��<e8��M�[�jԐ�������>�C��@tk'܋����5T��5I��GzGЯ��%'�T6�����dP�U�)zz󳦩t�����ݍ��Q���b���4Bn�x�^@���k���<CeK|)�P9���X8DW��$���?e��l��,�x���?	�!���3A8��]-�t��k��G�ұ~V����$���x��̽<�-	���˱���ď�O���x����~i�s�H�Q�ĠҢ�]�N������g�z�=E�$���i�S����g1�RC�w7�A���2@(�;����U�K�:u�:J� @�K_8��vqǏu�O3�NT<o�������C��Rp��D�5�)��z��;^������L*��N�� t�+E��y���ek�����V��|f幺,oH_�p�|/>�Ŏ��\y�2���\��r3)�\m2�S�fl�D��.\v�$4~����� ^U �����ft�Kp�4��Қ������'�*-h��05�o:��U��ԋ#��T�t��y�a����R���qe�2�7�� gex!��$������"�:�A���&�Ȗh�덋�����F컟jH"��;����tm�)�PLk�[���Iuk��Į���� �e�y�L^!�ñ�4 멟;��I�?� l�z�`��MU�>D�C�h&�H]���yK���}l��i>pO�(�!M�ڪJ�����oG��� <$3#����<$��2ͩ��:D�_}$��M|^$	�Z��kfO��iOT��p=�ÇТ�ȡ��J�ɬ��l$7�a#�2ox�?�y�֯�YR���c�6��J�nd"9�����B%b��H��i�.L��.@A�y�*�e���K���6�w����h�n�y�Z'��s�W,���X5w��z�`4����k� ��[@�_ b��Е=�u*����O4�������}{�ʺ/���x��~=3Ú~ܙ���ZC"� ��L���tP�6"��Zސ���P��L�0g�l�42��'zɂ��ӡ�0��pg&�'���rBY)(ѲW1���ٮ�B|�v5��sY�a��o���YV9�]�3��/�����ꆅ��_1��t��a�)Nc>��X���H��O�����[��UwMӢy��\��i3��o�q�IjzVIc2�Cr�`���=��X.?��%�Y��|\� �6<�+>�e�#�T�令=7ρ�A��?�l���<��ײ��Wŋ� aT7�3h!&I�Q��l|���J�l�h(������/�7wAGzz��o����B��|���`��9g�W�AQhL5��{�IJ?��fHo���[:ȁ(�?˾��3��
O��	�^�j6��d�ڣB�?�Q�h�wq0�_��T⻀zJ3F��l~$	#�l�aCG�[N��2 ��Xm
g��Df/��[|"�o|~�qP��o�	��"�y��x�$]�� Vh�M�g�e�m�}2.?���j~�A���(�q/������yw73-�F�ݏ�-0�`q������oNF�J����qk{�IeɞmT����'��q������(H
PK����ǈ:k���V�k��@:KV.��O_��>O������-��El	��3���*��6k�������̴ZQ�"\�1��X�O-cR�M&�I޲7/3D!��-,����-˽@�p����D����*�q`�o��iLun�|X�j��"dQ�l��e_?�GJb{�
����tlr�^�;��Λ��n]�a�/��<i�(�([lݎe�p$0l���epy�3�o�R6|H Й�1�WCwDfZ���m����B�S6i`�"���a�|���OCL`%8��I�v��Zx�X�K�ѾX(�ԍ`@@��:Y6ۜ��{�Ake� � ��I��V�d�/�Z�r����k.����L��`��\�BFY��S�a����O>�>"�J{9P�{���JX'��[�|����`G�|}_�9���I� q�U8{b6��ʌ�0O�Gq��}2�݇\����όĘ�уG+�v�g� '�L�]��3��+�s8f�]��W��
qQ�!]#t�ڒx�	�5f-.���~�2"��F<�ax)�/�8����:�R�]8X�\ݭ�n������$^�a���s�� Θm^�~����6���<ZC�"�n�[u��j�7}c�k�v#��Gڜ�F�mQ�T�oc3{w�΁M��V��x����0�H�]Z��ŋ��'��N(q��FiՖ��뜋�>£�A�%�~�\�:��a0�h��1`M	�& �7RV�+�� �#��*B)�"E�$���j��C�YB�7�~yޚ����?�u�d���U�r�u(��ݺ�"� zq���q�$�I���y>�.FP����J&ALR�XR"h�d&��5�?�]i|T��.$"�B��Tn7+�iM4�<�uK����P��3S
��\�c �*�/@�dې�Kּ�����Vˣ�S.��c�\t圯��4�`����L4��s���x������s Sdئ9k!�J-sJ��!�'�wkL=t�
�<�3V�d���*|�@����o{���o��h$.�4�ؽD�	��FJH����Zݪ�ם0�L�D�G�&vm1��Z��Hy"ďz?'۔C�15][��P+�gcP%����:"͡��#\�aLB��s���|i��`�,Y*����?�5$K:�G�^��9ITt-`�=:8��9l̃��;X ƿK�D�\0g �1�&b�m�HS���c&8�'�i�Ǚ2��ǻAm^-�4@��w�K�xp��<��фK/����l9+\��U������RG�vlǒJ��_�^%��3�Ô	�L��P���W�Vg�ǧ֤']GZ�q uV߼x۪��k'z$,9}1�N!�B�Z6�Q�V=`
P�[�1�24�Y|��B.J�sW���-&�biE��7�i�:����~����ѬS�S�-�̓'NA?�eԇY}e8��;ء�n�{*�~O�G�� �LX��,�w�u��m%�S��ə��xS}�(I��Ur���k��A,5ceP�:kh����<\�U���Ⱦ+(�o���|z
P�T�h=�0cg�CkzR��nŉ~�Y�?��U{�� ���u"�w�3Jj���0.E���\ι��v�Ҏ�� ��Pܬ��KP�����IW�V�bn=��[U���J�-	�~%]�s�Yzg<�uȳY�B�7#�̫�dZ�kZ���A;�}���7&�ѳ�f��mz9�0�";��0�CK��������С����>IKi9�:h�f�c\�<�HHW���m��=�&پ��}�:z��<���9��?�J� ݗ��J�	���E7z�Ki���9s�,�A&k��+�.�0h+e�2bm��ꨔ���՛KW ��ʯ���5����"�H7�<J�7�w�'��j�Y�Ȝ���T��d���U��t/oJ -�2�S;�׊'���9z�B�T��S���2� r���C-]� "�^���3���(9m�Vh����Fy]B���3>j�Z�5��%�����2��xL��?Kݺ�Y	yCᛚ��_q��u���s��'�[G�X��m���Gtc���]Ƭ4�mrS���	�� �}��^����4����A�&J�bV�j���u?~��A��ZR7>�p|����9Fԗ��ǽD*^�|3�8_�x�Gӽq�7x�|�����Y�7�[s~��)�Z�>*�2s�W��Cd�Tʟ 2:Vy-02E�0�C�3��ewp�cG\�d�MG�?c#�>����p�J��FМ��
Mj�$�Rσ��s�i)gUF�4�y��,e��L��B���@{G�_��[�'������^{�{a5{��h��wt�<��в�;�c}�td̩���qz�v�)��Z�>��Ⴝ)0+�A�! ���d1�!���7�&�	���-[���!oV�Q�l�b�奌��K�� W��霿a�urE�*��0>.���+	�Od�^Ǟ3�ic��8|'*o�L3U�RA�<&%��[k���M|S5��Wt��fԟ~������	���d��C�FX��z:)��~Ӣu��ul���d�C�F�t��um/IToyHl�Ӫ&vg����?0����'����b�BA-'G���E�o>�w,h7(��}���[)��c	^����ͪo����1O<=4	���������;Q�/��|:�5Ļ�� �_T�e�wyo~2?c�Y ��]��j��7����.{7K7NK���5Q�o�w�;ߺᎄj��_�r���3)��_s
���$��ʖb_.4Uܝ5��w8	28�A�>�m��;�D	'�uZY��wR�I]<�g�D��e甍2ё�Q��e��z0c�Bc�=�o�.Qisvp���L�[ ���dz� ,����Pc艼�0��0�=��Zd"��d�T��G�) h�L�C����1C��lwߙ�V�w�w�[�� �l#�#C�('F�$)7�8	:�o<�Ra��8#�Ѭ�$Աa|�7���R���y~jIC���	*�����\WEj��ܳ���+�| �5VE��G�Rf��J����}�^#��yi��Wg5^�'ˇ�G��CLū�%����.�W �	����=��d���6����I�'_B�A����Ǚ,zU�ة�h�)Jx��
D�)�D_��ޥz�םh�,BӖU��Ԛ��鑍��~�j9��I�G�1��]$��!�V�G!����[��ƨ�a�0�1��In�	lk��f����a�7�td1� a�h�~w֖-��|)m��\L��.+��eP��u���C����D"�F9��0�d�-���cO�6xH���շ���D�~�1���}�m��!�v��!m�E�����Ϩ���p�*��l�'���2��ib���14�	y�$�5�;K��e���P�7�����bF�����)�g����с��E7m��_~I�7 6<	�}L0��	=�p�=�<�=Hͳ(� ���U"�/�n$!�5��x��[T��ڀ~��X7�~��Íc^*y�`��Ě��1r�jUDI���T����:�H���0�)1a�d��;����6������b͡�����臗a-�X�9�YK���;�B҅���V�Ú˴��� _K���ڄ�f�E�P ���I�����m��D�z���}�a�k����
cd/��4����/jUH�4�EzE�Tc����TAC��ۗz���̑[�8��;��;:y{�G�?�|(�إ��S�Y_J\�p�7�