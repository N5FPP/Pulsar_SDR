��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5j jQ+���t��-�/����u��̩�Xc��R>G��$b�xA�Fn�z�F�X�Ӊ��q	U�z�qG��f;���,-vl��� 'J:>�V�	��0�7"�%�˝էo%���7J(]�7(MGw�rL�R���<c{��y�y$+{���k��6J?����ye�@��\��q3�!6���J�9�I�ʋ����K�e��t�f(��oǎqz':ݶ32/�.��.N�
s)��9�<�2�B�	>?�����V���c�Kz6]��0;YTHܧp��VS���J�0�L���<�0�q�j��`��Ѕn��-޾�Q7�z��׿�<SP_b�
teuϋ$y}�U��4h!���'N����F*9� z�[�����B�'6$���111��>x/�mD����_�X�5"���B��h�`�I"+F�8 3��R�f����<+:�5����]�-T̖�ߒ"���|�S����'l��]{�`!�к���7��*֨h��3��9v�w�'F��	�;����=6E�EfW"�UB�t ����Å��KKY��Q�&�5�c�Dv��7X��񋕲	+y��h�< a�D��Y?/��Mio��dX��vz��{[�BJ��?qq�:۟�hF���X<�:��/��|�5�9�_�'��0H#��丯����Ҭ���@z��JwHy���F ;��ʻ��ÛV���Q���>��{y5H����z;���Ǳ-�a��!��m�V��Q�J:p% ��[}���*�ֵr�P��ݯD�/�Q���>���ʜąïI�MH��V�"�HMf��$�o��c�AUl��K^�!�p96;�����Y"���p���_�a^!�M-'W�[�r���pU�w�i�)G��mr���l�����Ə�?��X8a�o$�P��L���'���_�H�4�>p���-�ޛ����Xyw'�(�ha���7��j�4��<W\���d�������B�?����jokR�'��t�Id�]�l.����3��K����&@��$ҍ���u�
 r32)-�6>�g����i��b�ҩ��u����H�}��Q��b]:ɓ�)֗��A��?"*P�	��,@�)=���Q���|NEQ2�����
qT%tR��5��7ё�ӝ���������/^�޿$_��_�d���Mq��(�=�w��=��츔{}�|}+5K���W�;�.<'VV�cL(k4��_�#��B����_P���Ч�^�x��=��Bo��T%�T�-�I�6\!.��:�P��UCT� �sə��, �ٶ[�hko���l��;Be�ZWg#�/q��,u�f��/pn�.�T�Ru�XS��-Z�hW(ڝP�LU���g�K�@���n�jWh�d�q�Y�!D?���"Dao�~Dhצ��xKt[��%��-4Ԏ�5����0�8�/(�9��ZҶy��	i��nu��[�a\	&Y�e���uҎ��{@��.y�7=0\B�M||�6��Z�G�W�3]a�^�P��1�����0A�2�r�u��y>�%��Q��z���zGhmG�'������ilŇ�CU>�v�>���_YK�:qw�+�z���P/rw���+ٹ��XQ~!��5��򂗢�n����B5G.��u(L��pU,-;y����"��yj����	�念O�����4g�7��`t i{�A+��!7���)���Je|N�������I��$�
�Se��M�l^�,h�K�0���}Z��ݨ��a���:Ci���Z�Znu^p�h]�ö���k�)P C�f�T՛�M�OI:;�#}_?nZK!�U!�����1�8�K��gik��6�dZ�	�����S�5��K�Q�)�v�`���!+@g�_�MK
�v��Q��+A�Pd�'7Y3Q/�eh��'q{x��%U���1�]���Ϣ��P�J����l��
2�A�P���5�R*�Q�0NڝI:"L��W�������ۏ�,>����=~��3��k��.U�
���}�[��V����}8ʰ�fޮ&aćޢd,z�߆f�瓅	��s���6
��hP}�^��ۏ�_djh�]���IB���lT	NB���L��|;K@
�]A�iJL���L]�@��5_�ʱ�,N�r;��K%��y���u����V���+���F'����.�^u~3�ɢN���^h�h����j��)�XNN�xB} k��(;MW8[��ѧj;�,����{A�q��@~S�B�,r��� �� �F0�{�gLWg2����V�-<�fvt�{$$uR$���+����4��t�s��QL��l&�ׇ���ڲ�����ˉƀ5j9"n��d�*&z��7�j���>\9�@��Yo��+E-����h�
V%��	����vϲ��H7�{F����W2)�'N�w#�A�����9k��bA������������s|?����F\.Y[��,�/��H�7�SǍ����E�\��ޫ���L~�����+���p�,��.lgT�틼S�eѾI^����a'�5��h�O�:3�'~�et��-0���b{������ݗ\l�D�W�mZ}��EP6o&��3w��x�!b�,)�iuf��C[&������[ҽΌ~�H�����?X�p����q��
�0z�".�n�BRx�k׻#�zrɺX�.}Mԧɜ�r
_��Q�y�6��M�m�(�hձ��,�#���@�o�=����{��c��N ��FT�؋�m5����^�o<N�mKlMH�������*�x��|rD��SL��;����6���2��Tj5�(YeXn)�u;xH�3a҄)�"�BE�/��������Ad�w;<�y{W�)|��Շ��P�F�|�1c��7�ȟ�x"���B����������/6��_nA"@!�)���_�������l=����\v$��n���8�U��tESY��.$Kl��|"��"�KZ+����xl���s/�et?@eG�zl)�P[_�	i��i�Vt?W���U=�H�B��(ȧ��!��W�<k#t|��7�l)l\e���s�`T�6�+mZV��(&�^SjB��%>�νN^2r�I�r��{]���W>����Z�e��͖���@#�5Q�K��?�S�����s��UC޵���Kz�l�b�q�z�r��@�$ܨ;a�c��:�(�'�\�K �]�a�3�6!�D`��t�xf�	�'=������m��/�p��� ��0ٽ�����R0���&��A$N��x۽�g��%%�^�_���0��E�*+��Ձ�Ϻ���a�	�X+���z��6~�!y�I'HP�k&̮mՕ(���k����-��1���5��5E��|�����`��j^P�9��3J�2ա�<�A��%�ie\yႏ5��Q���PY!�cX��0�9h""Ò�\!�;q/������p53vG䕨W���e~�S�K̮۬��2�c������K�����������ž�Ay���ɄE�:��8�WA��F5��%��{�u7Ş�ԏK�6E�j���ì^ĞJ��᥷dWcN fN	B�m����㏡䀬�<��+7�$H�-�O:�ԃ2+z�/�1F����1��i���)&�P���!�[s:4�����"4�D:�6�o|8��~�m�k[��J��#%�؊x7���mF�%�'?i�㥼)�e1�'�G�S�͚B��q�`&P��09���rk�����l���~�bp��L�"�U#'v���l��_�Us�OU�F��j%���e�n�V���O��v:M�����g����5in�����j�j��i�O�z��i��K�&�]�υ���ǈ�A������H�_��E��P�_fn��f������p�c��DV���z��砟aޯԷ`��ꜟ��p�ː"���{fx��7���������(�S��;�hϬ]gu8|N�z'�#�̜}��X�i�ޠ�sj�zF��c��e�t�XtL�40Dg�����#o+Y��{�J2��$Iy���tx#`���2a�$����=X2�������TR;�kR#����W3�TH�^s@�I�E�8@��^��n�r�b.t�ǠM�x�J��^xn�Onς�
�T�R��c:��H�9�ϯw�Y����������Q�Z���of���".vdT�2