��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��e�ik3�������w$����g|��J^]�,^R2�D��p}��"�o���$���8����	+*+(�`�ї����GOgu��	������< x{����8�L�=,5��}�1��(΢b�7Gs%�~����ޘTs��	��hÁ=�ms.3������NL��5�ճ�^�k�/���@F���MՒ�<�(;�{����++XQ��� ɧ���\H��F=�i�u���p�Uz���Ӕ�l�H���iYG�	�`ss�O0�>}QsE���>!EG�2�1��to��ei�k�i�LI����g)���Jg��<l�@[�;^N���l��5�	�5��wiisߋ�V�}A-���jA� 4��#���U�W���tW��� �-O��,�<��]��.&��l<�m� ё��Y���@��O��ӷ�W"�v���|��2QS㸳���Ĉ껔���X��o�阜����Lcv�=���9���J)RGspC�J�˨yM�ٯ���!���)�\��{?���­Sl�웠M�u��Rg�KD�sws_F/���>�������ò0��~ivӪvjk��������#K5�I"�	�C"	7w�ci�v��ʁ ��X7�N��˼�Wۛ1*l%4����B�+�8U��Y5A��jb�u2P�g��0�����������A��Y��A}����	QP&���ɝ�S,,ը�&��"����A+9~'Nón�E�SN$�F���Ȱ^LHA�ޜ��ܖsIR%�{�l��r's�ƛ���-&�����鈪��{5@�8i@����䌜A? �,��;��i����r���W+��zx��o.SKI�Jzm���@���6�`T��|"�JΧ������N��W��R'��dM��᝹~�O��q��*�M��n.�����������|
3�����\�?H&;�O[;���Zl����I�y~��0^r��'������Xk���j���œ]Ӥ��&����e�����ӊ����Ʉs����i�c;�����H[�luih�:�[���}L���C3��� rH�����Z��z�E�\M���k�4
������w����c�ف����*Xa��Cm+˟>�/%��� 7�͓1ܫز�y���dV�D�X��rp�h���\�Nn�H�,�9X��9
��/:�?c�HYm�m�E	E��3-�HqJ��QbI �
�ć7'b�ɒ�&pB��,�?�P5�
���[�pD6�,F,(�r���;��?Qy�Z~������̔�d�B]p�*m�Pp��+�x�-W��!Z��I?��}y f�zʬ��)o{b�9��Xh��oE�@'I���_�(tȜh}�m�9^}�s ���|f���۰V3�X�x�ZƲ�9[���`|�*!�W���
!���8�te%{�t1�x>���	�M1e�X�S���:�zw'!�*(�"�t��6�Q���Q�D������*�Qh"H�Q��;��Q�2L�����X�B�%+7o	�ߤT��Y���a�|�I�8J�He����	(sr��no���S����$<�������Q����Y�y-�%��2�K-�~���pV��mLO�@��S`�&�:Fq��_]�PکV,0��S��K҃O��m)h��A��wm43Cԁf�Sgo��1�Ρ�����I\�O��R�6Se�~> |�����0k0��`����NǷ
T3'.9��eK֐����,A
�Y6Ƚ���xvR��L�o�4������n^�*�/;���K�k�)�	^���H��^�ȢE2!��G?F=l ���`ukK
�m��h)P��uA�����:�
�@�V͊ӭ$LF�l��;ҳ/����y�_˛B-�hggV��(���"`�v˱y�~}r,�-KxM�f~�Ϙ��|�P�6 ^��JH�Y�Nw&�ƻޢ&@�ȼ��B�/H�v��s������x��7`ɷWP55��`��T:,�����a*�be]Y��j��� O~����\����Tx��Z��|��Z�	�k6��JC	e�KGaَ	=��q�+�_g��eʳ�T�oDg��#����.S޻݉t�߅��%�8�Xl�BV��d� ��_�W
;|d�҇][X����|��J��a�5$��d*4P�ׯ��Ҵ9K�V<
Z������·!�-:n<����z�3og>���ϷGmw��Mm띮�.����\�Mkt�3�.U�H6oݵ4�F]qy���lo&6	(�K�8z�/[�ccˠT��~@�9y"�jڄ��sv�z-�|Y�Y×ރ$D���N�	���t��3II�)��e�J�ٍ����?#"�
�y�24��k�%�ҩ0*R�c2-� ��"5KV�d��^�ݼ���axɴb�,οY�R�����%e�I����j.�5 �<VO�1�����_��]R����@'����{�pHZ5�)�g|���G��	�'t!�Z7�$T$�
4�|5ڥ�l���R-�dm��=�MB��,�"�y�3`�w���h��)�x��{���j�TF-�x7�hͥ�N0v�V��M���}��\���YR.g	`2X��ǈ��w�i�,�^����ƣ?��d�~.J�D��f���T.�>m{��8
���Ń.`�����/���T�Һ���-�"d�X�̍,�(i�x�l\YF�\�}8O�k�Zi/�~B�tK�`�3
bi�[N�����N��]즿?�D��t�����NW�������-4,١R�ibA���F���*&-���6�*d*���˫*�o���>?��ӌ�Xz{�|y�ᾌS(�X�h D�&���SD��iKlK��To28�'�"�Vfd��G;�u�F��_��61q<��kޘ���F׉�h�OҥJgq;YI5~4�Dq�ϝ���鲰���1�K)����W �q��ى��KqJ%a,b�����$Pk����h�i�`A$a��B$�g�� ,�/�I�N�-��Y�U�U҂8�2]�u���ʢ����h3&��f<@����9�t|N��"��5����Ub��G�b���3������:� =�;N�z6�x�ׄT7��EGD��QA�*(�W��R�ٻʡ�YDj�5��uj�>�1�Z�D��^"�� �a�L�;���_j�W$C��R���'Ŷ�E�FJl�m�T��Y߀��6��!E�Wr�u; ��?ë����b|^����6�"�8"?L�A��h�#��(=���5V���K���Q�*��!7%mPB��gGK6+�uy��?��o�O�$��۸"�2���:q�c[�������k���X$#�"�2Q�h�5��7�5�%��Y$��d0�R�f�I�:�J8H�w#����H���tz�����4���X��+��N�?�g�Sq�	�w>��ܒ�CnXY5w\�Y���b������[��(�$�<3�@�7/�����U�>�ϋҦ#B��f���;�x�ˇT�q��8/S�_yh-|a�u�����O�EHU W���8&6�TA��u��U�R��9���t��.��%㵅)9X9o����Z�gmQ䭃��K畏%	���uU��
��D���r���陘�dZ�
t��O*t��g1���
����s;d���,��t0��W3��j���S�Aѭ�V��G��6⃷�mB$��2(�����of{���?!�Ҙm�N�ˢu*+���G��7�H�A^�51��xq]֛km����ߑ�q��),y�U�v߾����im|�v����N����V��?�m��d,�uȻ,�!��¡*�� hl#X7ykj
Pu����C'sC�Z��5Dar��E��ܻ8�.'aB�׍�
����]�l�����ה����"Z��Z�0{����g�fX=����ߺ�@��*���M���IV ����o�ue��n�a\�_p��I�-Ӆ���tl�*�����A�UWL������WS�o�յ�&���=�����>=��Ӻ�u7������R���]�u �/��W2U:��OC%�rNʩ������ͩnZӎ�'����b0�g�^"��?[Y�.(/�F`(�o�>3y��0ba[]�;�����t������p��7U�_���r��,^ZE=��,���"�Ǻ�ŏX��ɳ6����)d��N7�/���Y�����`���QK��P�i���U��g�NA?����p�c
z%'��Nl����CS�j�����|�U�#?���u�{EoV������)ۮ0������_�c��������^���I��/���<g��D�ٿo$G�@p{��CZ�)P�9>��Y�+<�y�H뫏Yu�	:q����-o�.���ߍ×WY���0��y��^i-^��3}wA���n��aQ���g!I)���;�h (Wܵ\>%N8��"\L��^��_r�+�	`�����VH�ϵz�n�?_$"��|@�(~�� ��E/��QQ"��xz{���7=��L�~	Y�Y%.	�����&�_:�q�!�P��>F<P2��櫜�:װ����������'k�s�
\�T� ��(����z�X��{�����KK��kIV¿h���A��z������8'�:�<&ٙ�p��u9r/T��!��]�$fn�u�����D�ST�U,�j�&�_0�+��a?�Ɇ�7��iF�P�p&�:�ʒ����D��Nh�aӳ�u�p[�]ն2צf�8��'�sҖbjM��;�g���%t���2� ����sŗ����<�>�B%�zT~�7Xk+����4��t�\�a��°���$j;���͍�B����P��}�_ܩ���[��V����q�xӪ��f=c(�4�˺3�o=�6K��K�.�� Z��~�U�B��v&2b�/4���ӹ)E�ˣvʝ�ߌ�q����W�I}��c,v0�F�(<��F0�}�f$F��XA4�^2Ü��(���}r��l�a+����$__���>��O�N-Z\["��UpB��q����)p*C�"�W!�M��F?O\��i�و��ޥ����v�S�Z�� �ʗWjşw�+�U�9`��:�b1�2�-�!��X3�%��r�D�H�3�l�gS�%����o_��QSH͟$>��>�BbkwN5��H���l���@:nL"��ת���/}x�|��{W^K���3u��K^�Z���z��~��U���YX�<��D�W��f�c��Z �7r"(��@����5%� E�6AW�_
S��i���֑t��=�%�͝�gר�~j�f�T	Ў56)ק]��:������)�������%���.���Sc�a��P�Șç5�72u�.��AY���/l,� \#U!wSGfμ'��{RH��Y�K�-"2Fy�:J�x/��+�P�ة��c%�8_r7Ab	�>?����?r7��X�E��Sq��b:�� *쟤f&2�� �AtB��%�RS@�P�+&S[k���B΃�HNގ7�z�j��wL�ctB[
X*I|~w*�X�:�9>�E���(q~�h�p�4t��Cc!0Xn�tW����.Xz#Y�D�2��ߡ���3�!]�����mjj��<���(4�JW�n`Gj��\���3���<��ߦі��BZ`�U�(��/�@b>�y8���𗁷
�Al1G���J/�:*�[?/fl���X_Zt@�D��#�� � �W*(�
�~���Q��D��I�D"��"o�2�^���nz�68au��F��
*A���鮐���E٪-�-�އ���!<P�z�S�O�+;�^d��s� .�u�
�Tq|���8�]��#\��{vC�k�r9�H���}}�|?I짷�	d��3�N�ż�[�x��hI����^���J��%��oYL��q)ܞ��_62n�~uO�([=O)�ѳ�ܜ��?Z�x�b�#�'�sM`0�:Ӹ[!��D�������t�'N@Qc\@w�OL�$�>�ȿ��Q����B�X'��0�3~N|"Jo��I�;���`iڤu�*P�¥��3w�!u��!`8���g��cok�jծ�������b4���'(3_�r�I9�lB���\��E|h�K2P�+L,ɑ�����f��nF"zc+7�l��uU��!�9�����ӹ�m��A>�_�CV6��SؼpW��Y��bV3_�]2���������u��N�n��JR�P�����5'}�}�d���*:)qmT�@�0�N�/J����~�2�2�,,!"��T�&.���ucx����K6�}������{W	�*�ok����ͬl�*d�u��*�n�Z�j5+�X �ڄ�I!�0��������ف��9-���T��������(��Ӱ!�W|��zJR����/ ����y2���`��xuɒF\��/69,� �2�#���ֳ��6޸�_l������S�~b!C�W���ʸSeޒ���8���>V)s��-��E����4���:-�l����y�~���&&�������҉�'�����?��0s�vTT���d��q�b�Z{K�L3`����<��K���k��(�Z����H^�טh�4���� �+��a�S���u��@�6�ccP�W��T-�X�uք�W6A���T�����o(SS��Q�<Mo���n�/7\�3+l5&�����j�+rd�n�h����L�폾�������mZM8�b��� bO�y�;�Vp���C(\����_�lhw�7t��F�z��|�^O#0R=4?6���߹C��P��3B���/E�dh�h�r�| ����A�fiy=1m^����x��G�E'F#�ہa3�{�+��lض���#�I��_I���p��`�3HB�m�@��b�O�g�˩�uJ�٠M݂����@�zě�c	���v����N(g����{T4�#���0�����%&�1���MQ!���d��c�<���)�Ca3�ܖX<�c�\L��]lmY0i�{sf|�e�o�R�6i�Jr� ��tE��4�Ԫnt�ki�	*����B`��J͘.�
qw�×��:��Rn�荫�Py�(���{Vu%�S�J�P3��f���"����2u�b)��z��1�5�;���8/�ԫ�~W�(��s�z
�!`�7=ˆ��B���m��[5��Jh�	ı�24�Cj�}��I��T�J��쪡+�~"���!#�����D���@���j�o[%�?ը5;�ǁ���gN��<*�o�I�b���J���O6��V&�ad �涑�ID���/);�n���J���'/hA��VO�߹�\��/pJ��֜�kک�]�e�.��{�S�^`����D��r~2����4��Մ�5S��-p�"I$��!�2x�T
|{����`5+�Lu�B�l����΢���g/)f�`m9��6����Írr�hMC��[�H�XȈ%A~"�+�� TK��|�/�Lv��C�t��}���6��#�[#A V���`ٸ�N�YO�b���(������|����\����B�ܲ6��2BZ�juT�݈���+,��\��\ͽ[�.���w��U۵U��q���6�6�3������B��G�d-���0 �7��\�]=�4�S6��*C�
�qs{+�|��
<`�+�����I6禝��uy�~��5�$����䖘�2qY�˒r�ŶT�> �_��L�=���}W�b�.�'7ë�lV^d�%���d
��� �4�D�nX�
��k"�^�5a�1ʝ8�A��Y^�S��N�)N���بR�s����{V$u��`��X�P`���)��;��b�lz\֕� O]��i�i0�b{D8 �D��sǑ�T��)���DT�Q5��v�Z�!ŀt�d9ݩ����l5-Sʞ�cH��J�>F4t�F���H��lZ}�+ /����s�`�ս�3A�Z'�Kv�k�2|��{{Mx5eːio����A����������?$���Ǖ����*�#�D̎�)���Pp��B}W6�z1f
wXO�l�ĭ �<C����߻���h�@��g����F�9��H
�x\8�Q-���L�jO���D�\��?E�3&Ж CQ������g�-
P�VP�����gAj�4�ݲ+�.�Y$�����`�7W���.��f�|��bJ��n6?|�Q̡,c�;��8�l��=�I�G3��Y,��4��J	'9���+����t���$�۫X��8Gd�vA���/&�vF��z�+x�5kD.�_PːЇ��S�$ѫ�+������G=UD�2<-�qN�*R�IO)R2DuMNmPx�0Zot��E47d��!��^<r�� 9�Q�8��@��6�ŧF=�~0��$��98��4>~lqh9I���W�4>�� Io�� ��� Gm�2<��as����a:N��?Q~��E�A�ʡ�	s��ʀ�J�4�B���{�'NB,a8�����Εq�<�굳;�M�7��R 1����5 ���S�xF�m#���t�y�we��,�ßx�ۍ)�^K� >�Hn���{:,T��(���@��9ǚ��N�U����T`��.)�����Ȍ��a��6��3G�3z��Dd��j��t1�����W;w�obK����H���޻M�����H�
���{��+$�,�I���;����b��ԓ^��x�:~���`�B-&�^&�
J��hÚ��!��L�����ffa�xL5����E-Nߎ���b���o
O7z�e�ri���Bc�l���E _dF��1	ռ�(^7ʅ�O(o!�!��Zt�
F�r5y�vUr��@J:�p+|�+���2cЭ	�+�HHn9��=�yw��q�ג�$�a��9�D]dϋ�>�ஹ�U���y޹�0C����� v�=��tF�N���A��4ͨ��>:lHqk�]����{�Ԟ�v�I-_�|���L�n��w#�$	�oO[����5�dL���	��.�,�<��2��J����Q�$�.�;Ӌ���_���߸���B���$��̤���@���t��ʠJ<���Glw���~ܓ�M��Skr��=�d5j�!D�/��n�+Fn����ӛs�ĚF��x�p��ʊ瀅�T|K���{0��}k�o�[���,#���!�n�� ��к�J���[	��z�R'"�����g�y����fzϪ�
�$���X�Y:2�^�޳]1�"6����'�b��[f�����ME�'|\7a'c��AՊ2��9����W���W��|?�z����C I�+%i�\�2M�=3(*�<��U��IhSPT6��q��1}/Y��&x�]W�L��|�����Ż��xt��`N��}�t��U�`�TKL���Kq_n�d�I^�Bf���e�;p�Z��?yW�&�[H j�(`H�B@�I���&��h�:o��Rq�z� �^���b����t%����x���@�(O�&ot��p�rn��Z���cLo��J�*6	�����\>�('SI��A���]�*SW�W%"Fϛ�K(d��.�t�&�/Ɠh��o�t�֑ګN#a��?9��I5F�}Fρ�7ZW�e�,�W�cO����Mђ�P�6P>kJ�dD��$'q��>�����A�\&<� +E-n��nM��G#�s�y�')��*U�@ �s
=gQ�A��"h�E��`B���uG2y�)�|4,��.��ڶ>��{��ܬ�CP������`�"�C�i����a�?q�+�xg.+Tj!ƧyR �	���n�K*v�s�'̕;\� ��`�㶞-	�TW;�����G��5٥}F�$Q����ͼ3Nm0�b�7B]� sW�f�������~�CUI�{�'ӈ{u��Qz(Rۨ������dP~���A��Î$��[D��a6��^����Ή�)�y�[��A�Ӹ�|f�����&q�Z6:^�n�p��]8;Z�(
/j����W�_����'O�Htr��8�I�]���#c����a���o&��P:�P$ת����y�f���A��1��+��%eӉ�u�+�<
�����ӝѰ��n��0��2�KH>2�N�!8a<��CoavA� ��i�f�C_)B�8�t�9XQݨJ�T�öT}��"!�ؼ�u�I��Gk-Xw~0݆MJ�7��z,)5�m�'�@r���K,�㜁��dޅ7v�!�����9_�e����By�-/��JK/˰4��c@���c�v�ܾg�!O�Оq�$�t#p瑍�$:s���R➺��s§�
��.��\�3�� 8�ҠsFs��}���Z)Tk��t�?~����#5��H�AE����
�N�hq/s1��Zisq"��N�Y���]����9�;c��P�N~Y��C�ɜ�Y&/ 	��!�E5p�O%�W�o:_�#z�s{ˬۙ3Q���V]�[�N������n&�� |�M���C�f���P����_}8�:�QV/:\(e��DM�~B�'d�\�uU���Ǡv�h*�`nsޅ�@�L1��{DZh��t�ex��Y�T�S^���������]���GST���.����$���	눙��z���JMА��)�������P�i�{�l^i���\�h��dj)(�:ШNk��@�5�������s�>�DVL�ڸ�$3T|�j��.Þf~h(?w�ة_������j�[��6�h2�&'{����-�7~�\�d��5�q�&>�G�B(r�@���	=�nl$D ��_��MЫ.�*�;"�<v��^�iA;��N�D��%r����󱊰����}�]WDЌ�i�
�?�,M�ڞ�OՆ`�;LRB'�O��C-a��@���58v���r�gα�����}�v������7�0d��n��@���t�������~}j|����79���IKfm���`R�+�+k���͛�#y��2�KN)ݎl�+~���!�F�~�C����ņ��`���Z4gb��7ng
���Ԯw��\�	�o��,8&���4�O2ط]�#s���tS�.p�bE^)�)ɛ˗21R������q�MU L�v@�D�(��`9�-��-�0E,K�oGN4S}gu]�\$=By���v6ď�I$I�臞����{ꖭ�?��z=���LUS0�zp�����Y'
�ŚV�"̰j936U18�i������5����ز'�2$Z�o��9�Z����E�5�є��l����ѵ�����Raܡl�x���S�ȅ+_�2��W9�\����'���[f?ͮ�0�K����.9'�mZ�M�8}kaGk �:��Zpo�E>��*5�j
aP
 �WP�Ȟ�$����oJ�m�s��S^�8�9ٚ���ru�՚N9c��z���	�1�O�T�lg�rW>�z�$�����Н�P
Le���I�܌�3)�� %D�"���C{*Ě���Z�sn�8�F��Z�J5��A�l`D���ʟ76�SӗlG�gFPu#o�Ju�&�����Ûiz���W�R_�8���1L�&�/E�k捸����X�KLL�$T�����hT+]�a4�:C�m��2����x�2�ܱ>҇���~m���C����y};D���C���E�2�(>��EFq_WE��wn�����v�?�!�K������'��}���h���,v�H QlA� D�X<Q��N�R7lgB���hz>2�J�Ţ�c5D|�5%����V����Q��(/�qw�u`��M�v�L�?���]�J�
�������j֛+0A��t�Qw���
�C�[c*�i]����Nz��m�l�N��&� mi�@f�m�X7�E �R�����J�����d,�y��wv�8m�c�_JG~<y�ɩO�|ծ���$U��q��qk(=x�kZ���?"�CR�Ǿ>8�'�+�]�6.�XXO��F[��0�U���"����Tw�>o��},�ɶ�<�V����\�g�é� ���zU�?�����w����� ���JU�����51���[;rS�5���lv�>���X^�\�h(�_�9��7�DSiy�^j�j�2O���-���^��E�v�ׂ�4��_�!�my?�7[T1�^����*[��t���B��D�D�S�\$X!J�nϛ�ltx�7Ғ��v�$�3&���똽���$;���=�}��f�X!��w;���5`3Ő�a�/�b�f��9�z��vD�Pȯ�ڜRF�%�
���l���:�D�:5�2�)��&���r�����΂��K
�rhL ������@�QB���Imp��meN�'3����o��x*d�TIGXe��2a� c�jԱ���֧�8�u�`*}��r]��K�	�$�5[~L�q��]����w�����iv$-�:�L�0�W'6���&�����q(�
��P�\d�B��KAް&g��2[%ˁ�[:x���M�_e��xu�u��?�ْ�B�\b�>O�_�sƮ��턯�Z��K@j��HF���/R�0����0�D!�ujg�6���f���^�z�@�/�/�w0ưK�>���׌+����1�.��Q��ۉI :R;`
�P&i����ra�.���$X�1�o��1�ь�����<��-��G�ۤ K0���񂞸�T[�BF.y���ͶZ�ƈ�֢�L	P�������Ỵ�G]�y���ē*��m�Nlg0�����`��; .�Yo�֓n��Ӂ��`��nz�jR��s���b����ȟ���ɽ�x��i�+�TᶧO���7T7a�~��u���J� !������<���ϩ"�����X�0�)N����Q�H	[�	��vY���(��ĵ�6�Op�Vj�8Zj���"n�I�U�vi%�5��I��N����`F/M��s�T
nlh���3�ɽ@���,ǡ����Z���7�E3�f?"��0T���n(�as�4EGq6c�����o;��ԥ5�Ƭ������R��%}R�K�\r{�)�Q�]�^�cp��d|zWE^����kt6�Y��%Cؿ��s9�SYY`q+��@ �V=3��F����Ly��<���H7KrR��9�jk��?cl˚K,�^��0=2s������fW�qڦ2_�U���~Q(�&vu�훰7Y+sۯ��4��m�Ma�m�m��&;{Ԛ���|O���!偽�]�o�s�=Z�Y#�54������d�N��$���D���<�'"O����֩W�SF����f'�J#����i=����13&P@G��c���-�`8��^�h���/����<��p�iX�3�N����Td0^l5JcY!���(�����&9��=%����ض�@�W�f,؏�dB�	Ɲ�o]��WOb�u�*���9i t�������7s^j���{�n)(��2g�F�z<���8.�_���$��ъMT�mr��,1���{�8�4[�&����� {�2���
t.$~��Y��O6�qŅ��Y�O�df/��|�9�����	��H�G�;B�	�2���v=l�o{fȻy����H?�]��� ��|�l���H3|=�
��H���z*`y&IP$�����IZ����ݺ��>��%�4~5;��w�Ck��F�G��=�_ϕң��p��Їs�E�h�8�����qPWΝ뭫�d%� %�oP�C;��@�0Vl�'ӡ�X�3H�d���3�q�Ƣ����棟����57�h�\L"������l��?��N}�"���P=D��N��?��_.���V���0W(�rh��2l_�`.D����y[k��EL4/����{!�ar��}$r�6��|5�M�e�Q	�#��׻T1�x������{���Z�~���б/,�3 �/�5{�H�½�j�d��Ae�Ɛ��d�����G�#&�`3i����Z7��!�@�0�l�Xy�֍|���j�Ѩ�p,A)	<}�.c��b &�D ��8�e�o�3H��>UL�*�7s�Ҍe4��&ʉ�h^�a����R�5�z\�*	�A����^�����x��7���fcG2dD��|�SOk��tmz�=�A�n�:0r���nKS�\m�sY�c�?;�?��u��/��`Z�ꑆ��7����m���t�T���srD���SA�y�we���'��C���&�]��&; k��G��2h�q���G���T�?GĴ'd����hn�
��h�j/h\伨�{'Wn�H�;�:Z������Y<�KǾGj����X�	;��`�"�7��2�jm�P�h'��
�/�vc�a{�!N�P���B�n���Ƭ&]�!L�z�Te���n4�p�9���ܐ����$f���o�I'�P�Y�����y��H�i��ɮ�L6g�т �1�>أ��S'-Y�����.��#�iy�_�;O���vI៟eɧ�[����d�HoΔ�t4�����\?4��,��/���m��[� )+T\��7�jM�����͑����?��)%���V[����m-�ak���&��Y�݊0��K@!ύ�
Y�UVE`�����q����?
J�3���
���A��*��j��2�����f
es#b��.�~�m7-��/	�GM�^��zJ�R� 7/G����S�w�.F�:ZCݚ��+��v�U������>��Z�{�5R�4����S	.�Aͮ)C������^EIi>&�8��&Rp62j�u��%_������%M��>%���z���H���2�n�o� �����92p$W��ꪜ�Lt��C1zJ/�_�Б,���� ~�K@�?�m+d���87$@��!���8B�n{)2±}+�!�.@��_e{��������?��bM!��41 ��6؀�c}6FRs[x���
mn��m��(+/�ԸGq�l3(��+��Qa��}k�qK`�M���_���jמ��:����JՊ�A�� qi�Z?}��m7���=A�ؤPr��h.�nҗA��F���^��d��yo̢�3aK12)�lj�7H@	����Ĺ�i���M[{[�rXa���zܕ�i�Mn:vmu��������Z�MD�5c�m_u����e�Α�+��ħOs�)�XZ|9BR$��Y�����k��Ů-n��,TH?-�8�q�ǒ,�B����)z�o�$����Di������N6�hnJހ��(�_�tIyS��[�+F����bd�B���I#[���t�.-V<�M��Q�X.wϰNPY�� ԏk��煮��HX�5Z�S�[wU�).�-Ʊ�$��.�<���]�����m�p��-5��шC���3&�k��s����J#�b��C�9�͝�S\�Ậ5P4 �O��+�!��tR�$&�%p�����[�F"����߆�l�;\;K�3!r�����&0�5(_�˶c�Ip�WӶ,�Ϡ����TBgD���kC��[��O��H����W?�g�Pf���U4U2>���n�ǲ��Q�b��%��kz�1��橢�2��DҶᾟ�l�Q�#I
���Vy���5J�ɚ
��\B�H+U�/11r9�am��qX≺Y��y�vY@�,���4�a��z���?Ēd!D�*��}r�
�g�b������:�2����B�`��� ��4
��!ⅱ����'wx�C��A@
�(��ǫ/ƅH�������9l%���+�l��&�Շ��m�W�(��5呟@�[K<��r{���+�� ۡ�f,�����-�b��*���P|�p�@�;�Y��1gxiy��R�l�[�Z�y�x�c��o�(�;֮;�6|	A�ԭ�1�7QW�=��`n��BX	_�P5f���l�^���0���vۍ��ö��H
���I��|?�R��;A��[d��޷��b����T�/&(Z�t�8t�s�Zm�vC[��?���?�j8h*��e�؏����h=:A�h7]�疞���[R2-r1MM��f���\&:��޼�`Ă�H]T�wj[<��+W.	HnQ#�	�0/�6=��>��!5k�6S3�e����,�.'�rB��n~��	SEi<�A�����5Q��@��$�|�U_�<
���N�.���Dy�ֶ]M9�^���V���A���Mt��tH��\��)D�=�n�.G�7����[�_���r���U.%*)[P�u��s��X8
������d$��������*�f�R@9��ܽda(�^E�|zԠN���[|�Υ�1���z�{@��0LJ�F��J��#p�"��	,̅7�RG�s��0��C��C��
2�;>����+Ϫ��X������ո���^��j�F�S�U�|��H
1��3v�X=t�vqp���sZJ�T��ޘ3�(uQ�ԿCh(�Y%W �C�m��7Af8�R<K�R�L��P��vff��ċ+����|i)����˭�=39�IT�P�p_@��<�BD�=8���� {sW� �v����h��a�����h�ݑ���~������!�z�3l>N�!��2V����-�}��Ylhs;|;�M�����h��Cd�e�����sVHX,}\|�x	IT	m<
dXm$�^�ed��b���\��9p���2w�q��ڀg�*�r�f�Y��Im�c@�,��oU]=�8n�Ռh�t��@�h=�H6,^~�M������B���շB���P�b� ����l���.����E`�]*��=>����V�4��R;=O����aS����hx�;�} ̧�����O�n�$zf�t {Rݑd���E�)oY�8��[3}/���_�c��\�s��R|ۛ��<b$Z#�z�g�7���ؒc��� KV5��u17���F�?[T�䅔�
U�0;�#��Qb
�	G����(U�_YA� `�A�@�X����i�/����T�Ι]�-�N�$��搤 c� �"��f#O��"�Vֶ��wD[����]�����{e�ǁNƠ����B��~i�&O=5�{��>�CN-��
g��(��#��q4J���k���B~#�C��p��\����y���>�R�׌z�hA������.n��23��[�a+|A<�F������l�*i&Ěeލ׏��z�����N(���ԉ�E�6��� f���>V��dZf	��V���.N�r��p�,N���d&�<�}4�B��,� ڗ��Goa�.��=n��1�W�*��+@�����FA�o����M�p1~��fo��0�
$��C>\��IR���ќx#��Q��c�B1dp-�G-�k��*�Vv�0u���r.������c�R8�|�I��4�%*�Q���︉.	)J#< �̪H�2�VCD����?D����yw�Xꊰs��f�t8,�H��M���5�Pt�e��oQ��Ň�mb`jh�	�l�̀gY�K�a|=���ϝ�!=u3U;�]�#���<���˥��!O?υ"8�R�~Q��\���J�g۔�9̏����O������i�t��۸b��̄��,q٘��fT�����6�MR�2&�y�8��J'prJ�80}�����LJK��>�W�<q�b#ّU��r	\A'��,6C3�������RSR�7)�2(�4 �v(�`�Fx�A)�3�uꞟ�Bo�ٟ�B�ڐ����X�8�GW�ʏ����d5���=B4@�6�Ej����O�33�#⹦�쎆���cV?'k�*J�憴
~xz׽C�s[�\e:����P]�=S��JzQ�)4���X��x�c��W�vX�$Ч�8k㲦�1Cq��P���y(R�3�������K]KY�<�X!���
�	���=���ٝZ���:RnzF�2�����'���"��
3P���݀
8��I9��OD}<[�z������\������e�/�*V>�h(����gR��A�@γe�u��p�_��n���.��*��C>��p����_ͤ�ZyG��LL��63e���U��!3w�	;j9(v��*������4U5�r�1�#b�귡=R%�%����9XL�	�EVƉT�޻U5W���C��]��5b�3Oբ6f��L,�I������]>u�y�7��ȳ���\��e.��G���Jf���إt⯪?J�i�ڎ��V�Eo�?5�E��b�G��^�6��ꋔfF�7!�S�޸2�-;�DY��5fR���]���|V�l�}�6!U���n^� �ۋ`䴵/�f}�W12�~��0?=��:�MD]�"	�c�ks�wqDif��°H�
�NCe��k�|Ƴ����d�;�[����c���7Gg=˟��?�I�����y|��KS���8�v;�u�=5ߑ�:��k: �XI �S��XIūN��Ձ)�Apž��emt)�,�4y�,���0�2�|��a��ϟ-]�Y�=¥�d��f,q���6P��s�K�Ah���dd�A�\ϯ0��Y�y��O�[@I��`� D����D{m&�ٿ4\��[;7��Dv��ۙ�R6|���Ȍ�8��R��^C}X�WR|�'rP�_O�
�R�m��'v�C�W�aWp�߭�1�-�{g��.~1���x�m�,[5�{��)s�L�+���f�﹋�*�vl]`d 0�X�¤��TRc��������0���iS��^��[��1�b�����*h��]1Nv#��?&�9�S�]�B2G� ~Qfߧm��`��YP�ރ�x�%�, 4OQ���qAc�N7�Z�^��;��3���f(:
J9c|�tI���KYX�|��>B����roo9˺SQj��A�����ܟH�,����{���	a�_Y����)�Qd��
ݜ�,֞5����B���ƶK�)%*[n:��s6.�d����,>��A�Ă�rR��D���k�*E���]F}���"_p�V�08�\,���=!�1\�:/ۘ2��4:����&��J~��
X�,Ģ��?!�rNǩv��/�Q\-���2ԋ.�2���.W����[q��}�g�e6�!E�aD�����O��0�|D@����u=4�ٺ?v�֏��a#N��u�-�S�4]D�=��P��As��g�ʰ�R$��ho.�S̃͝~fd������H���f��SiA+����2)߮A���E3rm�o�o�B�YF�8OI�T�Q������d�@�Y�O5�c�lp��Oc ��	������9�<
M�o���+�����v���-�����diI]��ZÊ�c>A4TZV���J`Z ��v'N�]��~��ѭ�u�&	0x�в��i5�R?��'�T^��K�·���cq�'1�k�E&,_	ե0G���~$,Z���'IÜ���R�sYx,��ͣQ��SB�C#���W	�TW/nQG��� �&�#Yf1�g�,���GU?2.B����W���&�? ���x.Z/*�c��N�6)�<G�����G�,m��)d�R��Ȳ1ż{Ą��eU/9�t��^��y�k����vH[
���J�oA�=�'�ƥSR|��<g.��?�����	��W��BX�@���AH>k�m%tl.�hK��a�Pr�f�$�{�� ή����C	��ݒ�3P\��Y� �1�^<��ع޽U�|)�P�w4۲Ml	ʗW47,���Ϡ��@<���r|��=�sj��}���(x˺��Xt^W�쫝[�_��u%�3~^3��r�a7���@p�Ҷ.�1_�V�]�WG���u���O�}�:�E�|��F��L��,�d��`.Ug�0|v��S��4҇y)�8���aZF�\�<�4>�
�r��l�C!=Q��v�9��Qv�։$~��"���ĥ�>�֘@<6�=���,d ���֭װ�v(��n�y��nN�sy�!j�w�~��E
���SZ�|��ms�o!^f�n;79R�(Y��~6}��[�Dr-X����	a_��z����>��Cں�?@oq��g(�'0D����sO��/�0�Yk�`h�{�8�@�b8H@?naӎ)k2�J�xgi˶����]�ǁ_���/2�U���[�&7`�w��g9Qǽ���F�Z
�8~���-��D�W]�u&����^������&bPM�J4X�j�0$�i0��F���΄�?_��S��J�B�?��B�q�֩IzYHc���r�B��ڧS�)-l�<�p�L,-k�K:$Fw0�]����;�#NܣI;�V�H_di��� i���*ow뇹ٍHM�X(,�8-�Mg���;���l �&�?��BY�0n�"ݵ,�v�U47����5��<����b�T`�>�MYKzFl>�#+@
��E �kH����������a����:���kX����&�@a�+�w�K�ȍd�w`�ScG���
������Ll��V��bU`%���Ft��$�;����t�o|U���Ϧ:Ep\S��1{B2��nB���vDn�u_7�-�5ڿ���SN�>1��T��A��������K�Ej���[:��F��K��������u�E�i3�I��rKC�󯁒��F{o�����s�:�L1���lZ6B��b��3�z��a-sT���xAڢV*�����yg�.Ԝv��]�$�R%2������,��c��w�vm�[����Ҫ*��:��f]mo{w+#/Vt��O.��;g��N�µ>ƞm����wuA6r���t����|�~�K6��ޡ@^�����a�Y�4��&@|�dЎÑ�1�gB�D+�1t'ŀ�� \�y]a�Rf/h��o�Ƴ�sp1zw��t5��;�/��%�����d��nM]�3|�L�皾��c�[W��i۳~���tR�Ke�k��_r�E:[�L�ڐ��� ��|_U6Ր�:�Rp< !H<�d��2�$W��5��Gi�������L���߭�5b�@֨�b�o_)C8%����9�MC�����n+W����O��V���P�ì
��݊6f�JbU�f�j���&�*���E/�	$����Ƿ��b�+vR�y/�f6>��:e(�~p��v1D
��tO�H�����;_�'h���`"	Ř,��w���Z���֗�E ��!�w�����t�/7�z�*@r�o"b;뽊x���W�d�H��"�<��JJ4%����1ӛ0j��e�'�8����J���(�/�Ot���l\��Q�N���8 [ǕH��A+"�p����/xn(������^cj�i8R�-R�({~�!F�:��BS�2t&Iڳ��&�̀����@��.���RM
�
��XNk�V7֭���/ �*r\,.6���`��)[Ǚlz'�eY���2��jL�����C/,�O�<����w����bd� K�1B�u�u��.�|��; N����C�$d��NER�ɨM�0P�c���DOزc���9�$4Wh��jd��KF��S}pb�-ςqa�0�f@��ߴ�5�X@��+�� 1Ю��U\��j��E�m,XhoZI���m���:������P���Om���hL�߶�I#�4n$:��EH��\l�:�SiQ�s%�w�=������d��)�jiΌ�3�J��Dq�GB�TY���Nv�`|m�]�,�Ј��pc=�c���M�%LUd�����̲ �Q��ި�Ge:�׮R���}�D�:�d��\�v���5̎C��l��J��_�REv��])#+%l�ܕT�[ �Ԕg�j�_�d�^������vsb���B�2=З\U�� A�t���hٻ�G]�y��'�ؾR�Qe�"q��h晵�g��~�_H�3�\2nA_��Prb�_�^��
�vW��m��;�Ɩ��ZXƅ����Ï���4m��Mw�C���- ?Q؉pRe�����:�Z�f7VgX��'9�,�?h�����q\ȃ�؛�ѝs���VYX��Z�� <��A����e���3I��-U)��aA]��o����#���C�<���{V�����dC� �F	A�v��<�M�zW:TGM�[:�j*��I�1�uB��f_9~?�R{E��6!PJ+�nBm���`��	kȍ�'8�.������-"���lN�S}�Y؜�ˮ��X�F?qBa�Wh�sHդ��\8l5�,�vzь[�<>F���A��ve͠�
YJ����������7����U`�0D��Q�J�ٴɉw�����X�M6�lF�����T^���/�g�����zJ)F���s$H]����y�:�����n�y��¸`��[2��V�@��+�p�å���=5�Kr��O���_�,ڛ7�#�\����r�2�s��c!zi)�� ��)(�cu���t��7~W
rtE����m�VP�$��u=vk��+ǀB:3_�rUss�X^�X?�V��u�Cj�#<��æZ�C�O�g�TNL� Xs�H�Sp�[byuV�����gӣ@%B�Mn�`/zǰ2�)�dR�8����"��tI�&b߶���t$匁Q��K䵨�,w2.��ߙMaQ����/��twk�1P7`�ѷ"D��a��)�V?�?��fl���7�4������?�V�n�i��T�K�|��KM=�uݛ�r������B�t�	J��Q��vw�b��=� 8����.�i������uQ/5[A/��6m����ީR���蘦!Ǧ����`On�R=x��Q�p�#[����Q�eKxGxD�`lEȚÊ�_IA�Rzّڌ�K�1��� xd�z����x�Ǡ�wICJ֓.!�<��t��ɯ�G�|X�;�s�H�xe�z�$����!"����k���O�l؆]�8�&\-�v���rj�`)ݱ�9H$�Wq\V6��m�~�LM�!6���F��AaO���7�Gbo�����2���u�~U���NUw��hS�c
k��m��wk5/ wH9G���ig˰&�q��q�8��0�a:�X- WFG(�BE5���M7�+\['yq��b�߁�}�����~�:�<d���	�
K�R��=vZ��?��.E�
�O���Ճ����;��sW ��R���gd` ��w��P.n�p}޺)Q�8�`��?�W�9@S'����ؔ �JtN�	��C���F8��?�43�H���1������ҠW���P�NM��p�d	:��4F�*u�XS���.�V��4>���x_��� ��(�씱	���?ŗ�ip�h��uJ���F��π����#=W_x�9rO����+؆#��b����"�/2����,?���b�Jk�¼��j9��;<\��/.��7O��<�����JX�4������=5dSWN�@e�P�Y�/�0��ۧ�G8��u��X�-蕫Rm�({���V^�#�@t�!����y�pi3��r�Y��:������*�l�L��B�\�K�o�i�Z">ʱ��`�����P�)d�e�,��u=�if	 �@3��`��:����͂�z�����{ɪDڏcR���*��hYr����:J�F@�t��xә[�fםC�<otAD���,"���b
P��:�;_�L�A�لԊ�c���p�1㡹��>��f�#�ĩ���'�;�}�v�d60U��l�1��K��X�oo5k.��3G.�?�T\��=� �Hn�E���
~��t��d�/k݆7�K7����T������Gj���N�]��H�{���sY1��<5�|�W �@�����-��A��h�.�C���M���P䢋J�R��H���*���P'��6�vJ��� \9��	��U��$��(�K��?���u���5���&��,����9F���p�C1zH?�]�Rt����iV�5�Q+��D9���as�� Q8�	9�hP��T���
�+�� �˹��"��S�逴��ɋ�S����|�Ff�DQn�G��b��e���/q���8V�g�@�LF1KA.�*8b��"~I�I�w Lv��mU���彦����'7h��I�(����ote�:i��{O���.T/�g�9�� ��v��{x�V,���#�?S�
`:���yX�c���׸C��a7`��k���O���#nUV���{>{�5�h3��. ��p�7>=^�
��1���Ν���{2/�N�%(lյq�~��!�5�O
s��g�d2Y�����	k-d\������㭿;��Y��GG���lC�����W����{~ƻM[1�!�[@$^�/@������9{����n=��,���� s� �eX�`B�iܺ���|��� �B;P�3�6�+C�U������A����^�6�g޳���
�����7@�~ ����S���.�!� �����vD7]$�d��!Pi�X�����<�h��r,@�>�����V�.P����^�,c�\�j69�GAIE��*iū�u�,��7FZ�Į��Sa�@@\�L:��x�6;�-�!��v�F|=T��iI�8��'p4�hPߤ��ē�ǵ	}��Z1h�@�i0!����{W�N��M�kw��\�N�3u�$�vO�-"��v8t6� �7���f1[�JV���W*
4��:�ű�#�h1m�]L��/D|���[2��&�a��	N���ro̟�9�@���A�X_�+���֍R^R�_^�K���b�#����ٿ��W�o�Uϕ�ݏ�1�hB���_�����~�������w[�V۴kу�=wB�̔?JZ��AM6��
�thA��3�Fl�P�^�W	��ꖸ�hK����\�o@^sLǹ���r�}�H��P����|O)���R�x[��?�kC;�PᛉWM>���܀J$I# G?�ZSsZ^�}_���@�2?ш�:&^�nÆ�B}�ՅrGО�t�l�B�� �*��; ��C�&�ЧJ�Z�L���b�L��e�>�b"î�}+�<AJ%��{��K8~���apQ�(��DH�s��|�6��h�4ܳs�p�*Ch^�ޡ�Q$WJ�F;�defX��o��n�m�����ݘ��ϗt�$�[�m�oV�[y)��y�����Pi\7 I��n+4�y)I�T�����G�8���S�b�ke�O����l��u�!ؘAe��>;t6�p���Ũ�mq��7q��O�S������;p�VJk�`e\���DJ�� ��_-�4+�e�t��Y�4��X�µ:��p����$.+g򗹳)|�;y٤�y��@�N����5�����Ɉ��hFW��Ѽ�Z@��*��?��3��!U�0����ZYjU�̇Rz��Y����H/;�!Yp����a�vjse���U�'�u�p0B���;32�3<�-�Pq�4���l��k�-U��]'Yfd.�)�����!^3��L���_��Q�w�`Y����w]�.�I95��5Zp+�Ā3i����
��: �?�݃sH4������5/�P=�PQΨ͇9߯���f����ɔ�@PX�9�"\/�Շ�w=E��U���z�<�k���+�#���Cߏ��g�Pp]>������ʿ,e�`d��S�tG�hnWdƺ�pH�*��;_4*�"D
hk��X�������}���*�lOϗ���\0��+�;_�8*fE���+c�@�v1�N\mԒ?:���R�h-�_�}�I�ڟ,5��K�� eY��#�V��.^	��,'}3���)�R��bW��q���C�n�Ж�H �#��:8n�� �LY�������bҟ� څ��x��l��\�:��e������hL�YmK�����l�vR�&��՞ۣ*v����ݟ�W�ۯ[�`w�'d���s�ʩr��~C(Tn^�+J�[�C(2_w(�R+����vyN�ȑ���U��ˍ�BZːE���O�{��樰^R�6�V�#�ç��,�'��wC�����@h���q�=��.��E�;bo��C�d�Hx������ױB�(��k�>5�{.;�4ا�r��#y�c���1�@�2�0(��CG�n�N���/�fiJ�񙓎�;�+��#�qu"NbZl��J�ѱ.�8�T�@{($�})�KU7�;�<�c�Z��H4��kbV
��%�L4�eA�?1��Ok	\�
���z
�u��E�˅�!PM}�&�OQ�_&�b�"�����9��Tz��7�Z��8��DuD�Y�~�=���9>l��?Ĵ���F��]���
�w̶��F���J��p��F�@��˥�;?�q��j����B�1�ܶb�*��?�@�%��������^�|'tM�=jH�2�
M���Ʋ��m������]����\&b�����2ɐ��w��%��ڪ����/� �������ŜO��{�8)d��A*�t�Y�q"m�{cU�ʸ)�n��Ҩ/�c�"Z��D���L�z�?]�!��yO��5YV�s��M|9BM������*�d�����C�뤞��8���g���(�ƀp����l��@K?7`z"kd�"lM��4#��s!��V^�LDZ�^�{���@����A����SJM<�C�H�"U8��*�`���sͤC
��N����6&�x=cyd����D]Z�V|D�{�#�'8��V�e�U�ޗ8�-�g��.���f�c�K���7�1e_�S���;"H�����oxL�t�C�4�e5�����y|����r#�+a̩�)s���+�"j:��Ts�J]1z�È���}�3�&NsgP�+���݇Z��N"�#�Yޢ�'����oki��;:>���-�"^$*�"�^�kL��b��=VQ��$�7/�dG�l]�8�����T�o�D�9L�OD��msz���d�r�����`[�ytB�v�� ���̊��uk�s��� }!��s�.�I�)�����W��@<�Yg��1�_EƤ�K�{%��7miqz#�}����<�*=]�W����`��j h�`���j�(�+-�G��P��p2���<<u�x��d���fHiI�~�� �s>ݾ�������:8��g���Z�x�hs�6��Z��#N�fs�8br��e�[��M'����%����M��\^�(
'O?��m�f��ɏF�blk��俸�U��:�YZ�����U�Z�Ck���b�5'��c�6��b���si�րڌ*��3�9f�1�c���`cr�v�
l A�p@�&(�ۑC7���R=��t�����k׆om��.�E�G�p�np�	*:�$����8M��f��Ŕo�s7O�/���_;@�����aFQ�wἘ��V���Wu�`W%����CB�c�~�K���I��o��f��!ž~Q��g"�cKPݢ��w<�X��jH�����0Su�6�(휬�1*W8M��Oj�y~�^���q�<6��zk��u*��|��T"&������!"��b1^��d$J7��g/b�ࢪR�i���6A�N�&
�Qx��4��9Z�U�+�]$���9�p��1���X^9����k���� BK��8������)�-+�̜�r�D1|lb*�,#���t`�BP�~3��3�}/G^*O|��x���;�#��vD�Y�/���q��4�.@�X2q��2ed4]��z6+%:��e����[��c��r#�O�Hͨ�[��"[����je�V�G���;���v���El]9w����yy��
|H�:)h�i~�9y�][�l�B���ԭ����4)�ǧm�"y~2���������Ga8�:�f�b�0�����8���fZdA)��0�T��r�Xl|SO��hN������?�������@<� ����\Ҵ����ͻ��`*�m+��.��0{r!BUn�=1�����Ȝo��r���p!�mfY��qI�s62b�g-5J��4k�����d䨵�v�4B��=�!vc���'['"���J�_�Ez��Ȋ˗�Yn�yD+�%�[[2$Z�_���zYgl��3([C�9����[��뽱����N����y���ʹi�#]�pDsUaL��.1E2���.��zTh���E%�&��GI�w�c�-O�ι��j"���s�L%�/�}����g�ւET�򤲮J�ߍs��XB K.�J7�2�[F`����z$=�Pq�!"=n�D��G��,g7�B#U�8k��9��c�����?1^�S�r'�#+���H��:���:ފ*o�F7w�7�i�`�(�x�Q�3{��83�BP&UsKW;@&�]O�I(�,��~gfw�?���'���ʺ�{8�`G�H�k���ӋM���n�g,��{��	�&�<	.��52(��w�ߩ@$.�r��0����Ԉ�K�&��_[���y9F)w��.Y.�o�~}��1Pe���N,���I��EX��Q2ONY�J�d͝�/��J������w�%����ja�/�EѦn�g�5�6���9������e�B�>Rn�呪x_�Q�	��6���ង����u�]Y���,��ӀdH�j������
��*)�Z�G�'x��7�08$
Ď�a3k�ñ@��Qsht��Ib�,:/�+�oLtRԋ(0 ������\���SD�D4$�@��E��.��&$]?�p�- ��K�O��/:�
��Rr�;q�s�#�*�qZg �5hH���R�^�iC�F���A�rq*FU{Kx���Z��(4!�m�.�PGNɟ"s1W
PWw��e��V�cdj��7Ѝ���;qV�4;]�qY����@�7�VE�b�������=��P�9�0�FǺ���#�{s���`̈́AWgҥ �%Gy������_�����B82�t	����w�:��}ՠ���#�s�FJ@�J���k��k/$��Î0��E��b��Im��ύ-�i8�0��6f�/3�lx�[T�X�W�t���0�d,���r��Y$�A���t%X��-���/��i��[I����
�(m&���r�W�z�� �4��6"��Q��2f3r1
�m���Ue�ݕZ��+w��n���<$*rX��
��mA��� m ��M�a��uߡ�&��-���R0/)Mc�l�Vzx��@�l�Z����\p�HȊ]���m&�c{�@3�Gp�MT�l��:�B���D����	^}Vc�z��o�}�n��J=�':��|����iy%*gZ�{yn'Mu^�x9e8�ݭ�{N 1��7��&h�:�?��/%��@d ����!��K򏅍rivC��7yߴU8�ibD��(R����F�� |ڳ��ڗ���Ź��C���3#�d�qhC �]�{��9\�ӗ:t/"Ϭh����?��� ���j�a_�Xe�����,'�ӈn�9��b%T��}~hg	2 �v����N'���+���р/�~[�]=M~���p��jjˬ<Y��%��=���͓נ,�Pq&z:%��:�F���x"�Vr������VI�zi��c{gё>�/e�B<4f|O6�QIW*��OOX���d*a�k�������NhfL݈�S5g,U{�n�4����e��k�.E��ʑʅ%ʵD�����\��'��%����P8�wyõR�$)���*�di#�דl�4�T��<��$l��W��Jc6��.��Y�e��I~����<��Yά���Ip~���n�U�.�)��Kd*Q�Ob�y����VZ��s牸�&?ʁMe�CW*�2\�AH K�]��_���^����z���1����uz$�_�=bB�Ţi8��]�i�3k���>��+2P|c��"y��cs��0Τ�Y9bT�>���u#5<_���m�#@<�=���׮-�3r���?�G��֕�u��5���n-�y���ڝ%c�) ��I�m&�}��j�W���AY��?�j�*��\�$.p9Ż8
�;�.���)F������8g�(���	`����!q9dux��]1�]غ����K5��l�Sਆza�L�T����6�Z�b��[��*�y`yi7��R��f�X@ϼ�o�LiY�XG�I�b{�)���O��MD���P�.����hg�7���^�/�wַ:�$r��-l���l�N��1a���G[��Q5�� �u��X��✉�t����������H��:�t�Mb$���_���w�%�}�4�?Q�/{ߴښ�v��&�}f��GA�[ι��i�Pl{Fm�<�FZOX.9h"C�<�Mc80D
��a'�OA7Q_��l&0��o�D�ɬZ7e���T������R.S��6*L�1(]kF����R(���S��{�a#0-Xr1�&�䌸����3^:q�׺#	�U�5b�U���{�Y�5�hz�����bb�Ă<a�|2WOVa JSC�����.@\��9PRkr2G<s�?ET�j����TϪR{�X�V��N��X�e����R췎zD\r2��Z����<p�:ȱ;��qҘ��O�����9&ɿ^:Z���{��'=�?���*�&�   hL�`�kK'#N���*�-�Y����#|��a���sw7�3��R�K���*.2�o �F0��,8��I�������[S�3b���I�5"/9�~6�?��  9��+O|u��d�N9ϋ�VQ6>�̒Un�,>ė~ծy�����]0��̄`k������!)Ѕڹ����1'�ׇM�GYŗ�=X�����h���5�����J�ʺ���,.g�B��֐W��:��m~��=Y?mM��r�"�t�F+vH���b��o?N�"���>s��� ��ċaubLc[8q��� w�C�
�3o3��*�1K>��:��W	�Ƞ��ɬ��&O���<�Y_���C%�+�
R@0.�	������K�"�'�
�b�� D���I�}�{��k��L��1���ҽ`�D���R �y�XH�A<�h�	�-@��q/Dt+ǎ�|DwU�ܰT�F�jK|�DV�\���2�-5&ޖ=�0�u����U�R�>Il���6��֌7�l�9oni�֫n;��"�0g�"���v��w���U$8����WP(�~���e/��a��tD�8�7�Q1�}E��b�r��лsBޗ@5mf�ګ�^�Sw9���/ �`�i����UE�����fb.P�US��p�G�܃Zt�t�����|ʺm�s�&뿱Ymk���� 4
��f���Q%����d�MD)�K�ev��؟iB�����V��#�Dr����Q�q���V�>�o�Dt��J�������	��r|i0����p z�h�]��Ժ�+*�&��`J+Mj@��)�h���B��S%�Nt3@x��GLgi�P5�/!+�y<����p�D{	�F}��T�c,o�=Q-�L����^��|89�&��ѧur�Q��r�_y�� {�ʺ��O��B���D��F�t�7�9�J�����mߍP���(*1e�Xd�ʽF7�Mry=�<V�CZ�;�B�����"6�,�< _̗�G���v%�A����	ۄ�4�ۅt1��`G��t�u��=C>�"��z�wb�1S�����v��:vn� Q��fޛ���A��`��=[QuΏ�y����Ӌ"�	��u���z���t�\B;ndw�9Qs���ŀ���0?�ma3��EU1�'!���*A�A��������Ūd��/�Ň@3Ч��:�ˋe贰��i�@n$��s�_�\�^�1
�*A瘿����|v�qhS�V����{|���h�q�yU�
�a0��=��I�1�Y��9��ݕq-\ 7���Cx�3{؆�t.�ȉ���ä�[����� ��:`�'�����]ҾS�Y���ڮ��q �W@�߽���r�it���1Q��K��~�����>b�^�	ĒuG���G��`��A�ICro�P
u��>ӈA���J�5@�ĲD5f�F���%N�
��a��e��`�%�)2�M2�L�u�v=0ˏ��ˮ��w^Ȥ�Ҕ��0M��oR���P���絀l���N�^2�	f�mF1lբ�k�� �D�I5��vȄ�j	~�RBB����u����
�S?�EU{�(�M	O<��x�weɨ0g�F 6���k�����t�-BM�m�a���/� iX`����V�3�c�;�t�p��� 8'�T�F�A5?7�������	�G]ʗv�������9��Y0�m!�	����v�V�x�v�����ay�ր�����!�Άkg�V~hz1�-�4׊�ۖ#5��G7Y/0��t�������V�3�|4��m�T�#�[2p,>X�m�/
�~��S��je��'V�ξx�D��4u4���z�XNH��e�hz/NG�H�Nuah�N��A<��Dp�R6%ҋh)�1�rX�&��3h�e[���X�g��o���n����UM������q*���g��6Y?�\���"b�*g����)I~�Y�7��Gjr0��a�@�p��:�d�i�n�j����nrT~�<�`x3�
*(1�Z��rDk����Y�K(û0��{�S���`��*q��o^۲-/�]��]{w���c�?<|{���WX61���`�V���]�w�<7E�dE;�*�����5��`b|�k�,�u�	�?2�����p��3���J�c�7ie.�X`$&ݎ�a�U#���]!t,�]�j�C��h�wm�@��!�G*���\�נ�Q�1��b�ئѯJ�`M��W����џ��7�����س%ǃfuGD_�1~�Yp��l뇊��;c���Gji�_b2$��G�$X[��1����"���JK�_���;�J�`�x궱w)U�Ulb3�?�b�j�-����_J1��e���Fp2�S��뫃 ����G��H��U��@BhK]	�Ʋ�
8���(�6S%E�K�m�j����|�6���XT��]�Ǎ�f'Q/���+�B&s�<�J+�5��R�AM�&��Y�ϊ�'A~[O �N�>h���U�s̺z|�L�����\���D�4
�����)���T@��IS7g'd'6����{TOy1J'�9X��'#aK��.���9�ћ����*�ʰq��G�ת7"�h2����U���}-p���+o��Ȍ���;ot���Q��x�d�[x|\���Y:/�]�Q��e:m=����oT�Q?��U)GI1�G�J��k������!EQ�	�5��P�r-q_��X␣���毰�$��zUF�3�p �s�y�<X�<x���EJ�a�}�=�:,��P�O���t�K����<:��v�J!����f/d��B6@�^�t6L�ȓ����N]�>>���1���ί��U��%�Ү�N�/����ng�(�Rl��1pjm�SѠ�DX_@���g�Am��H�8R�V����}����U�oNc�I`yR�3N|r
�/�����_  \��L��9B�4Z7��U��!��S|o�P���D-�W�j�L��
��Oa%��P�V��u��`�	u��D@�+D��.��0��G5�����
'��<Tjo��~qYRB���F�J��}���l���ObA�2�>~�NQ�ck�"� ������. �1V5�E��
����4\������9[���3�;���z��0�e�m3���t\}-�9���+��\Z(Y�@�gD#G����Lau��b��3��B'��X������h�K�Xח�f5H�i����5�°	ڠ�{!Fw�� k�<G�"4$�A��!���ܠ�^GI���o)��j�q6j� �x�JL	47r�/,�@�P.��f�b�`D��
����\L��c�x��|
���������M?̑����b�Ge�F�j����Ј���=VPA �[�~�W��m~B�w���t$,��Zz�?.�굞��ғ\��� x�SbīNZ	��P�,0�l�y�>��:���'��:��Y��4����(� on�CA+���[�jQ*���ֵ,@��F(�{�2ν��ki�K���&���F����H�������(�y�+�$�`���K����:n;�2���J�V]T�����O��I��h��ר��!�a�a��X�H`:k�A�p[���uN�-�>����7>��x���uvK�.9��lt2�H����M�*�LN�m]gןԥ�1fk� ��p6�p��ׁ̚�?V�Ty �od�L�I�m4�X�z�=���(�U�d�@���VcG=hP7#�Rcj|S#jx��Zq�\�b4Ҁ �q5��ࡕ�ih�]���*�B>�4�$u�n��!������j`dzHq�q?j�����$�1�|4'fwV��u���g�7�PB�;��	����\�9+�,��>e{���˓�u��+���6u!<�,�p�����#u���y%��q��V#K��_X�yn�.j����#�FP�)�U��:Y_FjX
�wp�P��0([����ѿ��}�*�ŧ�ɌT+�k�k���jB�]Sc�3��eAvL⫅s~^��l�3h�/�#�-��N*rhn �Q�]�2�'Q��ό/��}�~�)�y�r͆�iq��`�I��o�=E(5���M׃.����2����Z�	ʙ�������t�s�[4�����9�ݪ�y�E�cKL�AL�Eq� H���5dF�:��n�/����i�\���Eb�L4�HmM��ǎ'���}uuC�P��Z�����$�`s�ū��.�d���1�\����T)�?���T#�c����r�&�*D3A."S�w�T���U�gu��OC������^�nv��0�68�w����0�~��fF`&'y]a64�LX'D�x/�����4d�����-	���t׫���������T�;�����1'�5��f^�z��)ah!�)ᓶ-c�==Sdi��#�1����Kv�^���
���n���	���>������'����J������wV�����4�8��mPǀO|��󽄬�@��,��Z�-Zgw�]������S�(���,���q�#�Nu[(ۘ���&������}��o�`�[ ���.a�z���[T�f�~Ե��k�Q��E�~(�OL^^g$�Vt wc�F ���~��b�Z�S��+�
�ޭ�m�!�Zǘ�G�����X9_\��6.�R�Is.jk�#;n�}AI��W�"�x���Qܑ���<�Z|68n{ն�:`W����:�>M�N@􋒙�TM�bl�s1=�{��p�ZD���L��f4�Y�J�ј'I)c�l����]b�x�����c	�#�q�%L�$F� D���Rg�p4Ŗg�����9�r��@%���� {e��̨�+k�U�\V=:�۵mR�������lj��}j�R��@C[X/�*�l��--SV�.i�NJ_\���F
�{R\f?�"���8�m}f��(��kƜb�4@�������[*Y��p(�u1Fv���S1��x,�"���쏣��T���b�ݮ>���X�[�����u.i�|���r+h�<)��!�j�xs
�^&�oZՀj�k4^� �1�~{OhѓR�8g��p�N��q�I;�N
]ڥ7�����pY?ݩ��hb�K��(�5�:($!6=F��L�"vƂ�W���eф���)������x�ʜ�����H���agJ���q���%D�!� ��hi���+W�o�nh YTXN©)@� �פ��\v%(�6�2�*D[�!�w��m��2����ir�s[۾:���GV��'�#w���� �k��.ˍ۞��U�&.J��0��.v���Jl��]�),��%;� $���캕ٿ�>s/V��}�5pȀ;�d$��!�t"*�F�30��Ρ��5��� T�������0��tl3>�+��*�%8���cd��o���,Z63C�3W;����:f�4��$�N�Zt`��^�CD�ca|�R���I��&i�!�#��o�,�i�@�+u!�pR��܂���):��	E���@Jg*�i�^%6�Aё�,�Qp���F�z�uh�ԧ���S�L��S�֫���w"����W���L)���L�#�����o]dС��-��J7�w���� ���Σ�T��˂4��_�WZ�y������?�s;�*�r0eQ�L$�n�C��ml�O�l9�&���^Z�p�{�e������b���,�Z��cBx1�w6*	-v!
�-f1��S$ɀ��L�Z9oŌI�ʹ�,��C,Ň`ّUz%���]�����9�
G{�\�����r�h�i��J��|̱Zi���K���{���b���~�������C��gX����S�5���OM�9|g�飽�d���B��_*�e����eA��	;J�Т뼣f�)��և�L��qWD0K�U>)%��ԽƅCZ+�ԯ�����p��R��z`��#�~���l�:���R����>�a�ټM{tn^�_J,�WN�U|Aa˹����U�_&��𙰝e��Z����Z
K���{�54!���2JܪȇC���׼�M�	�����n�0Մ	D�~ytWc���=��R�q�O}�W�}��.�ڪ'0����F�W�Z�������s>W���:��ؤg+I�40%�I���Q�����O���N��<��� 5��&��★IV$��b�Au�Z֌]�����5�̩��/�����F#~]O��{_�uԽ�c���X�$�p���N��ym��F�b�{��Y�g�cf�7ueV�(k�s%��9�c��ih�����4�ңC�� h3�z���0�Ɵ�lj��O.�.ɹ)[�ѓ��Zވe��4�๒�D�#&�j�a��mV�UĒ.������xUz�<w	g���Kd���z�2�5W]GنQT���o�h�A�U�O���0�%���1��4a>�U`�3=���h�k�@��
�i)��I���K;���6�Sk��k�� }��!��8�4��в|[%���q�R����,���6�I��g�2x�{�mj5�����]fH���Dh0�W�GLx�j�'q���s�Y�\����j��5s�kH=�ꢥ��rȓp1R"#Θ������AΕ�Ř�832ǐ6�8�ǒ�(P�}�W���qp��܏�����7؝����ӉZ3��A���l��d,�B�a�����"�$gǇ;�����F����!<�|���/36�|z���r��uO�Zw��`M� � ��^	���I)KS������V�x�N��BFS؎��������kfT����Є�.]&�:�c�U�bU!�B�,v�M؇	��?��D��*3#僁8���?�E^����gw���&X��,�3��b7��ۓ���y��j*�qm�Y�Y6=}n�I~�'!�e`��J�/�&��#��Ώ�O7s~e��{�}�L�?������8_���!`��Ue�F�$��1�e�;j��)7������0�a���#���O���:�CRN�$�hi��dG���r�����+Į^��a;6�N�Q4DBDv�>�冨�d�8[J3��u�����Ц̓�Y�Y�+�����k�E�f�V������d�8���i`�("cO���a����IC7��]M`|�9�(+ǳ�vw�\��f��ujP�pR��`�B�|P$�U���7ԽI��Ү������`�+gF.gL�g��(z�3T��kE\箿C"�m���##����lG�Y�r�t
2�J;�yp�,en���&�E|�cĩ#�ܪ�9���d�L��Nʏ�{�=�|�f��L����b:�d��EW`9[w>\6����MY���@A36~�Y,0����Ȝ�-6V\$� �C�mO�i�GHǮ�iM�T�
I��á����w{���Z���h,�Z�l@�	���'ޙr����)шQ��d7�w�̚�~bi��?n붇����9��)�Xr���\�:v���'{�p�0)1��6�d��3�Px2��Ik�`���|}!Ӫ5�qGw���_��g#7���{��7���od@ڻڹ���v)Yo�����1=)�`��ͩ�����񛒵��6:c�ʽv�r{#��k'����V���"�Z�'���u��!压q̀��3ԣM����Uj�&��E$���If���8�� ����-��X���V���b�4�r�٠&/����Q��]��9�J��o朒�SQBw�ڭ�sn���"dS(�8V�������Θ��*19�uݯK�>����{�18>�{�]�=z���qq�rL?b6�R�sU�L��.uؑ�Ëo��X�&}�pJ��pW�o��j�2������A�7� ��Y����f������y6FI�G��[�X���j��px�搚����W�۽ksR�X+�;��.M�(�b.H��<�d��K�:^a�2�[ºH�3�����g�l٤�:�Fz��.塸�H�-%kJ}(�喢6A��z��#
�I��I�H�o`*��;#����*]�PM>9��Z�7E�3t�/N�����7��=S�ԇ����w�y�� �O�����I��Kh�* �
�6l�s�{�Vx��)-�s	��k��.E$nJ���+�a<k#+����s���K��K!m�-����j��@���거2�v�2���NYk®��i�����_�Z~����H��t:��� ٚP� /G9�6��󚓒?^�FC�jA�a�I���w�Ǳq�u��9~5�:Ɠ-���T�Sb�Δyg0_$-����1��yCJcs��=���UKT[o�X�EC/�u~!Q������J"��I�w�O!<�jJY$Y̹	��d7�\MQ;���M����~�й�c`�K�,H�_�{�te�|��d;-n�Gw���V2~��_v�L4�Y��sc}$�}� �"���&����&��q�� ��T��d����d�u�.�j�o����@k��3Q�.aZ9��+�m���io�lP�"�����I�YE��͔¸�Jc��Fމ�c�̗�I6��x�l�-j�4h�F{���-�F�q�a1`.�e�����"��Rh�.LS5�ã���q��zeb>�+k��*��?s���E��pc@X�-�T��E�jg�u��Ly�A7�w�9r�a�M6H��?��g�b�-cS���������Kp����Q���=K�
��i�'L����e�{u!����:z9�X4�5ԉ��˰���y�I�g��-d��wl���~�|L��Q���RC�+��[�rv!0��-C̝Y{�2��)��R��������V�2�{��F��<�+�=!W�[������9��"n�L�ٿ���S�vSZ%5X��3��,ꄟ�-6@f1���3;
��g%��1���7�����oe�S9ju�hjE�!����<2��٥t�p�U!bv�w���<�P�+�\��WŔg?)^r|rgA�>����GP�I�d�BC2�S��j@%��M��}��pQ���+�c���	i�q��uEB1�rCQp�%��=C�S�����i ��f�ِH;�X@�f?|����d�����PR��V�{���'�*Hη�Dԅ��ʕHV#iz�a�<��IBJN`I�T���4@1w+(00~&�|�����5�el�f��#�d�I��}�[��W�{}��8I�&�ʚ4[/�t+MT5�v�O��umÐ�}y��(,nW&D�59ԗ�IK]���_�O[RA����>r�x;Z��8T�l��� �/�� 
o��%p��"�<�|�����y�,�w�Ѳ<�N,)����g�Q��oU�<A���B�+���$(��G�}K1l������X�G�<s�ŋ4�����A^�7��{�FYUx�j3致Sp�](��c�dg�3P�'ȺJ�m���\�G���C��@�{���v���.�
����i�a�8�䴽+�z���u9#���@HNF��4.��$z��pl%"s�.�#+�XL�Ͷ���BB��O�J)��K�0���=j�im��aE�q"�g����e1��]r���7E��ރ%�������>E��gK��k�o�XA��*I�)_�ۗ��Eր�P?TWp�n+��Nj�7<��tn;7F5>��-�όb���9��9u�>���Z��V[�o"���5ִ̲����_�0���)c�(Pl�	�}3�U��U�NI�H$/�&O�أ���(��D$��˫�w��2[W����$]����=S�����_�ya�б
N�΅���,A<RqUqZU�a���k�繊 D�a7q��Yw_nHHgp�G]W{\����M_�?�,�'���i��9�")2��'j3��8U�]����#~9���f�D·m�b)��FT�i�����D�|�OȴW���ƻ���ߖ����v�ҺB���������
t'���4tC)ST0�(V���I�)h�9�\%��}���C��zZ���J��>?���kh)׿�.W�H~�_nTf�a�$n���v��#A��Ω^�HGn�P-<�l�̺�v� ��2�Ow��tR⚝���Txbܹ{��	�*q���%��(�z�e�O�*mL^�!D�d EA�N�?U���;�.RKh� A�2(���K��Ė��n��>�$�I�	�'n�ۿ�>�Vl��s�a6���ȵ�{�����r�9��52˥�C�ˀȅdh/��N��ՖR������۬/+�/7�7���)��?O�m̫>�%��k�Sڝ�ļ��A֢J��/�?�5��G��QT�H��Oo�%�ʎ��E���Ƶ�������e�.䎽�ՠW�	�R��h=`<G^s�.�
7̮󦳍c_�ȩ�+�S���c/��G5�����o����Llo�P�<�{�E>��HXA�o'�w��H3"iʎ`�[F+�7�yE�j��wc�I�O��ơ��&��	���Zл5�^��$�#�Ѓxʸt~C��G{�>qo�yp��XlG��QS��FF�yT�H��d<��*qԐ�@�UBN��%� :� -�Ya�槞ŚTɒÞh'v�~�H�*|De�*Vb��&��Ƨ�?��B�GGD�b�|��Y�s��Q�	�p���&��0�׋����=u��@�wrQ����oҚ��;+�u�W��m��)T[�F�N3���7�T�At�O�rǙ�A��Tʕ�f�D�b�	y��qm�s�L�T��7���+| s;�>�K�j�������Gw1�t<��ܧ2��ȕ��Suܔ�/:z��M{�`�M���3n����gl��3@n������*����8˜]�7��f��<��ˋ<:z6�w�Yxp���9Cd+��xA�P�F�=25;��2�p�ϜR ���g���70PA%�@딝S�;�I~��Ba�����
K`[5�1�a��v��[�'mx���\}��:N�(���W�����[�����+(��έֶd�+(�ޞ
.p^l~&lJ�4�Ͽ"h�k��T ��f�93p+_j����ڋ:��4�A��"�p6uBھ��&��7>�=r�0.zޣ���߁�'Y�3�~��G�R;�} a���Ж�c��H��G,�|�ќ��Ux��I'��!sC�Z٢9�m�W����M7����=��7�7�d�D<>Z���եZ�9��C��N=�>�d��;�[F���Pp7�U��g�4�s��-55����ӝ�IK"c쳱�f��1KC]���ۯ�k���=�
~'�5���8dF�[�H�H&�uK������i#3f����;�G�v_�m��漟�2�%�v��خ�Y��a�\õ�J�:AG��x)�n|�&Ң(���_SD����{ ���n���#J,���=����2)��j�y}YQ���7L�\�Q�:���ڡ�%C�l�Wl���Z`�������6�@��ک��/ƌa E���yrT�a�z��hi�0�$db	��1���j�Qb^N�`1U��j�pVoh����Y�kP*Νw͝�;��TDI3M{���-q�~.A94�K��X �W`-j�R@+�cg��i,3\J1c�F���\ۗEO��?��7�c��(_�#)��׾(y'Է�T&q�.�á��<� n��
]N����;���1C�[���W=#��T8�L�h�{s��5��	'd�[ڹ���t��N�H�G���Cj:�f}�.�c���>��EnP�0��W�DZ]�h��^2��<�����E�{F��7�5���*��D����̟�)���X��� "Uzz��d�[+�kQHaz=2��o�t���[�}WK��g9л��ϗ֤%tw[����*Rv0�W	���w���q��Im�EX�'���K,EI�I��-�,g&|�IL����gK6��귈������9�ŗE���~���qU���SkX�Ȋ���L��c�{'���2c���]�Muff>s��Z��?:�c$����D�k�{����&5�^�`��cm-A-ܴ�pY;&?t�n���Oeb�xWͶ�',��4�{A���'m� ��2�#ً-��Ts���=���#���.���f��䠬�Y�@�"m{���.ɴNcrZ�\y7eF����נ�nUh�mC2��5H��2��+ڄ ?�xXX�n*�k��-,�	zW��N�gS����`R.>��'SH��*
�.A��C͍ըrF������O�;B�J>@^@F{��������	?I�Y��_X~y%�1�ڥ�q�g:g�������k���'�����{���f>`���8D���\+}-�pX#���������ץd��Da�K�/�3e�5]<v��n�ɧ��`AT��j�"v`�B�U��7�z�5�4a(����x-;�h@T.}g�^��c�		Yv&�G�i۠\s8�'��s�Ā,w�J���僋�bh6�`��dT2z�̲��8�������{���VW��"WAi�n���|�g�w �GOt=�h��3w��xƞ���sH)_��6�T#rs�Xl�q'��ԙ����Y6�����dw�x�T���|��K�M�v$���ZC�����j�r�$2de�ԟ�����:["js�hW��}&�=�mX��_������z�{�ֆFo;R�h</2�B���d��zԨ�W\*�Iň#_�,�O�H��m�4��ƨ�
� ������P[S��y�<)�eiw�ց������`QWo��U$.��8fl�~�cK�,�1�<5�U�9Z�)n���wV*���Ch1zv&� �lQ�J� �[��x�<%gi0�NŻxv��F���BPX�S��ߪ{�U���>p66���=N�^��ƌa��徔�OL���	�%�q�+e9T9�w�ٛ]��[C�ߧ�!#{S�x����C���YIf�7�Ü{TH4Н�b�`�ڎ���3\ Dmg���
�J�kq�����~_?��6���=�K�K����2�O<a��8P����ga��b���M<D���h��UG2q�~�\̧���������:��a1+E�f��'xjLT���*���D�{`QcD�@j��Nn�Z�m�M&����\�n�Ror�o�������M+�s��&�A����ꌻIn�C;W
��,¸je^V'��X�ߙ��x@n�,��j�3x|�e����1Ō�,�>�s������`����Z�aow>R��H���S�U�h�p�V鐱���	?1
�g�)G�W"�^a�X�)6�i� \8�����OJ���/C�T?݃����~@Z4J�]w�]�D����z�!��x���RsƼ̧��aˡ&��<yѫ�#'��V�f��jE�M�9�Sŉ�yC��x�_7'�R��"�����"�@RN�����.�2!4tu�蹳�'�_�ԙ�8鈕�K��JX���l�RGD����%�ʑu��
.婴Js�n���Fl�<�LVX�^d:p?����='��<�-�qP�J�K(O��dk�H�e�>�����Q?�{�D��KD�ĻW%�@��J̭Z7Ǿذ��*E4:۬Ϯ�P��0���D~㷖Odʴ��Pz�$-	��.��n`�%��#e
^�5���[��RE�!�[$]-:�؂?�k��)�3�]�ѕ�qsXU����<�ϰ�q��ʸK�P��Nsʲ��*
��Ր�Y��ώ
`��5n�.B�PFI�o�ns��N>#twq*�*	���*KU���,��ژ,�s�bw�&ha�s�e%K<v�y]G�!jaV-cճ�?�]�}�ze�X�:sM���zg�t�~�}�&9���x�K^x��3�!�����8R�i[ՙ�Z�a&��b�C�zn���r	�@��t�UI���rUB��D"��I�\*~��h���IV�o����q(�Z�g����g��v��1��z�5!x�yY�ys�q�%��s	e(PX�R9�}Y���Z��w"7�ҡ�F7�����b�j�=���Kkv����wh3���� ��J����~Gm�c^[����A%��𳑢��� �I��;8K���{���X�$iL�Ĭ��!P�Zh4w#ιLҎ]����LS����>DE�PS����='��K�ˈ]�l?�s#1K9|k$�v)�d�G�NO{I�r.zR=� Os�� 7w�i���@]v#J�ci�C����҆����[k_���7���Ƌ=� �G^�,��f�-}:��fqQ*�ˢ��~�g�U(�L:��j����]�^+n�³���"K�b�i�k����h��W��B{����s��ܻ�[���tK�ܧ��%���"�a�����o}+G��,ΕY���d��@���k���گu���ȅO�VQ�Հ(������A��������Z��)h�z]�v�8Q�x�X�j�N�r������{�eë��U=	-�3��o���pLf�7R�o�2?�mHr�R�Ns�PF��xZ+t{^ZC�Љx��Qkc��I��n8��AD�jv��i��5]4S�d|����H)��RT{ݦa��]9V�mI��
�)���_!�8Ķ�f�J���ʴ�c�d����ZT��(<L�w���P���»LK(OdW�q�����R�̣��"����N�����BN�Nc"J�S��RMSc��y�̉���#����s��7XBu�d�n�.��?hҡͬ�/)�+S`N�ƈTp��������Ü���iRzo/,W�A�ڵ�Z����90��-R	�L����M���ك�x&Z�����#5H
��?
�J��K9$V_�����2�f���R7�	Yѡ�ъ��bh�Q8�e�����)��&i�̠Ϩ~��!xU�s7s�L����9x�Ɨ��--�N3�'�0,��C7&�|�� y���Q���Y_�`��jx�Y�;�ț��ώ����8�ᯒ�~�_�/\MC�TA\Z��=�i����M�8��pS���$T8���M����`4AMc����YRK�����x��<�>������m�-�ǂ�\��LԹ}��O��S2mEte� Ϛt�P�� V� J7����#�1���{��f"�g���!0�0:6�/?�q�]�*l��pD��w"��NI�)=��!R㦘r>�C����1�Z�C��*Ɨ�����q�>��
�{N��������9^��\^.�N���)ǃ��!l=�-��h����E�&F��3f������a!H�FT�J��k�Շ?�I�DoL����:��B�-&�l���>d?;74��T|��g�����\����+�?GM��re��ީ����m:/� �]�3pF���~>�����U��J(@�{�p�C8(aOKi5�U4!XKeuc'e�g����"�ܗK3Lq��s8L�8?��g��J,G�-$6�!NX���NP�03�$쇇��k_����k@�[�?/����ş�����NIx��P9m�D����h0�>·͖ޗ�0�Gf�a,7G�bR�%��@���f['�������A&�%�+��A+OZνc[�"��"� y�r�"�Q~j�<�2��|Y�`�7N���s��z}e-7�gz�E2H�xNN���EŌ�@^l7�\�ɪ*��%r�T�Q���V�����u�Q�-ʵS���<.1�̮> ��T8?j��F�e�!��;�TG^Tz�8$��<�A��T�VY�du
� �y��`���RU�/��%�����W���} ��Lɗ���R)>w��l)�68����.>uG��ŀrI!&?��w��׷?I����-�<|�9ZȈB����$E\דraU`ۛF�')�߆mo�o�N�-+Cwu,�da�Q@�<T�^�#�f8���!Dw���_���mҺ���/�R�i�1ERB��젻VV"����Yn{R�c��� ��}t�1����'ҫrVc�7�����1�Ҟ�Ȝ�7G����龣�L�,����"l�/��3|/L�I�?�ǂ��
�`#�7�b+φ3
6�״����k �>���Mg�뜽�Rv�}o���h�u ;����5��������4�ؿ�J�O��#IN�����m�F��!锯��=]�&�z��R���%�����r���¯�m�q9{x��A:����"CRcEw�Pe�D� *Z�ݹƳZ��%��
��jtY��W�6�ա�-F�����o��E�p��Ĳ�v��������8���ul�:1!R-�d ������2��X���G  g' � &%p|\�y�Ã��q�çT���9����ݦq%�-A�ɋ��lq�ئ�f���xE������9���2��CЂֹL*cQ�ٔL���vb�ڍz� f3f���6y�LFb�	�p�h،W�T�D��/�{v��b�!��*����-K@��8���4�A����',|UI���5�/)y������VW|qd-:d�w�
�_o�G�)�G���I�\���1ַ5�m�1�����@'k�������6���
�S%Xod���WF��;�G��y��������[�*����
.K����)���N��fw
�H)�e�p��#���	I�6�ڽ�Jna:O����tlI�x�yuo����AҀ�w�_|�.�'�=�� ���M* ��8D�G6XhJ(&Ǖp��(���E���k�IY�0ss�7©r�-#��P�����>�53�^)�]�2@YuC�옝�Ez,?pN׆�r ؒ� ��[�'w����jR��/����;�d��BF��|�2�����,=�@�TŴ�~3o�۫?�n2�)�U��NR�@Y��X�$���	"�M�>�(�-1�����a�c�"�ޞ�Ul����Q�2*��2�_�i"�Ò=�����B�J��e�;� ΂��D��XA*� ��s����+gE �Y�H's�ܙXz���O��.�0q5*%r7[k渳���'����)�P�
��r9��j�`�U�\P9.Kv�F� 2��J><�K�$�֐2���Aߒ�O]2(l�|�\l�S*�`�u�1P��4:'p�23�N����K��f�
tv�Hm�쥇���ͭ���M�FO��x�]΋yP��D��p�j7�rf ������RXL:z�qb�<��&��V������=3U/��)2%7��1H��s�܇"!b�P�t��u�k��2����w6�((���IW���2�Zs7d�������{��[On�6�+H��Pz#.vEJY���I�=� p���,ֿ�^u@����<�q��b��?`�E�.�}���A��d��z����1W��L��C�K�6�ǧ�	��3��q��3l�eԸǞTh��.i�c��YP��8�����&��:��JȜ�Ǌ�^������s"�ݿ3�u@�	��U*j�vl�� <���Ƨ��ʺ~��9@wP����s4��s���/h@�prW�K�w�f8��M��V��������+�Ұͪ�ʿ��xS������2Tt����#�\�:�yGf�gs�6_�ػ�g���W���^l20�-��� �9?#��f�%����&�m�^�ⅻ"�Zq�E�.c� Bd����5��d��[��x@=��}��/��� q�:eY�ǹ^�y������D��d`\[������D����%�M�@��z��.��Q>k�L��󵚘�G~�I�Arbpy_�+� ?�4@�	ά�O��(� ������I��\n�f�.�b
Ǐg���R�J-��+خN����&����)S�ٗQ&W�������1�V]�2���L|�d�T*r�!��a�����3���u�U�3}�W���lؓ��#7N��Da��E�u�(Wx�s���{�0���H�
`%9`��=<�Ox��M�U�3���r�=#YKz�o�r���sӥ�8Hd�.r\���z ���~����,4�וM�Y�vḴR�?� ����G8��s�Z	*K7�SI�;�咒�z���'W;!��1��	є�&�$��-�^H_v��-��%ۺuc��ױ�=�o��s
�ޱV53�5��7�U Y��"H|.��2:n�"t�*��J��Oh�_�X����%��Jp�b5φ�Va�IgE�e�3����۷�}MG��D�ǘB��^��v��Q������Ïq�����	+��5����]X@�
^��Ƨ���h��F���Q��rn{���t�z��v5b������If�.�������%�{���P�F�^l�<��	7�xɹ9]�yՙ�J�M4w.Z���w<wyOq��"�d6�?!o��ķ��I����{9rG��9)M-��-�geZXѨ�cۀ�>��J3\�2~!иG�H��� e��ù�?���/0��m������X��w�9壦-'��>q3+��,pс�ߑ��$Rh�.�+>2�\[P����h�	�����ad���3�lw�����/Է����D����L��^�#U֌XEMhO���vF���Ǩ>���|�#�/ߧ߷�h�͎H��Ե�m�g�\n\�j�A�u[�<�`^[:p� J��!�������n��[���0��1���/7�_^�_>`�2�P\Vl$P����W�1����Xa��:�HO�R�]� !�G�j��b)Io�t~�Z��,��9'�S�77����6( ��\�k�O�:ob��p�t���b�^ޔ��D=i�|��</P��a��AnD�)�3Ŕ��`�Rµ��4��}&�������I�'��)��vu�5��\�$����wW=fD��bB��lP�M7�gT���.FCe�E�"G @VϜ'q52�f�͗2��Qz�1�	��W�.��F �vu���Zݱ�׳A�kLm��\@��Ε��U`�=��K��(��%����)wHB�ZcVɸ*͵x���
ӯ%mK^1>#�RS�������i��,��bS����PϘC�x�����	�»sY]|JD���&���Z�^r��hՆQ�x����?�qL�T�,��0�3�o��B����,��V���-nid����V-��c�
9��kNj�г�]]���L��.�y�[��썸m�$�P��}6�� ƪP BR!kj2 �==�p�bx땯!|U�l���r�#�p���'�5l�C��}R�`�,`S.�=��S��	�4�t�
�ː�+��-��|a���5L�	iT�+��J�1��o�j���_U܇��7A���������`Gr!�ly�K�i���d��F�ϴ�L�Q�#G~���[�NȶapT��[�]�2����#��rűP%�n����R�߿�e�����D����gkZ�B~3��G�m��8��V3}���X�+�Z���1���O�5�w'#�$���蔄ް}=�|����<4s���m�1��|��H�lmc�/ƉV�Nο�5�����Q���8]7N��,��l������ v<1%�oJaR�U��Dv��sB��+{�G4�j��k�nU�.ln}iz��>\�}lߘ��<��/�*�Ф\D�5�����cd������y/�Kht�=��F��Ǭ��A�JتL<Јt*}8s�
�.G	�ӗ-�{Ĝ�+^D��pW�������@tŦVY��d�)Q��e�`&���������4��"��v� >�==�����0�m���s!��� �鎭'��Q*<F#��=�����!gȸ��vE���+���3�3�iJ������R��b�yf��!��𧭊��`����]�bb����>)�x_�9�N�3bO�����ɰlf#9#A�~�L��q �c2���jB+|!2ā�{�V�-tMi�E��]d-!�zT/9ݳB���ˬ�\}c�&�rR.�J���3�%�X��a� ����NWt�WS �K��x���##����+�`���l���Ʃ9�=�v�5B��P��<C��]e�R��׽6،��ֈ�7��d�>�"Ƚ{Ǹ��u��w�b�2���
 ϊ\c-�#�{��O���RE#�U9i�l'��%R�-"����f��ǥ���M;��B��%�>/i����Z��J��4�}��=\#�$�U{U�
�f��wɪ*?u2�+���1�Z/>��,���s1��+zp�?xd$�X�Ae˓e�j�J�L�Oi��il��]���|K�fX���OҌ7 ��x{�d$�ѩ���-c®{�Dpi�F%�#M�Ÿ�A7��d�iG��*�V�E��Up2������>���8!EԹ㷙�;�-/�ɸms���xc���^I�^'M��c�3y�X⹱�)v�g���(�#Q�[�?�_�c�R$ac��gD�����#GKY��x���C� �kW�V�9A��^2�bsVoM��׌���f>�����R���h�4Z�^db����h<��l�m��QfʉNX�߮��ls~�]2pJ�=�˕!�p�_v��<����,�H�mu���b�ga����̩�)fW�=ē���%����s�lx�v}�w��
���B������H�7���d5����6sݱ[H���`q�k�3��ߖ iç��}*�~*9ݡx>�w[�(I%�02��}�����aw�ݽ[7�a�@�O��gďj�'g�R���7�P
C����1F��.��4˝��[o� �(��EZ$�& ���ԓ��Ɵ�~�s}<(M	��I}�t��QN��0'�B:��2�Pd'�VX��5��Ç~3F���mix��KX�p�V�R�w
�tF����'�{?X���F�s2Hl�� �k�@w/S�=��K{�D�ף�3iʑY {U�V\�e^CF���O�
di9�Z�c>�+���q�c�Pq�3ˏ����ƞOߐ� 	��`��MX׿�%�1����������Ħt%�B��;%.9��N�Jr5�pT����k��l
g�=�MS��9�6�n��k+B�o�#��!����js�&(����*n��[!���fo��_m>���>3?�w��F]Ku��j2".�'�H�B��i�L�����0�����հJ�ȌZ���jr��I�Pqn_��+���k�,h�[��\�+�	1�9G�w|��h�����^���R[7��h�L��#9��gFl�[J���ֵ�,�|��j��,���1)u�pK�8����hvI�=�Y�1��"��2]�/֜�q�Y�c�NG	$��RG���/�[���b��W�/F�RD���v���w����P�5�ו/nwC�e��������]c�ayTs���Ć�@�ԆB�ۥ<F�nox����Y�b
����B�{�_94M�.V~��hv�ޙt��ٰݖ��w��TLd�`��nތP����ʯt��VO���i�'�F.�Gp���tU���J�[��N�f���P�mDM ^]9�J�1�T@S���J],�g�������\��y�%�+�F)Z8�c���V��0i+,[G��D ط�f}~�a��P�����G�OQ�u��n�2#,e��Պ� ���	�]�w���2�3���A2�EOUE��T/+2=�Z��@�zҀ�Rw#��c� ���BQ�JF�~�"qUQ"H�"-kO���Ӏb���wG�l/}����b;N~�Ӕ$h�$)���V��/g�����I�d�Z� V!,���1G�߉O��^���7W�t���D��l���U���SA�B�(����ȷtB��`"/
��Ze�����S"�f֌BsY9
J�/|Y�_�I,Uv��dB�pJh�br���$~�j���}�2];w��Z��JsgXX�}�A|�UU<�P��E���ņ�ˉ��� �o�X9p�l��˻g��U�n�������q�_��s�	�A�/>eF��I�5�cAT��4�T��V3�k$j���!�'�܅�<x$�Y��i��w�L��wg��$�ƺFtR��P2�H�w�����P�Ԭ�"s�E��B9^`�X^Bl0[ Ϸ 	X���fRqX�u�4��	���L�\?�Fe���|��Lr�7����<�V�1?;-��@G�:D�7�؇�v�V5~d���ѻ^��j�P1���C�� "*�}�	�)I��.(BC�w�R2��n|�@�1��
�$�RWU�%
"�����2�Ч��1���6+O���ty���z�J~��c�S^��E��Pנ�ZX��*&]��R�)_�������� �w1X�#C��I��L�q��_����uMX0+�X���;Yƶ�hU8N�P�KyK&��:��1U_�/k��"F�	���
{k�PħO����0�tsW�{��G��((�4ϱ	�|��B�_�ϨW��Ĩ2�Z���O�^��	"#ܚ$4�oJ � �6G��<���K��VG2�ϐ�\���{�n����>לu���d*����T�j��Nj7Xe����-)A���.�������v���9�&���0���e��X�Q%%�\4�ۋ�5���X��R&��h�D�/�V�#�2V��hM-=b�ec�c��5���ꦃ|��s}��O��X�~���F�%~����<��с��9ʥ�M�x��G�M�;ݭ��V����H]�Y�,�%D=�g�K�<,��g�"�tU�PcҸ��Vw#��y`Fׄf�1A��yxt�ўP�F`�14�5Ę��$u� ���^V2t0�V����<ѣQ�]�y��"��4Dpe#ʍ��^0Y�Sլ�)�ZO�:4���c���C��5]}��aU2{n�[<3-��&a5S�3I�h%���6�H���wA�S���dxǣ�ۯՖ��2�O -����h���;�{+N�|�u]���	���j��� �WE뿿#%�&��^�%2��r֞��Z�6E����C�\�Q"�>��mQ@PC6��"Ke��4�sI&�Je~���H�|��x��t�p� �_��g���+q��D_ٶ
2�f4�T�����W꼏�<�cr���5 :BTKF2����oAC�i�'�ח�L��M2@�o�D��=�m�Q\R�&�������E���gH
w^�u�C���b,�N��h�����Na[����gs�����Ao>�rF;l��c��̝���L���� ��
�dJKXgi��d�S}]�H2�z�ƻ�&X ˑ)t7ft7R*�#�ڡIxE�)����ɸ���K��g�g铜��V�rm4�.�ޔ@��e�J���\@i�T�-�Q/�A9��rkuI��>�b#��q��ЍNX5�I{���\E��2d�č`_�\�c+���b�uc/���]�=I�����Z����=�#6�+��_��o&2¹'W�^�5H�h(Tj�g 	N]V�"�C��iZ���/�n�ʅ��z3Jx`� <p-���
R� b����%���i>'�g�a�9E��~�?����d�߈�lO&KN�3��S�~V��U�R�Ҡ� de�_��
xr�U�u�x�\1:�O��*��َG9�H,؋U�>�Yjr_?�nG���>{��S��K<���`UO\����tɀ�����ze=ޫ+�H����C^�w�O��F��o�����!�= B���=��^�A7R��m8��l�]�ķq����ZJ����Cħ�1���qy��4>��83-��񯅺����q��p"�m��-��8�a�\�:�Ӭ�i� =q ʥ�T!���_!$��_�r!o+�s�����M�?�w�Q5H콅2��'	W���E�/����H�C��U�R��g��,\��$r�{N_JS	y�����9����7#H��{���I�`s����B�[�3��u�ɦ���)Gwp��7}�OR��a�z��v]��6��~��I�f�c[VM�r8�  �U")�\�:�U�Օ����2�� ��-B�z��D��l�����i9��q��M0^�h&$�����e@��P1d�=��{ٝnx�*��u⋄�=�ٷ<K�OK��������)�V��y�%C��#�y\sGq�(ӻ����&I�F�Ǽ����X���/�?�"���p���*|EM�tB����_>��z�V�c,��zz�ِ��������Q:�̷�x�T9�U�|GT��W���T��� O�Im��)y���}
 n�0�1�n`�!�NT�Z���Ugb��.��qn6�>��'_�lS K�@�=�A6r-�-[;�W�^+�
��� u ̂���4��6����!o(�rD7��"��7�eZ�k�B	8U�3��U+�>x����dS��/b�\�R̂nN˖&�7�n�⓮��6�r�� %�|�DD3���]rF����
x��	�����,�tE��B��2�P�'���y�}�'6�\M�)D��7S=k�L�/a#���tӴ��\쎕�i-1�1��@��o��0J]�m5G��=�U�Q
�t�z����ԏ	���hz�5��k�F��C�{Q�3'���-?.ReMɚ�g�d�O�`&���IT�62e$��x{ߐz�[<i��;M"�'�>��f�Z�4�`����=���62EG�۠xc���G������/d�MN�{L�RIV�w�i1���	 '�7�����A�'c`.��$#S=�C(�FdG��B�tW�3�1=`�?Z�Bl"-�Y[E����R$ˢ~Q|e�|x*�h9���F��*��M鏕�<a�0�t�����|�0�ȳ�n7��!��}!Й/�R��t������s�b��b �-T��U3�AuZ*��l�]ClЮ�"X�L��Qx���$���?�a��ֶe�J4���䡳�ѺӛY2��@��q�^F��g�.���c�F(+�:b��"������F�"� ����e��Qr�#�J}��yr�]��%C3�׌�2��M���/�)�tTh�I�\�fBR�3� ްuM���`�#��+*�Š�ޏ�����ޒ-R��NH0$������Z�o^���� ����#���|���.�C�kP)�)��*|#C<���7qe�%���N�ԭ�@��_z*|�xF
�Qt��PjD�N�X���]�r-�C��W��=��7˯�� ��׬��OV�X���U�qv�D�������W�(S���
I4}@�Yk�AR��욢�bzp�Ոd�����V]o����NQ�o�Ą�.!	��kE$0}�=��l�zsW��p�0Tp{��ls>r^t,�8yw���C1gϾ��}؆��S�a��I~�WZ'��z1Ƚ)�KϬЦ����ȷ��ox.]��+�3��ߠ���P���{`YQ���Wu����7��j@�`��������|n/gY���[����LUG1U�i�LI�Nd�?a�"�|����,]�XjW�F���uG�d�¿�n�c�"������D���B�0�gE��z�N�j�e[�X��y]v�Íj.h.��G$u��2�aDm��`�H˙��NQ��5���K�8}u>n��4�'.���-`�H)b.����0������P�	�s���20aWp�&����Y��T�A�^}{Nc+gV���(�r�n�����_��w�0���L����k��~���Éo%D �<i�����	n%bp&�_�7�@tA���M�0�L"9�^2�#1�<i%��^H��^��sUIcц�!FP��	�󜏯�P�P���i�'�F">�BԪ��7�aB{ڽ�>� ������e\UL\!���ʙ�s�QB�Z���fʗJ9����Q|u�
�ÍX�$�B۴r�t7o�u]������<���sw���fJf+�)(��*_����t��=�b�z�c��"�l��ED�s�B�K+J^9��m��*еk�q:u��D�٩�'�(���8�F*�3�s=�Z��<��8��%��8�m��E�S�NFC]u�&5�z�	�iu^ìA���[q��<��;T�z�K��帕��G�ݗ��%fɚ�������kJ����8Z	d�&���}��j[���k<+��[�!r��𐚺"����ox��E4�g��:Z0��zT��>��T�����R3�����vS�m��7B#�%Wލw��p�㜲˵Q��w}�p5���1"�Z]� �(VA��0��"j.fVt���8G���q�鏆�ƴ�1���Y�@��%B�;�gI�?��u����+.�2�Ih��YS���C�cA�9��R�n�O ���T�[��ן ah�<��K�X���h �����ds�3f�c�OA��ې'G�-% ��I���x�T��2=mr��n�L�?,Ae�;^�yC��&��<�|j~��X
�v�����w�ㆡ�g�k�:��O,�߄ͣ�+1�Wi #2���7�pu��7S,�8o�F��H��2��L��eCb�t4�Ě�<��ٽ��Z��Y���
�lsP���K�0[�X��@��G�\�5u�$�,Fˣ�Z:�L�݊�-]��DQ�b�����t6�/:8�;����bz@�j��A`���i�:>�M!�RC�P6ŧقY�!�>��῁�ܞ�h��s���A��Nԍ>!�bP�~���'�LN�;���3�	
z-n����B8�G�J;��K�w�9;`{�2�"�R�-=�v�!��妿��7/�[��p�dN��60�gs��Y���o�z��\�
k*���0� _��B/g_�;�]�8.8��2P���a#I�JV�Ao��:fZ��������Q��1�lz��v?q�t$U��\����z��]]#��(���z
�9]e Uhk���M�9�(H��-��<WXt���%L��� ���<Y:w�x�վ%�q�p�5=ݡ���|Í�\ZU9$� ���%{L�x��M�&�����g�>�טϹ�[��D� d�Bp�t
�_/���K,ηyt��gޕ�$P����M��S������
U��e��@9HkB4rO(J��(jo�C���̻j��X雳�"�R��:F��j�#��`��y���A�t�{c+�(�����/֕��t�.�F,���p���(��]�����~uO(��`��~m��|Yu(�l~E�^��-�((���q_����Z�+���*�=ȇv�����H,����H�A��$�%���mE�Q�U�˗ճ��-�k	EfHvM��q,���RR�ip�2龝���p���������")����wJ��բo��^��A�řL&�6l,H�5��bn��㮗�dC��Y�qC<r�<�E�5�I|x|$�G��� ��k#�k�Hp�,��٩AA�e<״N���D�G����sb�4�*�^1���;�wO�W�3��	�e�"����G��%�UY�p4����P��\�>�T�����P9����mT�0���h�,B\��׌6�27c�����F+�\6��-#s��9�HK$GܮƵ���uMA��ʱ+k���D�%��9"3���Hd�;n���`��ʧ�tI�!��M_Ā�t�HL�v��Հ����A��  7����ɎM�,��
E�p�J炘NaK�k��wa*���N�
?�#Z��cda��A�d;Zr��d�5FlY�Y�Մ@x��	�V����Kw;|Ta�(���:���(K��A;�icH�Z��㵤��,��a�z&������pvn��q��'m�G�K�M���`_%����͵;�|?�U�r��YZ�+v����в
1hL��1�5s��? z�6�~�`�o�e,��ؖڽ�#���֥*���'t�-�<:����. t�r~�X��t鰝�'��b�-ލ �� �Y�K���c��r�q�3����2'+.:���z͵ ���f޼��r�ydc�n��k��!�P�4D����Jpch+����T��qI�o�M�"|�Y����`�iDۣ���_��t�Ʌ8�wӤ	��k����9�_A=�\�DйI����BO����RFP�(���Q��n-�4�Yfy
S��%�j�Pi+&=��w~R�B���,3q���������ɑ�I��KX������x`����`�:�IM!;�#�
K��a�?e�;B��s�:�5z�_�""N)�FCt���u�O�Bjtl�!yW�H8Kb���p��1܄���+�G!�!�:�>��'şd+��٪�IPߜ�@y��fg�Q0I�� ȳA[Ic�>#��lr%3ڶ��,$���?�1�(��N�^i����VG�
AӃ����*���`3(��-��ӆ鯋�؎�^T���!�I��0B��r`��%/-\9k[!����W��4V�0y\�l%R&���7��4���^�� �w<�e�՚�I��zp��pp�Rj7�C��)��L>ԥ)'�f���J�(P���$X5�6�7n��E���tEY�����!�T0����|Gw��������A��t���K��
W��|����7���5L"Ñ	�������!���!�c$�����Q���v����x��#���U1q���w=��T�U�R�VE�Pg�����,����j�����I1�;zKM}},k×]`��7�:쇠����~�V����<P|��|B&��[M�6�qsu���S�0� 1��i��/�8kª��h�:LQ��r�T����n��X:l�e��+�7����(���T=2|=��P��-�{�=�=��4�j"�^��[eI�S��������O��XБ���
�3�����O~P����������ﻬ��l(�ľ�$g�˱lM�Q�aV�	r�ۇ�K������-�f��э&i�V#��-�&HG�CV����*����Bk%����[n
F��]'�8���o���{�I�iy�B=�P�f�`��tn�,.��)<��3��ɠ�f:]@��z������iʗ��zNt��k>?��v����h�|�)��)V�7��٧�t�����&BE����gb�Մ�`G�E<Tp� ��(m��l)0F�ew��#��=BC��X7�gr���f���;o��r�(k[ϙ�3{������"�-�RG�9oU���<'��N�F��(*	S�a�1�����Y������ߑ�%�.��5)�7���ɀ�E��p����\�a�^<	]���k��ޯ��@�L~���1��0#�#���+�0�T�u���73{��Z+TB���i��v��{�_���G}���@��M�%�a=S���0��]��A]�;���Ws�uk��5hȷÅ?���?/��g����~6�K�L�@A��VxU�f�D4��wL{��ς=�c;�P��Laóͽ�I�{M�c�u�+����;��c��(�u��AqSa�٬0�mi�[�f��)+[���[����XB謹D�!/|��������e�{V]`��|�`nI�Ŵ��*8��`�ِV��/��')�Z��v�g��������K��V^=��6���[߷!��~��y<�����
��]�҇���#��0��^���q�O�y����̭<��>��]Ջd�h�ph��h1�J��z���qM�Xi�� e�5������F�h$2X?d��t6��!%���J� G��Pْ�����İzn��Bk��`�&�[�z����h�9c�2���dppB�Y��މ�xp6��rK���%KZ��lα��[����مs4�����5���,���\��"�%,�S�'.�N����m��q��F������Y���;��!*x0��,F�50�*���Į6���U�d
��8�h�'Pz9������l?�D;��~�2��2Oxg1�l��o>��k;��S���n'*J�v��OP7'����G�~�'�X� �q�#Gs<g3R̢������ �P�>=�k:Y�:l��M�2-D�U��Η��$�M,	�z��u�"1�ZHyx���A�\�Je8���s.͒(�-�� �����g��;q���Uy����^�oC=�ϫh����L7���Օ4N����E��|I��c9���Qs�Tm�O=r06�K5�b���Ϣt\��%L��s �)�z��;�閑9�r�|�=�H�匁��i�3:r��eH ��a�&?��Pa�C���� Sr9*���n�L�%r:w�h�	�#1�ъ��ZQ)`��i}Fr�[�o���2`)���-��b�*}��d*I��"�1�&��ŮѠdJ(QU�t,����5�.l������T��X	@a�iJ��!M�LûU��Xi5d+����l�Y� �u�4�LdC��Z�gc+��Z	��?�驨L�Աg�DR�5A�z�t�Z������J���x�mz/���Co�ڠ�I�۟���z�E�ǻ����	Bb�&�+��~R���~��ChMpd��Rx/:�\4���1�)�t��A�8��Wy�J�{þ��Y<N���cQ4V� ��q=�(���� (�0A{�ϵL�l��i�oTƳ�ӝ�	������	�(WAMr�i���5F���
U�y��|��+
 V\��$>Ź�A�m����< �������F`N��c{�hӫ�u2������Z��SF�%7����tn[%�"N+ �x�����f��˛hڀ�d�97��Sx�?�����)��H�5,^a�����Ku;L�p{�;jo��(&�:Xiȅ�z�c.]���$��F=�'�(g TjQq3���ƕԲ�������q�6<HAMKNm"���j���#�˝��	��)g�+��v���#Y�z4�]������h'R_�B���S�O|9�8�n��K(}�U`7?��JoϨ2|AEj�H�\^��n�+c�$ۮ�rO۞��6�{L�-uc�	���gy^�ĤU_���:�%9x�J�mjN��%�_s�jM�6��J��kc��L�n��=K��oqO>�Q�/�s�p B;���'gX�!�~,�t��|t�1x=eMh��N�䲝*���K���73�z�vkro:I�Bi��-,>�O��Q��h�	 �F�7�y��P����4Jfx����w1�ъr�����'��)	͑����i݇eZ`�,j�Aʃ��`'�ey;Pnv)�!j��`}NZ븓s��-@���_��+gu3��,�z�����/r�TG)+?�0#'����K6�k��3$lo��WCAN;+��ϔ'.����]mPsT5i6��Q�!�K�U��� :�L�U��q��U��{U�W��� %�LB��Q8�mc:����&�"���P�LeP��7 �j��������#�;Q���5a�t��bshOZ6l��c�P=
�Q�ϭo�u�m��_���)d0�I��ϿH�n����u�,�ODaI.�X�3�E��蒳P���%�K����r���9���?������'}��R>a�
u��)�PG��A��,�V�(�r�tX���[�f�=
!�I&j����1Io����1^�tł����CI�+��P�LG�y���^��\���x��N`Sc�~+"&��G�|B�ý�u��lF�`{�,*&.�}�@b�C��Yܱ��?
��k��|�!iu��~�hŗ���jsj@(�ͮ�A��ۗ���9~1��e)A��g�7��"K2�g�x	*~��#Y��C���mԴ�&I�@~ml��N�3��1 ډ�Q��L�^�+�C���+sb��H24���HU�_I80Q/��K6�o��%1��S"C^�'gH����� �+"DkRݘUg�_�%0����<�Cw��U�%L���ث�s����c�ڌ��+2<�ʶ��"��&��v��r��6��
�N�����3�P�^�e����%��j���a�a�.��)Y�၃m��m3Zn�%�\E�jN?,���Z�z�Q��q��ү���W�N-)I`�cyf;���6F#g3����+�N0��갨&�	�y	�DޱK��\�L-�B+My�� �y�M�U�1BΜ��ɝ�U}�C{�cB�T|��c�\AW�]Y9]#�*�A'�
��<����V����
�b�Z��F��I3����,����`V��zg���%��j.�ӞR�
Mv�'ɺ��"�[T�iu��?�I���,���/x�wXd�Y��##��O�}��A�d�p|�+�E��ܚ�Yr�N����.�uY`]`W��Դ�I�K�Zn�޽�V���\�ȧ�,��֏źcV�1ݗ����H�.�Ɩ��W1��-�=o�wc�w��ʷ#8�UFӿQ,`���J ��9`w�&�qʧ̽�B
6��eYL�b����V���zћ�^��J����j��^��5��W�/~��VJ~�h�=�{3g`�C�W0|��-�R5�V��Jua�r��z �@3vo��nG�E�p)�j��� &��cz�Cx\��L(��|�~JY�=у�'���v�����uH��iE	�?�M(r��J���v�<��J�E�d��ɍN�<h��_H�q�$�h�x���/v�Rd�K_��ѢO�,����������������!Vh�-W��Z�L���W�^���>���ug��	�t���fvV�T�@��� ��H1
��X��;�2�2IF\.�Ɇ����e=nT�t�u�J׎k�MA �Y}�c�t���"��V�$�R���<�9�Q����n�M:w�k;�[S6 ���уW���1ɳ�G�;n({��^Z�E��|֔`mLp�V�{�g�W&���g�!
���dV	U�S�CW�����y=��;���*d7gbKr�!���7��4�N^|-����u���_��l;KP!u#Бg(Ia� /���_ի��6�)[H�M�F�PEG�bD�7۵�<���S|�����c�f�zٸ�)�0ε�n g��L?��7>�����i���͚��^Y�I��h�Zznj���6w����V?�'��1�G���>�f;TP���,�����9�����Яv�-������B�fJ3U3�$/��U�P��Ǔ:I�˧��P}����E�A>�ÏT~7���AI����,p;h�e�3U/�;�	���=Dv�DTG+�y��TV���8�S)���ZC|���4D`�����A>yU=ŧ�w�����- �-v*gi��b�nF90L���T;)7�{���O��D����G�\(ЦǄ)m���[9^q�4�p9�_�,�<�G>�����H��ߝ�T���VBu,_ARL�X"Ȩ,U��'���R��4������Z���6�>���v�§P^�5�9m��oc��ē�"+�����P_vE>���q7�]�����[2a-?�!�ME�7�ڷw1O�_���0�ފ�l�6V^�CU5R�?y"���yg�������c���� �?�2|U�X	�U �`-ǂ�dk�З����"����ޒEѵ
�
�-5.Wf��~��`�p�Ъ�a�4�(sқ�R�]-$�u<̖���Ж,t;S9[8�w֫�w7%�$��G̲v �u>���M�`;�l/	m��&�Gj�4�^�z�����^p�(U��Ѫ�����;���y���v	��{��/�/]�"�����wt�|��D�q쿰��h!Ƕ°���Dl��m9iHA'E�XO�cd$O*>h�-�5"4�֪��-5�~�\o0�f��J�24\�
{\)}�a�u��G�x浥(�Ţ��������T@2���(*���͛���J:|�x8O­�6���|��tH����]��d����\�&��q ��t'V�}T�����oZk7��J�	���<��!-Bz�*7j�gvs�טF�<؍___ G+���k������&��ɲa���N��]���O��ݖ�'&���2[/� �l?�MY~���lX?��݃R����ܧ�BT�p��$�wƆ���\2�CI����SNG!�*�$��Q�=se��s.��Ė/Pj�?j�KsU�S���B�٢3�yK�r�oBT��V�RP%����p�E�	�\��|��^��+:a��Ub���B.+��m���?4��������Y��f-D$������M_�=��"2�(�rGۗ	��،��CE�>~Œq�������s���j�(������g}"��	��Z��nr2h�#Y�AK�P���yܓ>M�/Tc#?����kYw�Oqq�~����/D���%�;#L���7�gM�=H���"���)μ�T~~� =Dg9r���^G�"z`��9|�LF�C�|Dg/�v���{�� Mg�&0�E��W�:�r�`��y�bX�-�2*�ē��}��C�e��%��>��Ut��d��������T�����Z��>��-�ge�����~��dena��n�����f�K���"�$���Jtz<�A��Ѣw�4�ӓy�>��Ф-HJR�UЊ�Z������O�䀂��EH���2��kO!%��A�4 O�}O��Q�Ovi�����_���ĕ���N����+<�#F		�J_����(�c$�.�3Yg�eF������g���x:�1�X#i��KaJo4U1)LG�K��B�+�E?��c���Z�=��ZP�.������Li_ʧ,SMN1M���M�y�8�\�T,�	T*D!콷I�)�ƫ9�ni ��%��p!�����u���Y�؟�K0�`_ApS�Д�@~e��MQ��n���Z�"rd�*�2����ڋ]r����r����q�����Y"QMN���M0����q#X���j(�e�檡_z��J��bxEE��6[���8�=;��!]�9X�i��R�-�"���<c
S�����_p�l>�8���j�qD�ܲ�"���K�:�m�����R�����0�w�&��h����h�c�^,�E�+@w	��
h�]�A9�Q�8�^���@�t�*!1�5 �-�f�BE�K��bHw�q�_��[ͫ�[k71>{uN���@��CUX��߃ܦ���A��fj���[�D�+�o`�La�ƚ���E1<��D藙�A�'�>����C�}��Ys)[:p|��L�P�� }��	�ۦ|I,9bޱ����ܘZ5�t���p���,qx��� �k�P���[2��S�=���iu��H� ��B$���STL>k.��XF6��O��:��39�%���'ɾ����?M�5��~:�$.��s��Jc�ďU�7�'���<
�AYtm��B�1�pR���G��M�æ*h��I�f+�#w's����A����CϪ��,M��x����2	8�9n�UE�Y���P���y�^,+�*w�����a���F�s���L�`@(�'z������OH)9VD�}@qԕ�y��e2sB�д���`��S)N�@$~��x�=%�H�U�x���]�A���K�2�i��HI��1�U}��%q6�"�?�;ց�0�����|����q����H�_�ƺ����ùd���Aa��Ƽjd����
�s{�Bx��GwB�t��#5R�1�����h��r��d Sƺ�>C����*ZJD��nS�j[��Qǋ,`�Ű�vE�h� �+r6�����;bJ|���dJ�=l��p�W~�N+Q�/3S-�!�ڰ0�t��uTdN��A1q�G\�3���`��3ep��%�=.ů���gߚ�RYCv�K����_�F��hA�A�q��e����LT���p��|8)9��0H����5�$�YG]�X�IR���S�o�k������Uf���ؐem�·��-�U���^����״a?rޝ�-q�e��>>���V���pM�{��i��Y�l�ఴ �z&���hǖ�|1?�qV���^'m���+3��ܛ�K5�T�ݖ1�y�RiJrF��L\�xFaAw���!*��r"/���V�2G�+hi�H�>��G�
'���0"�#�Jlz��bI��1tnњ�Ϧ�܅���YFѻG[�xn"���f"�pn��?H���*��4�*�*��{_����]�|�ֆߺh��v��@�{�I���܏��KVe��� 9y7���1�����uu�P;*!�#FO��C`����t�%ƐN.�%��XR��]����w�����>e3�,����R���~�Z�So?�+�0�0Z�A��Lp߰����G�󥶞��VR��G1���l/��v0�W2��J�e�%�F`ql���2Gj�j�^�K�[WHȽ&���Ԗ3A�.��b�$���V�3!
�P��d���+*�	8)�]�!�멍� �O��9Hܘ�����ܚ�y��#M<�. ��z����=MgFY�e�H��)����vM$x|R�OF�p�Ug��V�����%�`��&�>�LR�Tm��.�2 S���Y��x�����_}
���!zp���ihN�R�<ܷp�?g�D|��>E�q�Dvb:�s5���w�e�!!��*밣���0��-�
�e)����-��>���}d�|s�fQ��U�8�C1#D4�c&��?��C��B�ŷĬ�2\��Nm�2��ɿ�A`��� "$�RB��v�3���yC�ޒ"�m�;Ȃ�u��;`ŭ��%��6�xh�-�l��h"�3a��;�2�m����$� ��r'�>��kʼ���~�X�<�x�m�ޏQ�8����1ެ�i��m���lBKH��N�d��%	�B��xD>���UB�j,B��lf��n^�h�o�9k�ڝz ���]�0Lq��.�U��9M>�K�s()(�>V�YS%$�[s��4�'�Ze���I�tA2�f���Hѱ�%��t�s�q�1�K��sN�ż�s�*�i{Dؓhn
���W�O�Bn&|G^�L@c+q�6:\"�ߋ�_�zB-���.�����'�)���
z���!�{�4�HP�B	q�:�~%|n�����=+�y��wcR3O���k�6��Y���5��o�i����A��= DTp�t�o�M��!1�&z�mY	�0b<~��VQL���E'N�^�ݸ�5�ߙT��T{ޞy���q-�sbKj{BBo`�ȯ�t��@zCͬ�R�dѦ�qM�ܔ^^Tb���]ćWd�YK#�V}>�4�8֩�&[��:$�����K�d��[Pw���KR���l���w��P�f3�#�	Ҥ`�4�3�Qe�D)e�����������ll�^{l ��=2k$lp�(�BG��m��	ϊ��U�P��Ȳ�}f�[�qy�'�������T�<c��u�V��ѩ��*/��5JlL+'����T,��7b�s��zc%�폏��L^&u}ur�"�X��gw���3�G:�~鈉��˖����%���~kl�X�1Џ3���{����y@H�zo���) ���f�8�q8�J<�#M;���q�U,���^x���p2]n�������"Y��$���>���0���ְ|M��ı�N�������P1�v&s �5��������lr���t���#G�Q�u����@^q��%����i�_B8�b�m�R�0�>-�kQj�GK�1�,Z��]7���,��XAvD;�D��'ˎ}qnL���'����rGw�PICD����)��f����EaxWq��k44�rS��F��k9���LO�-@%׳�y�Q�>� �w9-+QF��a)9*�?"������c���mY�0�_?R�W6�Q��D���^��qd�4	�U�˧����eD�hYR��#��HU�J�m��&���r�������K����z �@w�j��*6$��yO��r<��S׼��? ��؉$t�]l8�b�d�� �@t$5�)�/��(��lhr`/�>�e�Jz�M���.ޢ�WK�K�l��G�bK�Pm�M����޲X�8�uYpd���&i�XMh�4Ed� 8#��� ���"\���G���U�X���ᦓS'!P�@��daY��ٮ�kr)R?����8�Hvs�������`�S�)��إb�0�|�y�}�w�n����՚��|h@h�CɒNF4���,3V2�x��J� �
��Wň�ǏU���i�ً�{��!��y����Wp@����w��C�N|c?�A݃�M��ʧ��"����)�2i,]��ԐeMc>��K��Z�Y���7�؆�C*��ֱg{��h�+l�@=�2���y^|�����T����B���Y�l�8��e�x��?�J����vA��V�B���?\��S���!ԛe� ��y�A |ne�L9##��9��a���L���3b\�Z�1�X����D���.���OGV/,r�C:�sӂɦ�R}��4N��4^7��{(�w�)�X�Vud�4Ӊck&�U� @}o��xF�L��W̆L��}ؘ�	9��d2�1����ˉ�2<��KR�Lw�Z({�嗚��H��pd��~1}kr�{�PP��JQ�#�CW5=�7IjO6>C������M�F�P4��i4O<v��@��Q�.�\�c���3�Ѩs�a'�c�	�#��\�(&�?��/m��qf&���nb��P�1K�yԩNʬcH�nش��MlIМ�bfC����X�Z3|�E�Ѽ�?8�XU�u�c{�>ġ��)��O8���ܯ�e1�<Q�VL)8k��nXhi�ੜ�|�x�Zپ!�a(M�\3�w�^��Ħ��z�X�P槭�C�T~c�J�g>���vU���/P��u�2+�WY�c]b0�5��n<�E��YC�u�@��e�H�w!$��ܩj�aV�E��:��C>�rM�}����!�I��awǊ*U���Ȼ0�[1$��j]B�%r1 x�H��4<�iű�Au��@��6�ËbRN��}j��3�����*�hv��\��.(R��8�(��_[�Ѯaғ��Q�r#���2�c�PC-T;@<DmB�9����J�cf��oh̭xxG�ޠ��b�cZ�uQ*�d|�����̵g�0��:�6�g�V�~�b<��u�P<D��v7�xt�q-d���.s������3-1��5��Sz�/��B�5�p��7f&��n��>�KK@����0�W�V�?��/h�k״���&�h=�N�����x+�X���1e�=/����.Y�$�Hv��������n�*?G�4����I�Q�s�|�?�=�n�O�"<�k�8f7
���J��&��^�+��a�5XBAO��[=��^��PO�q=ۿ �"*t����g�H�ƣXZ*�A�������80JUcy/�5��M�:����{�p%��u��5�1`�6</)W�z�Θv����CE�	�G4�2J�O�@�~�27H��]g��f w�����+P��~]��z�C���U�Odf��w��>@�t�̚� �uXU�$X��(���`3DVhD�T�J�s�a޻�..<��\[��S��׀&6?>'���F絈�^�Z*8u)���Щ��܊����M� @������\��Ir��>2MQ����J�{�~p���A��X��p%戫Rf�B$�76�!B�������L���afw�d+�8D2�㉡Z�:*˜jC�r�v� I
��u�l\ق��#�ݤ��F��|���F�>[P��>h��A���l;J3� �I�.�L���=�<����o�"�`U�Y�Bi�^�2p�&��:ˇ�
�\�Z<��'��Dzb��Pd^C�vz3�O�: g��΢�!�	'�
X%��#�A��aR�9>��k�
 ���S��6,���i|�M.5�I�/݀fuԨ� >��#$�Zs'j����;�G%k���E��C�p��_�]cO����ԩ8�};���k�^6��f�E���«%���z�����X��	�6d�6@����G�k�S�Qu��3SH��}��%��*�E�BA8��҉�,#���p"4C�g�q��☀6�ɬ��Ś^VVRg��	Ef�9$�rf�9Y�Z�=I�?������}��z���*[��.�X����߭�=K���O��+�O٧_04^IT@h��~��� �jj�t����4۫�K*)K�[����2`��JM(�$��d!:�eH���}Ԗ�:N��wK���#l?&d�N�G/��M��:�<�R�gs�3б�
A�	�O�Ǌ�ձr��w�N%�5��U]6�H�ڤa*:�O8�Jb�]{đ]�����Ā���s���:���FjDCª�o�~Ҷ�\���ܿ�-5	�	͆�ďO���|�nx�}D�K鯱ď�^�u:G�,��^Y�*�Y�q�V&����?���C,-�E*6x�	#	�]��@%1M0��TeK%���J�}�"�X)X�Q�	x+��S��#%�5�L�Π�s��@ڪP"���9��&䩫��7����ǖA䗷r涕����!��Nt�CD�NB;�~-̊�jh�G��]P���hխG�o�z#2���x�r�T�A�k¡x�1(R� �O��G/��:�7�^��
���h��M�j��{�c�`�_s�ܭ�8�p�([��������ь��t}@i�j���t��Uޣ,8���`ⵃ�R_�r4"و{B^囮�-;$ĸW��߇��a#77�P�5��8��U�-�lo��jX�N�5�i:����:)�39�ʼ!�����s�ڗ^v7��aAh�0_wN�%�g8\�Wo���d��/8��;n���x��V����:{YOOE�����|�(���m��dވ��GǏC�R|�i�[Ec�|Aw��"��Sށl���^�L"�@�����s����վ�P�r�y����I���ZNo7�k�t��g�g�h�������܆,w�@���R'�����xb*����q�/��6&@�/Q�2�q4V�n�o��2�̐(��(�<QUV.'8v���S���-�5-
�>�rJ���0~���W:����*�*�%���(��KX���6�-⡀�3�&��ޠ]�[�H"I	���Hj�j����Ƙz1��L��^��E0�i�kx���c����za�m���!=)�����a �^�tx�.�pn�#�>�����.8 �z��Mb���?�ݏ���,�6��50��U�<��eQ$Q*��Tϵ����a�}��)0�F�)����J���;�F�]A.��)�&���b1X�d���o�Eh�x�S0��$����_"H$�c�Z@뀄��A�%����h�nѣ�)_�8d���N�9ܸ�h1�j��qSP5��R9��Ơ^ˋk��(M�h�aڑ���3~�@w�89��<o�m�HF2eܖ��?Kt�K�������Y|�)N������ѹ��'�D'U�.)H���jd����n�Yq�c��G|�b�<	�A%�z�`h���:+�=h�������;4ה��Y(Q�XW|uW�h�/v���̃>~�� 7��#�B�U )� ��V�!��\���n��"�j��(Ӆ'r$��N_q��p?Z��,e��������� ���&�g�\Rⷘ������*e �G��0����I�����0�?�8dE�}	*�ys�C���A]
BYobR��*x4<@W�'�i�Lj�%ɦ*��,Q\��:�@�����=�.��$჆�El�B�q��j�?i0��|�j0�[�l�V9~��/��?ѡ\9��^=��2Kk�c�Rv`B�/ol����(�Q����2�!Kf߲�?��f�v�TJ>Gٚ�R�$9NJޚuRή�%�t� �gہ�-��������R!��a:��A�>��vT37q@����6蔄���5�ף�zG�`��[��,��,�)����H9��g}�{�e��%&V*3�hb�Q/�[u����xX��iҷ�%�'A�K,ԣAK}.|&6c6�9����s������#E�4ڟ��MU�I�.a^g�l��	�~&���=3����A���ٿ�h���,������$3n�J���n�?��nʬ�Jّ�+]��9��K 0R�����B$;��F�h�.�3�2)�\IQ��R�a���d_�R�Ȋ�K�����Ս+�Vz1K;�:��T�&���c ?��5+���C��װ�L�o�	>��-`�G��v�����F�8\'�=mC9t ����E�J�V��)=Z���0=Í�'���߲�����G���n檬WyJ���7Ah#�/J�K���'�H,�{TZ�8������)B̖:�N\��ئO������l���	IPЧ����YB�:�#��׈Jy վ�3ͽ��l���T���=�'���H��c�a-j�*+�?��y�z!@�?T�۝L�8H{�o`���J������c�B#���Q`���魹��B��?v8���C����;�b�X^M�Z�A��u�Ʒ�C��u����`C�Ƈ_�I���VTV3���#�Ȓ}*s��8�>�����x"��O����alI<�W����A���q��3�NR��D��g�Ļ��~q*�(|�ݬ��伅�HT����dі���(d��h��`;WGB�^���b��Q���1��ʗ�O���e����$��s�>I��Izc�g�T&�R;��/wK $���v���Go��X�&�B��VMT{�c�㘺�9�<#�'FEq��q�V��%�@r ?28�g%���xal�����Wb�^V߽���-�B(oR�_[C�)��^����hz_�l���n�&@�e�nu�r_��`��j���(v�pSl�C{�YS�:)kݚ��s��,���j�����Q��ri�tF	g� ��T;v��hZ
�[>)`pf������x/d5�3|Ċ�D�P���2��l8�z�����ᚴ%z��hݍ���b�L��Ӗ<?��Ű� �|7��`\� Ǜ��ݯ���9�m�;O���R	�_s����h'_ܦO��R����=��G$�9d���#ܡiG�0�5cO �qvy˝�C�n�{��^r��@ͩQw�Cc#<�@�aK�@>S�}�В"K�>��@^'Fn��*��_|���.T�P�?؍��)�B���s����\�ǎްr��&��ؿ�ӆ�Ғ��]~t\,±.65S�����>0�M���/�~"��g�����X��������n��(W4��]��`��U���\���$N�� �J:��2��&�:Lm�O
b��*�s�p4��>IY��@��^�vͪ\b�V�l.��9DJ��}�`��wQ9㬕mE_��P^$���ح���L�_=�3�r5Y>Y��N�j�
�yE�f�����O���?\ g��曱��w�vi��e�	�7Z�����E�)�>=Y����l����!�ʇ/�=�Lk/܂�vdW�u<.�,����eW�!�֏�S�S��O���'Ĩ��aP�$�N�����ߙd�=`��+U���6C`��Vq��o�� k�d8je��{��(%��X�>�8�B��3�V��c)Oq���I�6��{��lo�4@[r�Ň���;�p�1�ۑM��M�HĦ��mlg�Fn�b�P,\f�T�T�̭ʒ���gT��CBf�ϝ�����f��p���M��B\s��w�Z_����ݡ��e����sc��_|�ɹ
��;dx��k�]r�d �G���]�����iʫQ7��NewT�s(�3{�+Mn�*^"�X�mMk�W�@~j*l���"��ֿ�d�[v�y���]B�mo��6��[W�wYi�)����խn�ǀ���
B�k��c8&�RHT�g�z>�fbs�Q�3%g��� �Z�r*{��~型O/��oێ�gs���z�}� �٧7�� RV��A�ꁫ� ���1��K�������u�����v2����#lL��u X?x�m�"{�j��m.���lҎ�VV��Q�l�A~Im�����`�R��J��{��j�����#g�yV~M+}�D��c8��˙`��q�{�Fgw�T��_E�v�
�~�?��r��D=Q4����q��O?/�m'vTB����^|O��@b��O>��ی%�n7�Ѣ�g
,�݊��D����������m&s`}��J�xs�	ާD��U��굮v!|w��1t7JE�D��#�U-P���%d��ΆOv����^��ɣ~�i����vn�ga[3�R��4�:b����1ʪ�"�*q<i)��@�5?��2�@�C�y�����f�\�$�,��l)���dmя����WY|��I֙�!��d�PD�E�;����y�#&��U!���(/^�&�?2��5����%S��X�0�����P� ᮇ��)�o��Ӭ��oz����Q?����dTLG���tZ]��dͦF�Ǥ.�l>�t*���8���UWM����@�>�����8�i�,����%4G}x�]��aN@�B��ߏw�Y�k�-	Q�#���u�([�s��(N����\QƗ�>�i6�v�O��8�m�:���3v���z<D��ϣ������?�������Қ�wO9�:�~�zj�A�ޘx]��9o�n�t�����ٗd�"C��T���A|7�Z�'u�=~S����Ӭ�!]ŅL)����Rw>�	brT�ϧ����t��?�SB��c���lo���v��+�&��\��n���r*,��e�͖p"@g̾��w��cF�/2�~���l�� 3�9���&�Z� |nba��4��l�K���F������ow_?�	�8�M2����@ԕO���Ëe����`�U�ri.nl�V,D�#ŋ�ME��n�4Lgr@n&2�����@ާ'������Ӫ��#��;��Jt��ZO�	
 ���ڥ�'ҷ�Ɩ@�JR��i�fs���#�����tZЄo]�k�)�rE5�P	$Q�ͻ(��7q"u||#z�Yl������WR���.�.8���|�n���@�z`[��ʑ��ͱŃ��pT��	&��;�|�v�gNG5p�4�p�2Yޑ���-d���r ?���Ο��BFQ������}��wȊS�k<Mz�j1��v�*h)+t4r����ߞ^��p�� )���᧶`�81�+�t�;ô���!��KT��ܗ�d\�%��UgȔ�iW�s��?UAM���K�&��UD�qƽNf��My!�
�C�h¶�$�ʳ���㱝��^�c�?]'�$�j(mg�!k�k[?�UcK�x� E�N���v�����F
A}@7��P����]��R�B�PWL7�y��vY!#���fB���~��w����TT���
���ʹ7���m����ͣY�R���<�uk��_�Noz����Uu�A�{��ޒ�&�����Ĕ�:W��I>8.B2��ϼ���V�Ht����������ͦa^���4o��KN���_o��i�,�+x^��3>��~�.\>��̵ûr�&���"�����nby�g�v�e�u��W��Թ����(Ծ֒ک"�2�8_d"$�����6����_x�$̶^ef.����.�L�}�ja[��v}�7���	��MZ��m[��۝^l: �#\���t{9MGˉ�6Y8�Ξ輓&3��"Ưy��h48!�"Hf���⾀�f�n�o,٪0�A��NLZ�VY8`*7?#��^���NX��A(-w����-�*_�h'��8y��c�V�y�)�첱�C��D<�����L���:6C$��r��r�.����Y�u`�u^�򜎰+7@(rEc�ɿ� ��щ�B�DT%0Y��/ԝ�B�dt�!
��Ï	$*�,��v�=�{Uj|}��xn��������"�K;�ߥB��?��g�1���R�95;=�T���>J��$�}��n7��5
E�$7k�%2zR���R'2�8d�n��ɳ�2\����	F�#��qD��'�Q%���_�����J@��+/;DD+#���qF���ϔr�mA0�{-�o�ݦH���duoWi-�XZ�{�vI��80~MJ_T&��Q�:��!���|8o�������{um2P�3��P�ʪ��7��A9��ޜ��F�s�`��kݨ�S��Q>N�.����� �M�w���fv�\N�f5[���x�?�squ3g{>I�DXĀ��rc�>߄cf���c-M�?�_9=|[�(F3��������X��G*���k��Hx�zx�t�tꎊ�zre� ؋��w}g��'���PR�>��{�w�P�v��4��9 B]�5�t<������,���� z1`9�N5��*��3G�� �B�w��P,�C2a��4K&�?8N!O.�7�4�Nm���%%�:/�zW	���<q�!�p"�-̓��������a~ W�c��G,q�/��N2��������h���j�1���T"<��};�!�zV��⠪���?�^�	6�z�}I�3oNX�,\�� �ZÖ����<�!>�K�7:�m)_�)1:��t�Zpnc�j�J/���Pʌ�?8��S����{NdלQ�h��ZDe ���8�m���v-e��s)������0h#��0rΧ�}3BW��P���J��5^��/�b��X�=��k��Z��4� �$��o<O(t��ҽ���*�C���F��ym'49�.-l����}Pĥ��M�:�g�}z5M�����Py�9C������+��_IDڂ� ��t{��oh�(���1�ڙK�y���(�����
��^�$
>[煳}�u���V��V���ނ
����b�pG�H.�56�ӑ����bI���(�-cM���E�����(� �C�S\�����o�B3D��Q?l����R�ts׿}�օ�{���z�5��-/�>.K3VN�]�F{�`n��LSd"��V���E*o�G��S�4Bws����]}r��}�7��^��J�Q^!"�q�AnV��b�I�7/!�(��Q��8��ׅ���1�av���cj�:z��!/B"��B	-8��ֺ���8�z�!'��ݫ���"2Lu9`�湨��G�\����=��>Y�K(/��S�좹$�,�0AI�81�v���;�vT~6�w���g�!�t����`��!ݗ�E��oC%��3�S�K�ad|����.u����A �}��,���c�ڸ���}'���y�ܻ�Sډ�ES�gK1�=x���kg،��8�}�Aڞ�;��xޢX\P�R&ދ4�K']|%�[��{O�k�r�YRjDr��*��w��gq��;���	���j���c>��^L���<�~KCڸ��o�`P
t���щ�x�����˴[
!����]>]a�|�n;�����_@`��������@d��� ~�n��l�k���H���	׺���g����UDV���%k�YQ�?�p��Z�U=o!l�{�7��u��z[(];�|=$��H�pc�W�(ׄgpq�����!{�n�C�_��1��ȔPnD�صP�D�
���n��ȈZ�	�@<�W���@C�n�ܓF�{w�iɃ�SA���'����=ڋ]�[�}W\�	��c���=��\����U�i�O}���#}��qh�mj��G
v� ��9����F�n�^���h^�1�u�j�nam[�h�1YE��F�Gˆ��������S������3Ti8��\v�������N��}������.�n��{<�deЧ/��*�G�Y��
�����|]	�������PeC%�ę��y0���E	QS K�87;3}an�d}}��>���g�S�u�����h���4Ř	4X�e��,��x�>��������)��]w�X�6����}�b��c��h
o��E�Nܡ0�p`'"]����+ns�yG������.�K�5�`��r���x�Ke���<[w�\w���2'ݾ��7T7?�h��e���)��(�*X�O�a� #(��8(}}�c���o�����Û0d�e�|�a�����"]/��pM�s���W��e�(��Ʀ��Χ>dd⧓f�0+����Bei�R�G$B�ߞ�|��c'��U���UQ��T���e�Kl��ڡE��v�n>oJj��X:�pR�qb\bβ����'/��mߙ:�,�5�b
��S�wU�=h�q�� Y��?{=l�ߙK~�������i�e��"3G:��g��b��ծ�` �m��}��[B�?�Xa��Knߛ4Ƀ�Ű+D�#�{R@ih+�qNr?%|͖�@��:�b��sz7� ��Ɣ��4K=ȼ���U��������+�M�]�F�I�v�?��I�ӷ��޺�HQ���%�Q����ӉYHh"3t��~� (���0V=� [4&U+W�w���b���Ls#8;��iw0��u�J?0#�	��4 y�2�n�T�A������z"oY,{:,q��dW(��G��{}�U.�KD!
G��9��Ϧ�������s�ڰ�6_vix�[�gN�#A$�+�_��b������lf� vcy��4}}Erщ�^�l =��|g��C1{�Z���[�����m��O��b����H@"a
�z�LI8�k��x����6,|¥������.�]I�.����莽�dө��}�\=�[�ǃ�G%=�<谁�Q����X'L���C��4W.�̔7@�?��8*ü#���z�>>.�0%��}"�.3H8���f�w�Y��x";�pRIj0��U����.�@4��'�%��{CI5W^�_�-�������9��#�(�	��2��%�F$9�"씐u�@֋Q�mV��gv�R��:�$:F����R�~����y�Ӿ:������J��Q�?����Fsf�ӎ�$ɲ~p�,�?���C��� ��W���}�bh�BIf�+z��6��Gjc�����{'���!��3$� �*蛧�[�����0��(�L>�YY!\eh��	��0�h�cH����e�`V��{��q��֬�,|~�{hd����ZZ��M�-��hy�.IJ���E
EA)�kύC>r�%d���V8��@����I�u2]�e�6G�ZZ3�vM:����L��'Y�ĥ�]Sa��B�Yhq�ʇc;�t��9��?�a��ahH�V�RȗU@8�buM>�j��F���>�*� zZӦ��D�u��X�DF��B��;���<�Wh��K����}�MWv@d$U�(��Jj��y7��.��m3�<M{��g�'>M�iEq���������>���r�Y���ƿ�!�8�@;��!�ն���+Ķ�h���C�W��J���Ix�~��,}9S$��4Q )k��ю��b���F
W��p��֪�|�v��|^GG�ܥ|�B�Qm� U���W�h�.2���t�W�A<	�!�E"�_�HPF���I�@�FKn�$)q�����k���^�$�Ōe��N@������� ;�Y���Yn�U�Yf��I��F�r�x���K��#P��Ʒ�uw{�V5�f5�`;�L���M�Zf&e��Sͱx���вdY5��0���e��wT�`�V����t8%����a����ʸw:F�<�|��lYk���gC�
�/�z����e��Lx�@^�BQb��q�Il$�8�wd1O�#�〼?��Nfb�t��q��C!X��m��غ͏��g�@M�;��UzӲ\���T��qP�Q�w5�>��o�9���Q'D�V�|����'VUL�!�}����l�A!���\��>�@з_��N���'ZN5-n�,��L�Y���� ���74�lU݃��	u|v�3E��4��o�~��;1��7��b��YA���֊$��|�F���=nk�>����?��{d?�RWw�>������MrA��<�&����L��;u��f�Iۥ`���L�A��AdU���,$��t���;Yꩊ�/s�zf�G�� �n�zn��"S���I���V����j�u�X�WcGDp8�>O�+4`Ϭp�/��=��t�&�({m�"EgH���r����O�gƱ@EN0�P���Mj�53E�$tE[� g
t-���
pb����tA
���<��]..���l�g��g���޶�n=J�t�����B}2i�9IB-P�aK��y%�vY����ͻ���h[��0�v=�D� d#�r�����{)��$��ʍ/��q�e�]�<`�b�غA���e�������>�k��M�����@^�b܀�Y1�[%r��o-J�vO9��u8|"tq������f#�T�ro��c�m�,_j�ϭL�؞qk
��=V���F���3�w���O�2��_Ǯ��h|��DϪR�
����2�����"g���V6�l�tY�9�vs�6
����~�<���#���=����❭r��_���_�0�����)�����ώr����
�c8E�� Z����W�L6������tj*�1�,윩��4�Pb��:�>$��1�0��(��Kg���Xo���f�G�� $�Q�PB�m�������*���u�%�xDWf^�q�:8�k1��mE?�.e�!�c����~p��Yh�|A������iU9I��)p����e�"mj ]*n_~2�h��1�0���҇���'8H�D�_!�Bu~�p#ǙX�����Y�I.|9�E�/��ha�Z�xe�yp�X�C���p�Q`=����/ԙ߂��A勢H����U��8���S;�@{&��\�����H��(�q��]zg���	B��mP���4n�8���.:(v���y1
F�<'^��{Tۻq[x��'�*�k�� |HhPGu�,BD�P�Ĉ�
�%)�h>�	����!	T��7�������X�]���:�d��x�^�N��R	3��O�{���ꫜ��j -&����/�Q