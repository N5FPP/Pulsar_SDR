��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>%��}w�K���ē��fu�}vi��U�㶘�ㄍb���XT�$���sݜ1�=�5ޓż �+ןp����,��K�D�׺[��3�m�9N~�H�&\��D��>�԰vf���֘N��s����7�{�Wy0��}er�)Ƅ���4���I�d��<�MM���l�:-\XgdJ�n��XJ��������@����!���O�����e��}��~�?rt���v}w}F����Y�����ʎX���Wx�m��;�f��<��оª���k����sYX�f�g*���K��������*�@�/����:�J�p�m"��9��#S'ʛ_�#�y�ϵt/����K�!8J������Xa��m�Eg��t]p$� ��L����C2�|W;��.e��5�ШB`��U��dd��0W~eݍ�#Y�TX͉�R~zhb� ��`9h�0к�$��h8�r�_�'��x��NFR��P?O&����4'
��q{���8����B���[����(��M�<�r�h�D68N6�ءh��&��jnB�Ld�0�fx�,�:��ɮ���Ş�]���ĉ�V.KɰE#�(��z$h�}��)<9���u�)jV*�d�	�lf�6c�.iP�KM�~��!����.�ڣ<1��%إ�Sf����h�[{"XP,�����l�#������БY�f�ٞe��
o�[
@�U�Q>ï�8=>Ξ\�kfp��tӟi�݊X�a��8%�}p~������9~�6x���D�G�x�� FkPP�7��cL��i']�38�Nk��-�X|L~��9��@.��r��x2B:��oJH�X>��<D�.��#C��S�񎴢�/�z��n�g\��ʙ���S�_�/�?� ��K�@/��sxs<%�B��3�qI�������9w+!⧞Y���R�wWG�]Ϗ�j��&I��Bf�D���T��Nr�M2�*�Q���^�D��j�k~l�n�)�N��_ȗK@�%�K��b�W"�3s�}v�,��1��#3.��jԠ�B5�0&�ޅ�T�@�թ�4��0&�!֖����q^�<#�+_���N���(6.��$�����ց ��mA�n)��Q_u;P>8�T{Ļf��i��ë��J�Q�3x���n`�phg��^� �����뺴`��T�*��ڃ�J��,l�|A����*gl��R9E͠�>�b���[�	վL� 2G-~��3K ����O#��.:I��	ηM���Z��'�ֶx9w�I�e��9�=?����CR���*"���,�d�흉S�%�8m�K��E�H3ܢ'�t�����P��d�X3o2��v?��&m�@�c��]PF*MQާF�����*����r5$����4���
ۉVCčb̗��Oၪ��@��X�ם5���aׄ��>���h��Mz��x:<��d&>n{E�޹HI���}�z��m%�|+1o��դ�fc�MUu��B�l��@	X�5�� F>`L�zkX ������'��`��Z-�u+ll��r}c����:��~��֫'x�GK�>��\�i�� ������X��\x��o��HI�����B������9�dp�#�r�M���	v�W/��0_I�����G5�pE�R����H���=^:�;D~��uH����6��5b���L�q�/2 �C�>�$6$�Ҹ�����R?J�S#$.��a�G�:��<5��,��_6l&�1~�\'8� ܌V�­0e^0+�� u�g&��c���ѷ窋j�ϩNH��|4<K����Le�딷c��|_;� ㏹|k��R+7�1��N��I)~�y��	:s�71��	�����xd��ۖv�ww)��o�׻KK&b���к=3s��L��
���j0v��^����ίY�559�U�]8�v��DJ�&�����,o�1���ȹg���skca߇M16�smq���"�h��2���n�����+�����]i;���!��hM�f�&u�z`�T��1���>�!�ڐ%2���Aõ����g:���"1�E�s�c�\6�`l�D�q	�wK8�X� ��/cS�!~��M΢���o�s����v	�?41�x#�>�e�����걥��g@/���d�J�fK'�B�w��6� 0j�c�Lǃ��5�D�9�IT�R\�	G������c�Tڠi�o"�.���W?vJTL	&%4ϼ���t�����w�)�%�K2"�VK�H�U!�Ϝ��,����sY���-^Q�����+�F�d'^������UY2�����@���x��ð��O>R��Y�h�;E�q݆M,EU�R���8T�G���P6�����>��Z5��6N���F����BG�K}kz���wk��2����8���9�PI��V_�.���Ei>�q�l�$��|��fW���쪬7�B#�}���P>���Sc_��z�[�̜�5/w�B
�	��6�����Q/<?���+CS_����u?���A�=t|Q+�[eu�%<XC �%l�2[���'��oF���He���?�a�����l�D�C�>|�Y6=(�z���A�N���Ls���Ow���c��>���[ {O26� I-t�S�ZN������G"�jڏ8�($\֘"��j�����}RB��mt+��SN���:].B�Ñ�#�Z^�v����9W/]pC"�i=�1\��-�����(P�5"�ж������Ĺ���E�Ζ}{k)Q6��  �+t��Ł&0��v��6��BԱJOX1�&=�����Y8�Ϟ���(��-��o�o�wX��@`�bx��f��+�J�3�w�'ޛ<�O|�;�l�~��Ⱦ=���J�	�	e指U�'m�F���:��IѰ,m	XˤF*D�r���DN�������.��	H�4�����;�{^(	�1��g��Nc����e�-��9]3�kVh����׵�
7v��ɗ�b4=�����/������#o���_WF�i�x��� � B�����'_�8�-X���Q�?���Af�M�.�b~��Н�e�~�������w�F�gO}��y��Q��ʒ���Ʈ�Ma�����٢Z ��gV[��1�����Uhs��󟴮5/@Glx�-N@,����` ��	�����V>(c%$R�d�W�������_���:�C"��'r*&�� ���\�	��ַX$��6w_�]׺�b�ǻ"���t�k}^�B; ���_k)+�u8O�ŏC�Jeb�t��}�s��^X�_'���̹k�n!�q�����o}�9<��
t��L(��<�W8�����]�f69+&��2=I���{�2�3�_r�kY�A���)xT����SBRJ��hb�`����i�o�O0�ߠ|$�QZ,�^������ �ŗ^I\��g�3�z[Ƒ�w�Vv`�G��Ġ	�gB��X��QdG`غ�n9�\����R�^�dS�K��2iz�V|6퇛�&Lg�h�3�۸�n����˺&6r�AL[OZ��!�ܰJn�^��j{��*�ŀ�(����Q�%�եaɳ�x�z<?�d�#p�&I��c#���Y[T�$��6g�e�W�����B����M���/6�YxC:���Z�\�H�n�v�=惞>K,f�	��։>�B�j}�1;HǞ�N��NdW�,�U�)����[���"���(W�x>���e_�ImWP������&C�&�����I�-s��� 픷��<��ۋ�0��/�� '
�V=9���(Y��]Lt�I2�9�F�!f�U��*x`f����.�{��7�)���ZOk�4m30���"��͆�6˦��:�oW�e�edZ����y<U�=+����Ίd��Shw���E"w�Hl�N�'w�:��?h��e���(�K�.���Bs��'����9Z��1�̯��<Frm^�N~�֟����.�=~�r��	�#����=S��:!"�qd�q��8W"�	�k�2Cv��O�v�����`�l`?�������y�Mܼ̯w�B�%�����]�������۱R���b@R���)�3��;m|��gC��ve�J�k�^F�������Qd���E>�`8�����u��`�@HR�/��j�ЧOM�	z54ŤT�j�����s����%�є���tM�����L�������b���yf�pJ��e3A����u7B3�t���8#�Y����>o���]�Ұ���0?&��{�B�6�
Юw��D�G[R&���l�X���Ro?4E�KC��D�G�a+5����	2I)�2f�M��A|�oӽ� �u�Z��Y�'���+��S�o��
�91�e(�9�S`f��OV�[ �k8��V����7��x9�|ob�2�4���j}�1��t��j._E�������P�Z��y�����f�CL�Xh�"I�
�)�55\����&�&��w�lx�g6k�����dX���\ȥX�lV]0�vU��\O�u~D$\���9g�'�F���в�+C[as�b'A�%�$�[�r���6a�A�ƑS�y��5/�t}4�]�T���t������܉p"M�-�X@I�'ۋ,�.kd�}��.%��f�m�w9�;����䷋uV���Ƃ6�-���{B;���^�9N��6��hO�rle���p�hׅ�rT˺�V�B6�z�zϡ�#���1�@�\�
����J[l�:<?{]�����ں�^�/�XC9m�-�zѺ#�`|���^H����oڪG�6'b���۲bA�$yO����
��?�zC!���s~CqP"cO:�5s^;�@������C=�Ln��؟��m�.b�y�����p�,D�i��_Bxy�s8D�$���/G��n��n-vI~R�a��T�ɚܥy�����p�;}��T�̰���:�e�aw����Hе� W�o�����㿽m���ˁH��:W-���tGxC���*A-�';,4Y��!���3S�h}��f�;"m����(����b$4�7D2wl�Omp߭ =m�.�;)K�C��Λ����)�$a	�h��OXt�<Z�h���3`�X���K$�%��捷i��#F�MY�k�Bz~��/:��}��MÇ@hva+��ʽ�_���|z�ă� +��IA��- �B ,���)�bqɡO>���,*p��}G�2ŌA���q.�=�uՌJ8d���	�i�º"|E�3� �Y
w %Fla_F������ط���_��0����:fd�oZ�|�J�x�JPN��ˏ�TvG�f���M�Ї�Oߩ��9Կ��12��������+#X����uw
�����Ùb��D��O�a<wK*�����֝�4w@G{�[����8���Ov�+�Ll�nw�s�T�f��k�PW���pd56v���$�l��r�ۏ)�&�i[}/.\Ã��q+����N�#H�a�� g(÷k�H4�TJ�A��zjJ*%����Fh��V�C���֔�Z�4��|��]�6.�����<`^}KeQ#u&+�>z����.��D������`��/B-�ʊ/8W��5�¡3�$��b�����"h��hA�b�Z���x_��I��QB��i�rk��]
����/��@�5!�p�p<�`�G]20`�HA��nk��`9���
�r�B�߻5rߟ�QW+����U�5T*�1��>	�M��n+s�2��d-wpɫu�R��(6�w�V��\*�<�C0�A�F�z1���-vCiUfk*���N;F���s���q���I2�ɹ��E���$�P���k^���u��h�l����v��w|����ۤ�j���=�\�WTFɽ��>[v�o��/��񑢒*�N��n��d�_Z�rH�Z���A�;�ґ�͎U1?â�7s��:V�h��⳴J.�{��{Q<�k�J:���AZ�(�S�O�q]gԃ�Q ��O�{���G��VH+���+e��XӯL�R��LV._��P^	%Ă��"�*W���u�	߆[8��0�Wq���b�����cMf�y��J	��x>�qp2����)HЎX���0D�Tᡪ��-�Pj��n'Q;�?c�3�e	�3^*�xa�665>_]2�-���#Vxd ����c�WLP�-�2x�R$�Y�_�2'���E��Wy���`�zQI�Sa���U�v7_t��Q&1f�>��頷�i��B@���K��î>��E�d���C��������Θ�i�ս'��+/�x�C݂T�A���S�/e��`� jT
�-�C����5�#9��(z�=�-��[��z_����G%b��Q��#�2m�w�cɜֶ�˰����RZu�Fh�0�H����W�vv�܂��odXOj��@F���h*\4�r>����rs�q}V���"�������NW^�ƱI�wg�;Kl�a��{�������Z�2C���e��ſ�S��P�*�Vۖ�lq�|�W4��,��1��K^�w��m���^ ꜽ���rӰp��^N���_8s�	�Hl��9!w�
fXkAz;349��~	X#�͞rl�Ɩ��7Zm;g���J�a�n�¢nչ�"{.&S�D.������4f.��=
������>�ϴ���Z?�MH �xjhk�j���#LE.ޑ����1����S0T��fx�)"���Ag�����]�mm�6����={�Nh��o9����W�K]�mi������!_S�m��}�waBHŐ<��=��c'�߼w G���'�>Үc Ѷ� �%�j�J԰���-����*ۅ�	.*J=�����r@Ӿd�RW��e�Xy���O�h�]����L�u��jO7�$<*��AMF�\x���q�і�hܿ�wr'E{�a�e����e�2P�u"ǢQ!kcɔ��v��垅���]w�h�v��]R��I#��^�Yč�t��,�s��4�<���C����F�I�s/��4�Hc@8ѕ���	�|���}�3�U�xe�kW�S�;��|�tZ��r<RFZK��t�M\����LZ�ZN�A(��S���2j5�"�X�h��3�-H�)��������&FH��_`-�b{�I!Y�Ҍ4m4�\/�Ӷ�E{^��/2�
g����a}:A���M�����&E����TN<ʸD��[9G�����nݫ����H�X �w��;��w__�$Z2Ы���������-H�e��xWS��B-8�8��y[7��L��~�q$}��V��w9ށ}�i�n91�b��{��j-5  �6L��x�Ss�L1���/7d���E��/�7��?6QuP���t�Ί�B�c�}xYĄ8;&�4#m$H�=/(ʮ#��4d�g�����E����<��2���˳�x=H�0��Ŭ��R%!J���ߜ�r��9�/X��*dlʒ�Uvc�l��9H�Va���Z���-�9Ӂ4<��PhTG��|��N�|����m|M���.mhծ��o�nZ��4�A�W�6��4 \J{pIҟC���85J�E��3���h�����E�t�9FZM��Q=�q�S�����o����ܥ�}�*}�u.�l���#�<{JH�;?u���������*�R{Pl�=��A����L>եJ�tF�{�B-��t�+jO���O�FD�^e #�_�W�#L�9r�ޟ���������1K�Lh�.��U���[R�t~�n��Z)�} �FƧ
'@���
 �f�P�@��(�)ۍF�ib��;$����"�J�;��݁���unϥ3�TPӖ&~�Vv�S�ix�::�I��r�(qxg�;��{����n`_6��If$\e�7QnV�-<��U�W4�{���;57F�;��R3�>h'ή�B�]��)mo���1j�=<�Dڄ��٧��:3L��g>��j���h��"�Q�8=�o�W�)C����:�ShbC��daý��'���p�r@`w���u9X$��+�,�V�X�D�xo�A]�9����x��N����cm�Iؗ�1�w�R�0d��]�1�/ l���:�c��nJ�@oiYE�Av�F�}P����F��&��@��jx�3r�*�������pq�6�[���Db��M~e�����:�S"g/o9�T:%6
�uk9-q���0(�a���
7S�B�Y3��_�?��i��f��L�{ܰ�"Q;9�īl4>L�t�e <��+t�k�9#�����J��RKU�û�T͌T|��l97zn!�5�ڐ��_?��-�F;܎�~d'i����P ����7�ʏ�7�$l�b$R��4-��Bcq�"��km�7!\� #��t���F�o:L�����C�ߴ��e�Z6��{bs�3��S���t��������6�r�y쎲+)2s��j��k��w��ӐRd[����J@z�w�U*q֭Fl�A�M��e35:�B��]�P��3���Pt��ە2O"؏��Nv��x��&������2��՚w�t�4��Q���J��.�G��k����� ����q/J0�~:PC7�Y����ds1�SL��&�Q}�9Q)+����}T)�v�Z7z��y�GMv~ �a������
��
/ �T�k�I%t�˿�s�t
��G!��o������|~�Q��]�R�������x��2�|�n*���B�E�7p.�����H_�'�⪉ܹ� ���Up!>)!D�E^�,)5���i����n��6�,ߡ����������f�}H���b�8R���@��H�{֏d{�M?�P�wj�~��a�}彪q�>�9��eG$?~��x�4�����˖�\g���r�Ϸ=�mDȁ�l��@�/���"���ޣc�����5>~zG�o��������[���V/����Df������]��h�%|=�uU7/^I�=�!�J�����75'�Z�z�<|�b[�^���F��������*26���(Ю�O��7x�����A��!ؽ�]� U���X %�q��LV�sIk���_Fꊽ���Ԭw��0�r�#�۟�<v��[��ŞD��Z|J��焆�PEKA�qaDp)�؀@��᪣��3+7��]e=n�Gq�1|�2�c-��Uze��!.�r��?�z���U�+��>�j�}��	z�&�(i�q4ߞ�Ql�v \5\9��7������[�3��w��Bry��៚t&Ȫ��׭S�*�F��ĕ�o���.xgu�e���v�ˏ�H���D��S��l2*�Mܛy>�����!�	1��|�D�EeY�߸G)����U$�nb����8զ�咛��#s$��K�,��y)o���<�|1�2!�7��sJ 2r�Q���r& �r=f�����lz�Ɨ���B3��a�C�ћR�9K.�)QO��ڒ �De��M�&qo]�wFS A�8�IZ6�{5^Ԓ�Wk���P�.ΡP�mM���<QR��S�vo����}��\2�K�3�u�?vQAX��� ޾%=̔D�a��ə��w@�h�q�#զ�q����lu�3ʖS��y����vՎA�Hx�6��t dz<���)���7������*.���Dy�8���S�ŉ�����]���{��V-�2^;]��8Cy7D'RtUP	>�?ib�zYA�?�>$+gj��B��lk� ��� J�i��<���ːi},O<1�|s�w��M�x�������>�X�=�*\w�hk/����	�t}�/k$����Z��tP��Id�Z|}�>���ADwz��OT��wskCL1��/�'q���k�	%�5ɴ9'��:�-PW5��;�����Yǵ��D)�ږ~��Ϟ��@k)�45ɖIL�l;\"�ӴO���P\$��t�Ϗ���s�9;(Q�
��F��������Ä����˟�<Dg������r�J��%�
ҽ��e�|\���'l��B��6`%����"��	M�Kjn(V��N *���k'O=�Jł�a��X���%��9S�r�V(�#��V@�w�pF'U����-m��-��r�$�L�����x�޽����O�F�;Q�.�J+�s&�8c2��$��`x�[���"����<~��2�bS�?�roKùsS��}�1����]��bͯHD�#W�*c8�C��J���~ M�	��]�rr~��)���U����Fe�{�:�8ǹv�i��h��q��h#�e�!�9O[J{�,��p���uR�	�S����<S�b���J�L��m~�����q��tM���N���y�c+Jm\H|E�����L����E;Z ���^�s �>�b�߽�L�jx�Ky�P�B�(d�qc��a�[q��A2��u�,�4G���J���3���gY�ͻ~�%n^\���e �89�a�ii��yƯ��$VX���D��l��U�3j�9�^n����I0�{��@,^��r��� $F���gŖi��=���+��a}or;���Ƀa�C�9�2}�]��:��(��JU*f�*|��Ӂf!��h�Y���4�����	{O��WPxo�Ӝg�J~2�󡛙y܈������M�|K�4���K	�tb��I��~�t$�g��>O����{@y���(�C�KGҰ���g��SKa��Rf��l|��)P�+ܼ:b�C�a+9[*������oɢ%0���L���(�������%3b׎��Ai���&%��,Ɇ�URLHfZ_=ևHm��Uq�l��u�
]ݕ'��Oz��yM�yl�[qJ$���
�.�}�qj�����%+HR�ТU��$d+�z�sC[�s������E��H$͟�/5"�;}z��X���!"0�R�G��K&%θB)������9F��P���w�A��Q� �^o��14�Y8����t���Ӌ�M�)�n���V=S�G���"��(�M�u"f�:I���n_����p�b�	�xC�lɞ�����ąW�������)(0�FR�<Q�%�^����M2�t�$��ˆ�t�}��#�	,�� ���?�O�t+��ϟ"�R�>�iK)t����8�
?5E����/�U� �1<�D�m�+��W?�MGy���@�B��"c\b��[�T�؟LR�5J�ʠ���l�ƨD���z1'4�pN/؛���6a�G��֐j'���pH�x��&�w�L�K�Y�:��v���!X���]��ĥ��˔E�Mc�|9�2Y����#�"�3��n���J:�ס��.Ï��gH^�~F�C�C�CqN�*�"2�W͗�W��B