��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8SjfSު�U��c<�`|�g�J�@r��c��W���J2iO���7���d��t�#����3 �SF��%u�l�×ElM��{i��O �cZ c�R�����+Qn�޻�yv}T�m�O�D ���@.u� �[���@�+%9�Yف���y����&_����$�#sɌ��Vqp��<�/��X܏ᢒ��/����]��e�Gc_09��v2���;��Ĥ#q!� $̑��r��@��-�J������ꫮ@s�t���b�gi\�{�%�;���Ɋ��8�W��V�>�lj��/���5�E\�gl�Ħ���S��v��V�pr7+��H����8ȶw���m�u̗�_t�h�%���xh�
�t����<��
��ܶ�GY;ۥw)?��tO���d.���k�#U:��~B"����2��Ef����7Q��YZߝ�����k��euh�"��}y�'���ܑ݇7���{��&��B��8���V}@͒B:TZɖ�Tb�Z�D�$� j���D���\Jй�%��?�`V.�0G_ N�PPͭH�εb)��}c	�{��i�(���;;������85,@�i�|��~ڏ{Jo�$�u-�D;�X���i����_�6�OK�Oߒ���˦F���if@T���`�=� ܠ�4�U�lZ<�ZA��`
�R��N�̗E߆#|���D����EE�Q���76���ao���ލ�<��.50O""C��ѝ���)D���d�X�5���m������D,��pJC�`������)��1D����NRv\O :@�m�!�tz�0�/����ţ)CճG��y�}�����.�]�l�'�^��BP���d~%���#�E�!.��"́��($<��U(�є�,�A����H��;��ߕl��7� ~�����(�E�ٟ������ӑA��p&`�e��!�E-R�*U{���H^!�rYo_��x�"�ٌھ�o�6��ԩT�V��b'�S�o������G��ۿ��� <O�j�#?�.��mI�v-(��T6�d"+�b��I�1�҃`�{�g��n�(C���Ҕ���$h�|��9�ں�dI�")#2���v/���[&�`t)�Ր�$a
Ӥ��E�����Ъ�����اS���vل�$������Ը�V���7:��[�ʅ_�F@8�~b5����3����')�L��GJ��Aڙ��>���%�A,��Z�@G�U�ǹ6S�u���V��ǝ��=I�8�Q��� \=u��I�X�[�yC��'�1� �y��b�lxx|c��d�l��]������]�Z����5�m�L��E��d>�@n�5/u�����杲/W�6����ׁy�)7bC��פu���$�.��V<4P|q��+���x'�|[�N����qD$�X���0�2P��F]� n�IG��P/67l� A�P����Յ�v>�ҋk�Oջw:W�kj:U6��v׷�"fA�Ez�5���8ᔏ 4�s�w����5� l�U}������D�h��z74�3�(��'��'�oOcKj��W(*��\0^��z�ɜ
�>�yY,?�����2��a�R|�P?�}��`��{�b�������f�� �2e�N���~ߜO^�u��Ӧe�'I��.�Wvz��=m�L�3�-�������M6����~�7i���a��`vm"�RxC��.�#0��Iۑ~��7�m=�V��a�b^����F�,��L -�����ǁ�b<�H��Ż���y�\��X�	#����
�W��m��'���}�Q�^E~d���e��7D��P�hr�����3.�I�� r߄i���12+��Sǧ$���J��]<Yu#ݔ��v E<.ʴ��V�Ʀ�6]DS��,�6|���+7�J��]l�2���4b��-;W7Y?ֱg��9�Ne.ho�(�v@����m��&��(+nҁ�F���|W����W�xȬH��-�0cH4�A7����n�SS���~�|ݱ �m��~��K���}�7K�U^���
4e������f(�x��P �=�8����za�����1�J�?�����K;�X��xܲg�F/U@Y�4��}���GF�++�@���9�:Ơ�o�J��@|����kqY�OQrwj���=:��ǽwC4��7�
PlBo�{ �E?�����{�y�D^4a	4���!���e�8�1�"��^����(�]l%
�w��pa�<j,Ed̄�]Ǻ&.��Mq����aƚȵ}�3��O�QC���5�<"O�_ACtT�"H1�i�=&���y���e�to|�9	�ъ^^�-U�_͙\��qe�mr_zK�$��K��Y�m�%R�g,{CK�3R�[=!w>�4?;�U4�&}mm4{؈u�7`�+�*�Y} B1�o�P`�\�z����3%Q�?�'�s\	�����TfX�z>�i%T	;*o|�Mn���F�K-~���3�Dx�NU!����4��S֔= �j��i�*95wy:Դq|�vq��!����� �3�^;<�)��p+U��@}��4�i&Yz�9�%-�Xq����ğ��Ο�s��D��["Ɗ*@�ۘ2�
��Z�l7{C};��$�Q��]�&B�Y�f�!���x�i�WG�E}�(�7E����1p��d�*fd.��`����������
|�mG*ق��b�O9�8܃j%�M�+�3�;\@��ԡs�Hb���v��C0\��?aз`Z��H�✜\?ƨ�i1V�T�?b<UU����ĉ�=Y&���'���z6���Z�)���%�6ןU  �o�U(��V���&,g<��R�b���Z��F�,3�X�����;[�e� �e������t'�0Qaa��ޡ�����{5zC��C�K�K�`9\`;u�P2�<�Fl
'Ͻ4_�/�o:y�V���%�j�m�v�1��� �M$�J��	������%+m�����F���b8�=J�=�x��7,�Q|��s�
I�釷G�v�(wT&�9�l
��^%ުPi�q_��P�2���i%�D�1�p��2l5*�����,b����匂ʣVz��zj{37{5mΪ8L�/�>�:}9��p�4�w�cX�;	��3��)��)�����7��T
���!޽ F&��L<jLT�s�\č�D�������Ϸ�'���u�a0�q�;=>^H,���sf��u�fV�����N���ao�0�W�mr��	�t����>��W�
_��[.?�	�K��es$��J^�CĬ�����6��1�������~��k�(6���8�m��֡ʸ�Q�g^���L$�'Oـs"s��|Ql�Q��7ܑe�u�U��1ϴRO,�&�n��=#/�6�[n��<4�`e�m���~M��ZVUu1���������W�0�J�\
tu�N8T�9���lF���n�ac��c�K��Qk1�8�=� �q?�tG��zˌ�\������n��﮳qN;KN(9\[F-m>G@�����K�'D, ����r��2�&�1�`a�3�4k_�Z�!ܝ�6��@u^7�9��?�0I�5�}�jV�I��s�V��Κ���4"Z�m<�M+Q��\+���$N^L�dw�����V�M��L��ɾrg:�f��z<�j����Q|���U9��O���R+�$ȷ�aۛ��SP�rK��]
�A�f�{���4(2`{��[R������c`+w�t�8[_���P���Ac�a��04��8��4�Rz߂����FY#��!>G>>z�f�b1���P�H0s��1�d�b��d��"����C�cPH�
3���Z7��+ $�T�)��%�;$���d��C ��+�$A�OO3T����r�MgE���b�1�^Ad1��AA�3�d��T)�3
��P�Q�>Z�I�xv��}��J�,w�5��;�z}0?��=��8`*�F�z'���rU�I�se�m}�d:�D��M5p7LJK�	���e�9�ZRW�iw������SS���$I�n�3]��ܤ*/ӑ$�&]��G�;3ZK�?Bz���3�����v]���]�AϨF�ڠ��̏�ȗ1������ܨrAl	`[�'��wo�q<�[8>���Q����&�`�&L�s����i����S�/M�Ҹn]C�"S <v���l�#3�`��U�y/���]�g\v���[PIX��ɃR�X�L�h=O����(,�@གp����eId�^�R�����+��a׫�7i��Iv�SQ96�>�������8Q�%]���x�.�w�I0S��Fn�v'��R�"xDMp�����8w�z}眤�bu�'b���\�/���{�<"J�!����<� �0���{��/�ӏ��I/��D�/��_�/�H�u�llq�
B����=����E��KP~�2��z0���EV�1��!�7�㍒��p!V�-'A�Zʈ���7A}�1���o��Ґ{�h�-��~�$NO8��Ә����Í�_��[s�F�8���#���C `��SV��}0��?��ŭ(�/3J[zR[��� ������/�.ژP����:�@Jz�J�3V1�Ґ�*A�=\<A@F� 5�c)yC��J�l�$�b9�S	�/�U�SXW�OӃ�K�F��� ��y�A��
��n�q�`�5�pi�_����E��sЃ�Kn>�#��M/K�ZzԆ�ߙN�)A�LC_�ܦ��򀺋�KEM\�;�����{r��D��K�g�kӁg��&�����R�����5�����2���A��Nԕb�X���.�e8��mD�V=��O��p JGz�UF�	��b����axg�k�tF����C���]y��z���(;y=���2H`�:*x�xо�Zg1dZ��M�F$2lNǌ�6��	ۭ-�"�����-,��v�Fܕ#s6���ـ��%���*zY��a1�Gh#���v����1mr޳!�F�:�ZC�,z� J��^��,2l����v=���7kPn���	�_Y]������oQБcx��}�q�i���I)�ጄ3'Em��[�Z��(��iD��Q��Պ�V۷I��biD(�r'cl���Bm�'�^[�c�R5���A���heɨv��J]pW����y�visv��u�W=/���c�M� �=O��fvc�`�~���v튷�Ҁ�<�c��ȀgM���0��^Rqߚ���R���,i#����h����(Z
ш6��;{�؄N]&=�~(�"O��L>d��A=�8��?W�a6XÚs�
j����}f��C��\�j���\�ǋ�!W��@bo��ahČ�E�%sO��U�@�QJ�.��Ӛ���_S�ֵԜ�N]'��|rN��7W/���Ny���*�W��6���ߘ�w���rV݊(|�q �=>od
?�f���b�~S�@?��FG=�ٷѶ������4{�UW r8��0�����
cƥێo�xZc�e�N���S��ta��=�w	���QPG�a(\�9	 Xx�j�nU�<;�L��bN˵"׻Z�cFca�A:Ea"��\�QpO��0j*K.�za���@:5�2�/6ڰ%���M�&�2�lN��k�N*7wRK���³z�U"ds6�@�@��������5�12Qэ��`�jο0�U�-�
*��4H�n=��ՋTV^Ox�qs#�ܲ%_n�R�4����J}"����h{�٬�k�a~KE��_�刉�����cij��ˍ��)
��]Q�U±��T�P]�O�����J'��PpdҔR�G9Z
0�Yㄋl�5�I���z<7ݱJi���p��`xA[�>�0'��}��4/a���� ����~Ĺz���16�e8!�����4��VI@���$�nq`r���}M"���?7��8؞��q��;���a�Ü��C��3��@�4��L ��m��3�YQ`SGh⇘�P/�-F�KC/=b��ןj���^�t�i	�3m�����_�U��Erf����0@jspr����5?�3��6�yp�F˵CK�
 b���{/y@�Nc�W�����ˌU���E�[���D]�<�l�C�T@l�G�����l\S����Y}���`?�,��S�#��bc1�ws�8f)\bx/*�פ-���E�O�trsx4 J���={���a������[.|䓌�4�p��
�tO�Gg�]b�)Ț-h���'n�{�š�@	��b�-���:fA(f4 ��J�D��R��*�,�
����#�t��K��(�:�`��D������k*7Q��͈ew��!�����jS<J�Ĕ}�д_�����Vu�͹�`�Dw�]Vf��1��[��Z1�Vvo�1\FJy��{�|J+W]���ŷS�_�Ŷ>%�.�6!�����ϼ��L�ߔ��Y��<��!r��df��]71A��,�Nak�:ޛ��/Ä�Y[C��@�I�Q'�8���bϺ��]v	��M�6{tL��txĴ����sʰM�����b�,݀�t�w_�(:myTNkX#sI챔s�u(���N%����Q;y����V�-��M�z�(,M8��c�nN�V/l��U����p�� ��W�y�X�c�ts���"�))�v�r���b[8�<�&�Uė!���QAnՠpG�Ա�gv(�f��#-v��,8� {�A�E��Q����F��>���/�6ճO0Ie��R#�ʶY���$����8��1ך`ޯ���Ct�F�`6r���/H�B�~O�Vak�0&���"+�8(���H�n#����W.bE��z�5`���dU4����⏁�w

!�g{�c��e���T���Q��Qh8P%��*$�C�{T��<PZ��mJ|���U���^�mNBz����^��|��k~K����:�o�	��=�N����y(�DP�R�K0����p�c3�lS'�􆞿A�#r�������}U�����Rp���j�����I��:ĂY�Ik�0O��~�|YЀ���fMV��c](��^�*�F�ckZu�p��y�j[�(�OR�B�$����AQ�T�,N����m�:2w���ьF㬋.��4c����n!�{ɫ��rԙvI�"@:	�[�
�����.���I���ǅ�%����(.BS_��U�� �xj�!<�	�����S�ܒ�
껶bC��C�c���<P���C�b�R/]�#_�r�
��$O1���S���{�B��`����~�s���/����])L����&D��X��N��%,��R����BRxWN�*������B��B�o��oO���X8���ˬ������n�����ʁK����4�j �'��T<l���� �K��ZK��<�7��,f����1���F[l[�R1�1������q�#p�IU �=@j�.V��e��9y�i`����������?M=�:����%���9��K���o��}��X��V�ǯm.RzR��t��o������/	a�i.H����{�!It9���|�u��@����]��v�{O��@+^E��7Dsr[`�wl�E��Y�r��4_���(�"�#g��.���M-FV<�g�9�YY��r�3���7�G� s�.�E��lQ��\/�RS��D��s�OgTo��'�H�&R���ai�PQ��6S�L�NO����G&�0`�y�g�h�������\��p�Ž��d�F���q-����O�=;����V8��8����k�U���T�i�=���5�*�_�%�k�HF7�9����S0�L��.)�.��L�}��#	KڷC���\�5b7�&Rr����IW��2I�*��>�<M���
����l��,c�(�Dl5'��ć<��CB�f�@��J�D,X��/1N�G��ks�4<떕�N��ڍ���/i#,���t����5��+@j+�� .Y����a(s�}�P������4g��ل�h�e�`�A���BR`yQq���2n�� u�o�z�2�;U0�����5���"���A�V�ߦvv�wp]�_�bww����:��K�o���f�0�f���Z�M�� )ە[B{�rg����ͻ�(W�-��J�#��h+pB2
q�Ct�c����0z�)ۻFE9qYC	Ժ��1�^f�c�#t�:<�o�hKQZ��`Ts>=��|Ys =�$c���Ψ�v��$�؃~�
ͯ�%��z:�����w��a��w��?[]!�A���p���E����0��(�!�r��<U���$��l8�� �Kfk�Ȃ%a;@���S�XҳF���u�n-����1��1�j�]���f�~��K��A�A0 �)Og����E�˟s��$+b��s�vB�=��]S/��{F�4�?])����GLhhW�n���9vm6,���G���i�T��֥���@�4_t�D8Iÿ1�q���H���i{��睡fKߌ��JDB�@pi��{	m���Ê�������D�0W��������r����6�J��sD������ʊ[�¼7���\iD���*��A��K�`���Qj)�k�:{0��w��j�ݧ�c�����?ʯ�d�l��]�̳L"��ID�Nl|<U�����+jvuGh�;9��zL���φ�ԛ��B�.�;YZe�h�k�A�����ըZw��$m�~"\�&+�"�v 3�`�Eoj�h��.[�M<`��"�&2@����3)B�����
������{�
��D�'H�����h�`�|��#�ڔ���%M�>�(I<Pq@�9!fʋ��Y���Ё�[��^��p(Qİ{V25��D0��Ea�SJ����2�����}(�s���s�� ���Y��Y`�X��Z����^�i��@m�[}4����0*S��bM17S����C_ˢ�X)fh8p������ +	Y%Ni�@�:�oȥ�f(i!%IY}�����^��#�L";2䕊b����K�<�|ˆ3��lC��67���-���	PXn�*�a��A��L7Fۣ�n�̡8p0���\hs���a�NT�{<��T:ve�|/(��w�t�}��
Q��6X�}��@	�-5���%�1���'{��ɣOń�Ce_�v>�Q}� ���|��t~����(��t���E8��x�¬��s��*��˴��T���9����Sg;�J�DL�u�`��p��/#5�z��]'����\�]Z�5eR8~j���Dc�c=��(��ňrĉ�f��o���/3`E�NF��'ou��/F~.4�\t����zZ���"\\�G�U�@��s��
=��Q�
֝f�M!�����}q3����jj�mv��@���0Ǚ��&WR�P䥘�M��T��zH9ty�$���:�5j���N"�s��TK+o���W!.������۫ǖ@��>�����;�N%�~&�
��J
t�4,�֚��(*�:�W98[�8� +��RR�k���L�	|��PΦw(��\4�K�@~�+��#1Z��?���ˡ��D	��	��B؅��e�e��;V���]`�;�eJ�l	ۓ�`̊&�6~@�p�"2o��Yڹ��Lik��w��QjCL�I�g�Wҏ_Y�â��̈́�%TT����7�_�2o�=�|��@��O��D�2�^���)�Y��rU���|��w�e�K��o���$�?���DR�$-H<<_���m�
������l$��-i�OvI=����z��Dȸ��3*�}��6z�s[۟��ګz�n�ß.�S�1����Hk�W�
J�>a�S01�P��FY�'W )ɵw�jTj�M�&,b=b�cc��vYXOf�%�ݡj�1��K�	SxA���JzD�����\ߐ��u��Kg��7�w�o�:M��|�P�P.�J��c(��^�g:.{舻�{����z�^�i��T���YM�5��U�|%>��R�^_w=�NGlN����3iHa�݇��N �T��o�k�>!ɵ`D���8�_�w�=p���:��2���nN|�i�ql7���+�^�U��c:����D>]V���b�(p�����L,�65[��뢽@�����>���̄7���yǈ�75�O����q�(��1��C| 6��_�W
h'�Iu�C���̤D�nE�]U ��B�গ������)<��j]�M��1�c#���mv�m,��ތ��zu��,sj(역��á��,�0�q��j*~g��^�丅1Ծ���l���K9�HG���@��Ft�O����[wH�����`�/��Y�:X�V��q����J[m`Cy���2n�yC���A��m�d�q���|c!�=�~�?RR1̮�l���x)��kkZ���Jw@zp�E��=��t�C
�b��Ȯ٦�����E(U� Gˡ�x_.S�`+�`r �;�_Wn�d��q���XI���!�5��+��w��W�4қƯk��!1�-�8�z�1I���L����Ex���J]�Y��o�X%3�(᷸�:P��1�+�H
�<	;IH����W	7�jsL!���St���q���C
�G;f@e,X��)[�C���	GH���w*��Y��}c���Q֐��!��fn7��)���9n.��~��-f���}r<���x����j��[�>]����B0�e�rⱳ��
����ۨ�*L���ml���A%M���B.[p�4z����-�"��")�+R<�~���q�):Lk���'43��v#lGM��XJ�M;��%�0��>ȟ�/�����8�^���$�@$Ҵ٥� i�/����q�zT�j񷰶�-t��̋z�Y��rS�0S��@go+oV��	�27"1%�h:i�afAfnk�8���%�)�)5�]��|`=-���K)��O|&k��רZ	aa��+���A���
��Y��G+~�:��$��C�Z�{�����1{\e?�wv�ydU7}P�q�*}�T��u;BcJ�6�*zI�#֥DSa�A�&���v
$���j%f�탹��^ |��Οz� AAN��a!���vg���ܧ鼑�#@�	"�',�Ѳ�����:\�\�7��?�[^O�� 2H�����/�z�m [h�j%M>(O,�Ɇ\71E�"�����	�+9����5�ƣ�bV�-����pyjD����!5!�e�����M��/.q�D��4R�L8J��TC�YG�k��Q[�IpS����(�Ev"���C~�Q )�ו'<�v)�_I��Hn�T��F��Y!A�"�7���~%b24J(�>sT��j�23WP� �\��D\�@�%׵Xf�!�.!g��+4��4E�XQ�b�f#�}�
Nk�������&ɻAN�p�Ŧ��~���Ln曣�j2��Kk=��gڷGf){���ӥȋ����M�s"�|�u��a�����6:�����X��cTo#�_���d7�|ȕt>z���f��0���xH���C�.��^#3[�R�i�EL�:7�>c�r�Z2�i!�B��R�C�a����.�����:��CF��W�<Od����-��j[��X{\���.�\1��]�^go��#/ۜ���r#�wL㩿�/Ũ�\(�+Hoh��`����4R�G&V�!s�pҡṔ2Oa�!>����]@���:���Sm	�"�9f��ES�h_p0q��A�l�A�~�#U/t/������(�������$���0j[�/a,RS;8Y�$ry��w��`ӝ���Bj�L���"rZ?����# ]���A��I�u�;c������|�sI��-��\G0�%�S��ں�u��Yq��N�Y���Ȉ���7\\�+X_II�y>�5Z�S� v�d!�-l�� �𚝿J���yƲ�4A�G��۶�M��_9��9[��=`��+i'�x
�U�k��?��Zѯ��˯MM�)�j��f6�/�XF&|�09�������>�|}�2	�{�%B�n��o�4��h��0�.�H��s�5��L���^� �<ރl���9��"~zqg�����kn�P�U͏NE�ƚMo��*�� 6�A�gSW�[(��o��S����?|M4�2�:-}\�%�՞i'?о�d��]�#.|Vw�$��[�;�(�uĨ��0N�����5�їk�qԹ�a�M�-�B`ib*�M�[�E�L�.+F��o��2Ѵ{�S��M��=��(;P7�����^�[=P�=�����X�S.�e�Pʛ�s�}I��HO��Y�ɰ�=Cp��H��ؼ�%sK+7Ms�1��}��ڗ���˷����A�mP�.��!����b�]�B�u���TTY��<v8G@��c#�6E%0��r�pV��#��h�V/���t{a}#m���;��JM�����+���8�S����������n	�����GN(���l9oybk��[eN��}=<cY~H�����W�'zQ.@��`��4[m)$��S*�i#�{h�yw��snP��f��u+r�G��r^�*�V�VXw3����흹�*�%�"
D��꺼#��OU~���d�	���7�Q��۵=��'����N��RǮ���_���A�RȾٕJ��_���[g�n��%�ŁyV���l�'�Bl��ư��OڍN��k�:Z|O�/v�x�b �B��-���n峂'�}~�?�nTD$������.�}�Ի0�?7Ʀɦ��ߎȾҥ���Pt�~�/�pD��/}x&i�f�������hf�l�������\@}���_��y�MBkVQHLÈR^y�Cd3�㐑���Z�Ή��'bwߴ������(R����c�,�Ŀu%�.������J/�p mš�������C�f�j_~Z�(	�R�,Cđ���#j\P��#���آ���Q�s#`_��*�j���Ld�y�� T|wԚJ4-�F�CjKÄ�cy/f��
ew	�4y�u9?g���K�>t��j������Fޝ쇏)q��'��&��qP-N3�zyu�s�n��!���G�S�5�`�}�;GR��������x��4�5ksr�=>�'Q(���]5�*�Sc4��ا8T��T�ل�¦[�
��#[3�(�f�H�����B����*�pBų�x�q�zRg~2,��+�-f3�f�a��mSK�tU��yŅ��tX�}k���$',�5
7O9ί ��[a�e4ZV��+�%"���x��������b�
�.�6ۼt��O��;?�&��h��So�u�V{jR,?IG�u�#�~�|hiۅ�mAQ6��>:<�w������\(���ӝ����˭�X{Lf�Ƣ���PZ\���{f��ҷ
r5����7��dH��}YHm�Z��$���J�F���m��;��O�Y�\�)@k�59�`��B��8<�/(�,w�_8Ao*wql�ܓɃ�3b;e�xK���~Ἅ���>&S��z�b�x�`~9@r�NI���
���*��K�k�'s�g�אR�k����"m������=�<^����y^gw�圙ނϡ7|+�{��P��Z�'0�:#� ?����~b9g�E>W��]�4�1da�A9�7Y�5SOBO��g\��s�|Ԉ�'T��о.��TT}��k�:QzJ�(� ����� d/�B��L�& t�'�Z�	O����<�oG���� �3w0ݫ���]��q� �7����W;G5H9���
>�Xc���:����̉o$9�)ߞ��T�����<��S���E
Z���1b�p掸�b�	v ���h �oJy�#&�jJ�|(�f�E\�	"�M�uF~x���e�k��݋Rd���6xZi׀䫥S�v�q�@��xBI�*h�]fPs���e�w�3��=�4ؠ�xx�@|&�
')�"xF�p\B(���+��h�$<j�}�C�7UU�� N\�<<v?9�:��΋�<��yKz8�\�$e�Sqo���é)����o"r0G~�	1o����d� ��a�3h&բ4�������U��~GA���l��>WX���}�ٷ
�Ok�ܞ9����Uw�È��}-�Qlc;|l�h�I�c= ��m�]���P�o����@�$m*OD�M"&�OL�q��;�)�_Z������J7�GS�P������Bj5�8x=v7�4��=W-Ru,nd��Z"�@�