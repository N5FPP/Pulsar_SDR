��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�۫k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A��#��Hb�а~�g����o�+5FL�cu�ȗ$��ƃdY=�7?��ͩ�Ɵ'&]��ƴBAV� ����n��z<�+9������<�쨝�$;j��2��6#׾�9�eîᅱ%{�Տ?���/�gɤ�g�w���$�	C�Q'��/��C�cT~d�r��';I�d�?�i@��/����)q�Z��C����I��2�[�DDj�����E8�J���7�~y!��sh���5_,����?� ��U����t�4U�	Ē�����F#����Ӡ/�9M��G�N�	��\\q�GD�Y�ge��G{魖��Ռ�ٳ]_-3<Kx�R �>��:�$��{��������^`/�0:�~�P��'��	����$��*WeHH]h�}W���-�� ��ךSlQ��˷#�C[.�/�ټ,۷Xl��oY���������"i�\����~��3���s�,��ao���ܿiZ@,�RV�5!bAL����U��aK}��9t��[c��,�b��a����Ƹ�f[mӾ_�qm`1ca�W�j���:U�v~0pi�omo��/E��J���mN�;�����7�8� D�'|�n��Uki�6���F#9�q�@��*8�(�IBha��Z�O�L�k��di"��S�;��3T�袉��8A��:�t��}=ˉD����k�d��3�Y�zM I0	�z6�ߟ�[#XOt8M5'�y��e�j��`RTY���}�?;�Z�κV��1��`����B.��mw��l�H�au)�W����'����R>���,�$&����yD^U>F���K�̾���6�؞E+��/2�:�!;�f�����Q=�QF��P*�p��oۧ�H����:N�����}
��L�G�"\�
�i;U�;(�u���lVoS()9;��znTq��rT�Le�oVȺ��?�#�{�\K���k��v�cJ#�A68ʤ��t�m��!�X���T�{�Vj�����R�Ծ&����fP5&�-��F��b��w��߄�2�Ko��߽/9���g$�$J%�#q�����Yv�	U�)ڂز��N�ˤt��~ǫcX�I~�M;�T�Ͽ��ؖ��.��yv������'^a�TN),&�k**���0bD@�~�F<�Nv��\r�e��s���S��o"u�׷NH����9֢���mL�s�ͮ�8	$ݰT�K� �7_	y��P<j#����ճa릤����X�u`�gA�TY��
��uV���2��'�\^Q��
� .]:@��HN���z���Ǎ?�.�۩'��V�-C�S B�Qw�ꈋ%��V��L�����0����I:�(7p��c�f�j穮�/��Z����o�9벩�d�E�A���ݱ̮.�l���F^��@��4t蘖�%��+9D���Y���S��y�A�%�qyz+�py�x َ�' �C�:�!k.�k՘��;<&���Z��
>^�?��Zӿe!$��~v�r���/F"��rV��@id)�1���HF�
z�\;'(��jD?g��1/�N%�k���{]褉g.�����+>m{�V�m��� �UЌ��w�Դ��wE���/c'�`�������V*�� n"�DA�������^��m�SZ��q�����+d�;N�8�4!���	:i����ͷ�����ų��=�TT>��$n��:�U��}��*TZ߯c���Z��9�@jS�E��Aw
�nBVF��|(jI��!�&��c��A֘�S�؄e���x���䌇�L	��A�ՙn�m�c�� �f�R���?w6����.�����ſ����C~��miߣ���1S���8;������ �/~E�&0�$y7��)o�&�[&?�8ﳩ��W�~��_f�j����N��R���7��1A�J�z_��
9���8ϟ:����M����~�����ߐ$Hy: ��T�d�\�)�:E48ޯP�|;�XØe8^�m'�f��g��\��~�G�m(�J�����Go��`a�����#���{9-��8= �3�i�[�5�q�Zh�b� ��kD��{f?�r�����6��-����x�!��J���+au���4�|�d$ޙ��@?ܤ�dj��dLbg�*�*#�O6��T��pBR3�s�*��ƽ�{P�t���N���f��]@T%����Bԗ.gIG��M �q��H67��� w((���M���w@���?����>Q��GY�[�u��"��q�hi;U��4���	�1�v���NI�]Ƙ�����d��h5�gbQ��"zl���DCT�/ʠy��j	�=��8���d�S�5���3=� �p.:�d-���E�vӽ�ћ��]Vx������*�D~�����b�ӄ)�����h���r��b;T����U4nH2�z=<�,����+�O��X����5&
�Q�f�]����̙�{��!���(Q�q���-}���>�bc��]ެr�(�����BM��8y���
�E�A�Y�ҵZU� N/�z����Ǻ& A�7k4�2�d�mǅ����û���2g��n.�H�h��8�t^u,�i��;	Mɶ�]�t�1��*�D\N�&�~�B Ѽ�{�~��+��
�L�FHclt�o���æ�C-�6b����f����dq��O�n�45��z�>�7�q�$r��.}Q��)<Bw����Z����Ո%zE���Qjs�T$��sU�z����A\�`A"�xsMt�0椏�W���b�=��̷@����e q�ĉl�0L,�9�%���J):�l��� ~���\�*�=^�>����0ZSꊪ��}<� ]+΂"U����;�ʤNN�'HL�J�iP�<��l��L�����4��t��.�P�R?0Q@]��7O��G��n�N�#�'��ɮfBCR�Qp�5���_�nvQ?)&�U4��� �|��{:��/��!� "�=��w���s�^�dG�b͏Q��J,���S�7��}�fj*�e�Pw���n?P�e��?��o2�kU��Ö��x�kv��!�?��!Q&/�CEP�TZ�h#r�@O�!��b�&*����+�/s���a���I;���(A�,��n]4�S��A��<���}��N�M!;C��w���|6����id�)A��)?�_�#i�T��s���^�:�������]�-q+@T�Z�lg�^��\�k���տD����l��E�d����A{/��ۙ>�bu�����y;d��
�_�[%���1!�U���a��� ��O4ӟ�u��*C��CS���Ԋc�Z"f��,�C9|�;��Z�Ne!�3�r���D5]���AoC��m���l�l�3bl|˘@Xe�l�zX���\Mv,`Pa�=2a&;��2yR��Ԁ�r�9ד�/�S�i:�g���x�B�?��{q1; M_B����2\l�y^���}�R��gy習&�۸�r��[�$XI�*�(q��)�kW�ց��b�aR�jɝ0��\@JqmTk�r��j��?���89|�o��m��,f���4:H�/z"���I���B�w���)�3��� �x������p�_M�X�S]����f�˄P{��WN� �[��6��xLgJ�V����p��Dl���X�RCk~�æceA��L���9�Q��el�nm�oڍW��
�õ|q�ӄNz�eg�(
+��Q�7
Z(9���#�����vbj�;����'����N�������#�O�q(;�ꩩ��^ Bާ�O	�[r?�S�uE2�#�!nN��Ti�
�n�V��y�cmJ,(�Ц	(�^A�Ce��;f ���Sa��D��ٌz4_�٤���f5H�e���:��ŉ��Z�R�;u���(W�l#���	ۣ�����<	C9^����t%d1J��_���4��H�����(JJ�h����H�5�8��:IǢ���.�4��[��� �j�NE<��8������w NS���o��/�*9��wVY\�P$�q���𮥾����3��c�E�}=��@l�*DߣK��� ����w3�/�����_�v��k�W5�t��i]��"�j�U�� v*y�QU�4�p�VDNwg[d;ב��$#�^:�1�i�"�������}Kn�}�����g��l�jVV.�]�#+X���F��0��`�e�K<4��"�T���"1)��_����5�,�VS�����QK��L�e�K���z�xP>A�B`�%I�.ĉ<��X�1�T�U�np�e�E;6�0lpkȞ���mP�j�����z@z^���%�8��qq��)HD��
�ꮯDx���4�Zӊ��`�xq�.�g����~>����/�q1�o�M���Yq_�]�#�r�5Fj}�tvjLi�C��)W��w@��d��/�s�'j��f�>=��wE����T:tH�H�lO�8yZ�Q�%����o���o�(�����)���
��Gej�| �v0'%8�K�y�>���(1�:��/����4�u7�eb��ek?KV�7�F��̫C��q6ԏB ��k��W���Ȳ���ʩ�F쟛F�b�X8Ր?��ˤ���H�3� U��VŞt