��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY�Ɗ�����B��L�iD�Hi��c�->!*I�4���_:��L�Ƒ���&�{�ۥ&,%��p���8Á��ys�o�ȓMXˢ|~\�<�%-�RhN�,_>�"Z��Hs�(vb���"h9ʦSEe�h�1`��
��c0RyCV�4����1�^z��O�� ��צء
uߙEՙ.�$*��@�1P��ȣs�Xz
s-��&d�9����W�W����64l�o!����$�j����m����p�t�n�j*�;���2�c�d�&<hc9%R��8Y�lR59B2`��[;/S2R������-��[>�-�kԣ<D�(Zw��P!}��L��&{���`Ő�r����xD�
���[g�3�A�?�mtU�S⧡>1۠�PK��
�U�B��a��)�Y�_p����k�l�?�l��,��jϯ�p�ֺ�������4v�#�_�M��xВ�g�[�ᗛ�W�j��ӈ�V�����N\8��l���I�ێ4"�?�J�D���=�<�q��)¼��{�j#h���b����c��hs�����F��;z����� X���t �5��>�u$(� PQ����u�[���������w}	+��*�`�V*�6&]'A$*f<VXhq� �LO��x`I�f��)��/��b���ʖ�Р���/-G��@��oG��י4G��|~�@ۥhESNJo E��P�ܨ�uDo\S7@�sHն��^�|lT�'�Ө����3�_�%w�y�萸�1.��j?�r�pI\�bF��<����쳝T���HδS��{�w5���Sm��m������%8xhsӴv�M�<��@sMi���AT�D!7o�g��p~��ngB5_�����r��,� �	4��*j�Q�#�;v5�YL4�~�I�ؙ�g�s�"q�����p�$���EZ��'�#g��(K�o��b��gyk�Y3G��l L/�����C�����&%�T��X���w� ��N���� �Yč��c��N} �2}��;��z@��61QķV�7�Ff��J^�Z�B��۔��I�CLy�5�y �Z�0٭Fo8cO��D5Z&#�8v>-p;�'����u����s�<���T��Z�6� Ex�t�GH�0|��"iл����]!��Tɖ��h#�Iz�A�<k�<�r(:�%���'��dL�oL	 (�>�`r�@�b�	W0<��sFV�t��|;E���؈U;����t����u���d�	j�[� ·��	]�^:cA��Ŷ�C�;6�������;��l�e�=���T>��"�$�<��o���#�_�K���x�K�1��M�U�k	dh-�W�����082Couŗ�h6�J1���|��smA����%��ltV0��C�jf���qh�����-�|[ЧM�u���ٺ�Y4��5,%)!�T��ܽ�Bu�e�����a�{�T�b ��k����8�jɍ���"4I��ܳ������P^ƚ<	��<�4� ����Ō�F]u�6�J����t���ڛK,@M�uo�[wOa]���"7���V�2�O`�${�ܲk0��]��Æ��� F��� ����6�C�YV���C2J����b�ҟ�,}������>�P�ʩ�$L��3{�|.΅�a�rGnZ���3�����p��D�R��f(S�o�&�m,Nz���/��X�+��]a�Y���X�.���f��&��L���g���j�<���賋����y��+� ��[�h�y;e��壟qj������껫���K�R,�A2X�U��%�ш l0!�^�8�!����'�ksV}��=,a��,�d�]FY������y�'+��P>�����@}�l��⩁<���F��sT����rT�0$�����;/6a���!!�Ǣ&����țܙ�����lZ���n\"�RG�(^9�y&�_��W�2����i���[��nt��c�m�%ZO��U;K�~��E�f��I_ �}PGZ3ۃ�uf��u�k���v��Qvy�f���!)�F��]#�t�K~��vA����Vz�}.�£�*&7�$�Ԩ�:���_��mϢ>���k]Sѳ}��ۯ��_���k'P�u?�M��M�5�737'�k����Y�m�d���V;���w�J��	���nY��&:�&��~V!�@�� 3������h�/�P���L���&�@a~N�g32�M�q���,C(d�ژ�y^FJ�1�����ւ��TԩH`,��f+��6�?W�S�X�1�r�|6�d�:�i*���O�6iue'�4���mpۂ?�lv�CN�u/����Y1C�H���HH�	�q����huǋ{E`�R).�:�bH�8�����*��5%�?�t�x{vp�y3���h���V�����B^�{���wm�+�_��K˳� �\�K����8��wA �R��"��&�T�浱r��&��?Y��@Y�ݣ)��5	e��`9�������Iq��x���ƾ���5��\�QՄ��2/���W+p�e'�_�4W8s	�,�	4�"���q��41`� 1a\Eyn�w?ơ7ރ HX:>�}����;X��g%�T�Kc[�����qrީ��0�m��qh�>���t�7��ﻴP����v��)0�)��Z��`nu	�$���X}$��?O�R-ZJ��e��b���U�	Y�;g������^�֐���1�z7'k�m��x���㆜ҿ�Z����~d���Oƺ����M�I�5�f��\6L Y��J�%��u6�� !6A��sÝ�bW������C��:`���(\��41��R��^�_��?�dq�6�5IӇ
ɋH��$|6)�9�8��D��J
�*x�.�$\g��.Ip�K�E��!|]��K���X�y	$���������ظ��@�jgqzǇ���(��|<׾&��LlSv:u��Wv%/��J�u�i� ��&��tMjV�&�r���&�C!��z��n�1�6�Z���\�H�7 ���e4�a]�0"2T�K"h�o{�E��+�]E-�������V9�xF��vM��\����z��_�y۞,L�t,#�6�߇�a;��K�1���u#B������5��̘�)j��w�?��?\wN}�u���@��(�0J��W��b�uo��u����#I��]l�/�4t�mA\.q�q&�0�nZI^B`f�����Im2_Վ-���Z<̯�g1�!��T{�+�uQ�[c���/y����
oX��i�V/��TJ�Ҧ�����(V��X����S���C�}�{��4��e�p�ξQѦ	��˵��5k�(R| �>�)ͳ�[�k���3�O[F/�����j�[En�:�d7�BQ�t�jÊ��Z����1�*��b�O��p������A�e�ӧ�nX%�uT����m�''���q��D�4� �W�I�}����Qz�ϵ���8@\�-{���=�o|r����x�� l�θ�j� -rX�*��5��/)Ǽ� ��y�YR<y��@&?*����Ҙh�>t�Bf\}�[Y�����GG�'��L���{�"�:^��.���]bW�p��F�6Լwg�f�X���;�)��k@Y���r���a�cŝ9t���:��P�eb�0�FA�����������*�iY!�>��	$,������sk�=wC��Hd̺͂@#�9Fl�W^l��8�q���N�@����2*�QE�~���ˣ�g�����&���ڿ!@;	�	*N��n��{��n�Bv�V�[S�?"2���%��
1G�D���#�hVX\o<|�l�w'!�&�}���bQ��d�\v� ڟ���|���4���#ES��?ds]!�-ͼ<�E&؀�AX2@B���_�4gm!Տ�Y@���a���<֠j/=YȢ�]�	�G���1O��c0"Z%̵�}y+)���s�MĴ���烈q8+,5F�H�aC�R��iꧣɮ���.S�}O'>hf��͵������{�)o`��,�W5�����3ʟ
ޚR�	���Mz�gl���Ɔ� *�h��L�G�� V�"�PX�"�$��L���'Ȋ��G��]n��[ʳx�������%Oᐣz�6�E�V8�:K�[���o�����&�f���D�����:��cF[��[1﯂���p�`�0A~`ǝmS���4sȆ�� ��o�x��-�iW|p��t)l��Ƅ��@�T!G�95������� �D��0~��wf��jYd<N]uO������F�Y���>A�[;��8~'�Ѱi��1���ېC�\i�a���_�0����0�?'�kM^��+��%擱E?*+��][_�i�C�bs��ͭ�,�V\��Z31R��c��Z��hA�۴)��[T��o1Ǻ��HVK{�����а�fc1�C29�Z���.�ɵ&ù�2�~GZ��V�4,C�����T���C�Cι-*J�"r���
�b,^
:��?�#ZE�[q��<�f�����N��LT��4�]ҏW Q�ym�������@`#!~���0!�oR{w7���e� 6��[�8̵>��`қ�(�1�.���Y�*+���Oػ�,D1Y2o md�3:�Ԗ5R�}��������H�� )r`����<�>7��|IX�@c"q��C��K���^�v$�K�N�+?f0���,ɥ^�쫖hJ���Pi�A�����V/�� ro�\��ij��P7w���H�����"���&�Q���`_��:���~El�k��=�����rO�����<O���e�xƚ7�%t����͎t�"�`�d��v�ɼ �4�!Z����HY��ş�O {x�&^e�	:C6�ym($�Qg�p� kjC�M�m���8�R>�5ve�j��F�"�/5�eSm>���u���!TE}�����z�k���Б�D��?�u7��E��f��W�J���!����d�o�p��͂U�=D"�Z\��7���_����$2HC(Q�Q��˅o������V��~��\i���X(���6���O�g�S0�p([�[�����H���N���C"�V6.�a�w���r  ��;56{+Q8ܰqTB������"��M�k�ZN�`7؍
�y�+1I�l�t;
�02��.��@`�x�S���Hu�Z��e��a��@��mU�`��]pliRt�V��se�sd�	H�$Jȩ�q���v
OjM�����h9���$�w[\��ͮY���1���������4K�8ہ�w�����7W ���4�[�8�Ô�v�՟&�A�s��ǲU؂X�U��
��a�!e�ȦL� �ʲ|> �\@W�F>���-���笙'ך7�I֓ۮ���nTF/���^Љ]���C��>�`��Z�؈��'{"�vt�t��6�͒���M�%j�߫�Hr]���y�	"�Y,"�WW����ԍE�͌؋eJ�5<iJ�K��bS90UQ�ٗB�7V�U!�S��l�P�?�v�zA��VW0NK@�b��Ԇ���]%��*�`���[ϋ4�oi�	��G�B�b�'�8#�J+d�kP����)NZH��>��{�h��E����C�G���W(ם��62:0�2�$�m#،��u� �on8���b�/�� ���H��Fq��a���Aw%R~����9\��u+�3jB�`#Ɉ��6�=���>���c஫?;��ց����Z7"���	�:�e�!5t�8�QE3��x�jTu,2s8����K�B)��bM�8�Z�+����<d��d�n]�F-��P�FS�ɽP�=��w��vɯ������AU���l�^�coZVɂ��YH��,���'���:�P�Ԡ�����L��?���msxgB{���.�g�ԃ_�w����Z��?M��3jJ q��P��f��}�ָ�iۯLg�CCK=_6��ϩ>�k���-�=e�g\4��<)�M��OU�*�b�%Q]�5�ك&Q��F�3%){��=ğW=>X>ny��D��(V�&�=�y;�l����}8>���=�J��Y�Bx�,8����\t�Ǽ�M���Y��>� ��4�K����Z�1\z�Z�*uCb�KTI=��kb�O�b�F`���ƣ�3Xt2��P3��_�\y3��+6߶�p��ٺ����e��bE34o�(���չ|����°�~f�q�?s!Q�5������n���]��N���>V2^��*
�!���2r�92.�|�]y��������Nҙ.�YaX�w4�5��
c����A�A�5.1��&�U�=���cU�Aq�8��0�A㗳����6Qdke�Y��yνw* n�q�V0�`�5v�ذe��.�[�&��걲*��j|����t����`��-ra��S��K�E�5�1���^$\�YȮj��9*BjA��x1g#�OA��X�aQjT���P!a��8��[�q��.!��#��Bv#��r��_��z��h~�^���!^�z�ꌄR>��B�����TH[��Ѳ�z�������e^C�M��w��_
S����$<���'<A(��7A�x��	"�-d󦭳�H�S��vJ8�Ez��C���.;G��<Ӏz���	�Q������]�˖�������+	j �Z= �H5G��O]��T�
�?m�!u�*@�P�$�u%�d�fk�h����y�DlOpj�2s��L�q���1�lPnщ�� ���jN�Vt�2��=�1����ŲM��t�V0|��5S	�^	����5�'�����s<@p
Lů`��qV,�J\R�|êժ�f/[T�P�D���賂��f����x;��)!g�u[�ʿH�:
-iY,�S��\d
Z��z1p��+B��
LO��
g�`�E�p�n[��\o���X����.1F��2(���5�����Kv�b�e)f0�r�
5�SL��-�R/�p�4����!�a�����z��=j���.���gŌ�#�X�V�\�p����7'����.	��װst����*�:�؍F�&Gҥc_�����s�	�4w	�0���k�"{��ɮHx:�N�{tkC&��)y�<XMW).��U~�x���8� ���d<���h��Q(�O�?G6G�]�������ȋ�����d�c`�=_��j��RqE@p��3�_������ǽ��:DW]F�M΢�[�ơqe�T�_ۧ�1���9�K���]���9%�qp`���G���ۤ��i}pLR��U������_�e�[�6�T�ͅ��/��m7��X#h��7=�z�kk2�BQ�]y!�����.��+��.��'�b̅͛F=�e��ߵ�Bǆ�24�e�>���E����a���ә�P�S(�si0ތ�lC��OŹ���3p�9����*��8�R�1�j�o�O$GpW��(�X(�ӓݟ�q�j�b�:ľ���Ї�K)��̎m�(9N:g����r�7ߋ��5�����߶cL��YQ�/�T����lqϒIx�!��;v� �����͉���&R+�������Vf�"�ӝZ�G�-A[���\_J�Kf�q�0��h
a��v��z�|j�dO甆��1:�F=;�P�_�eau!�8��n�6	�Q# ;��:��:S3�B���U��釘�z,=��7��-���/n��Kt��m���a9|
o
막���1H�ى�P���6���@i:�"��`*t�|xm���B�����X:�S�����>ؤՀ�nÒ��4G��4f7����*��q]��8�l�W1��ƹ#6��$��,0�t"��H��x��I�,�6�����rnn�ӌ<�G����R�&�iZ�>z�;�/r���uW�솶�3��m� E��f�i$N���*�$���^�Hꁉ1�c�g� �e��<�䪧ٸv�k�pꋸ��'�fq�m6���`G�zR�J9�d?]�"�O��w{���P�9�9a��5+�I�1*F(�O3��Lr/��YWr�մw_cw��[F��3�_%�ȑ�4��+'&�4K4�ٸ��
Aى�2z	�����Кk/0���TT߯S���_E�$C��k*+OCNak�>�Eߝ4��؏�2�}���I]���2�5V�ŉ�!t��n��2zl o�o@�w�ގ~��?f���?�VG;c�#�����\y�vNU�;�,%�-��7{��yXN����k_��N,#�p���,ɸ� ���4 �z.���bbP��IC���G���]����'�T��79����{[b\�x������H������ڇ^�d�� �_.jj1pPƼ/~hsW+��LօR��5��^���P��8���}��J!�r��M��,Wf�/hEcR��n���㝄��Dҏ��JkQ�UqsS�+R\j ���"_�ƣ϶���0��%QNa��v�U�H��K��!I���[������#}��5^Oh{��}簊aK �M�R��F�X�v���\u��ׂ�.=�|,��lu!Y𓂺u����W�m�+���ԡEJ(�5�e�޶�p"�W����C�a�c�?�/��v�tH5$��;�B	��℣t����"���G ����E��r�(6�sR��9�+�w�w^�J�!a5�D=��%�NF�O9I��x�w2Mj�P͘}X�R����J����ZzVk?Y������	J����s�e�#]	�dХ���$��)ʛ��vW˒#��9����P���gO�^r�qr��⟀�����)��g��s2�,g��6�D�wD�3t�f
JaD>`��V��%:�������j��