��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 j���αee��X�@���
�M�p7�O� ��`�Epvm!V�U!V;)�����e_8u�F+wy���\����X'��Զ?C::2�5�%��RĨ�/�A�M�Ʀy���*0v��ut�2��<�����vU	�v%��v�I�j�L������@�@���,�2&��6֓�įj�&�����>�nn*3m+yp�.D�G�)�	YUO��	/��)Ym��Ef|�m'R���*���s�x��,��f�������))���k��Wv��$���։���,g=�k�E�����=\Pq����ʌܗ�?%�L1��;1;!��u����]�r��[ܛ��~ �iwl�:8a ��t/�غ&�����%j�j��zV	��9?��4�+r2�������C��m��ֱ��V����c�G|ߤ3v �� �����/@;3��3�����MDb�)��Hi���m�,�<) I�G̜k��;�7�^[Sh
9��#��!�E� ��P�|F��֞��0�#�3q�,y�,��q�2
R���61��l�%�����Ǿ�m�^�7�;�5̶
rڻM��w��
<��q��l�^�#�-�,����$�������ή���>���,Gr�䏉G�P��(��ɼ	�8�;��s�����!�`��Ѽ���H��>a�MUP�Y�۾/3y�e|� G[��������+A��B�,!�t��f��t�%�o�gb<RUf��<&�4���p缃�5/ӷ���o���^�v"sG/���)��w\ގ���Q�zrk���F��2v'�5smː��䉲����#�/ۉ�.�+n���e�WQ�i;��p�%�bw���2��m����l����?��t3)�&��~��[U���yZ��ZU<��
׵��Y��ɥˏ��_��]������ )6U��:�- d-ǒ%�u���3A��R(�3�F��S� ?�|���x�,�iڐ,k�l����N�x�DA>�3���=��.Fi��O���k�9\�1I�����&������8�S��x�St��akI�!�2�`rF�k|�lh���z���9VV���aH�I1	�t�e_CŎ|��债��鹇����qa�G'�]��%ev}��L��;'&V�ߠ>?f(��Cm��&�:m@�m�u���Gi1�Y�=��GV�!;��^6�܃�Ã��"d0s���%Rd�������(>�<����0p�RP�Os��]yH_I�	}��Y�����K��SCN���q�&zBpY'̟Q�&�1��S}uM�<�]|�Ĵ3����c���`e�������وTb}t��0n��Zk����&�ȓu҅J��q�}V�9������9�D구����X/�|��*����6{�T��"�e|s��<�,h�F��2�R��3r�qu��}�ܘ,���,?u�K8�)��̫+8{)(� �m�����e��v1e��a�Ve6},͐$U�����u��K����ۓ��ȿ����WPޡ<�{|�-�}��Y	*X���:�#�ȟ���qP��x��2�C���t��.H�IeD)��'�	�w7�J��Wj�%�7�~/����<%��aݹ
_5�M`�SRH�$~#����$��TW`b����1pj���Ɯ��7��H�9c�
���[)�RW�qZ���ĵ���e6i���G �|��Y;��ڋ�=~��;���%J-���Q|�$hԃ#,���!���^߶�J�C5����B��|^�}k+�z��T��&��0�@2|ͺx��yEc��P�:/��L�����l��n�*gۜ<4eˡ��3��c3^o�8�*���3py�ң �����y�W�uGu�>H����L�=ݗ���n2���������c`��80y���Q8��z��U��By�>�`�Hlf�Gؘ�T��.��?ߟ���[�3��;���NA������t?��t��RQ���7��搵�ZH�t��S-�E$,�J�<�!ղ��	�} ګ�!K��1hK�K���Ϣ?2�E��Z�)��u�Ttr��p͌�.�7� |��N�.L�>���c�aEk/�A���Y\Y]b�# �{6��u��Q�DI����i_ bk��b�W:�P2ȬڻH�L�Y��ߔz���\��&*���S.��D��y�l:�w�ڐ����F�1���$F/c��6���%,a�F�QS7��Z�������{�0v1�ôQ4c��Ml���xr����M_j6��7��/�1�9�_���6��߻��<��𙉨Vdc�������(Yn��S��}�Loܘ"��?P�^��� �y�p)��r]D?��E��e�q�!5��X�Qm	H�;��� &J��vCS����Ly�~�f�&�ҝ�-�Kc�Z=qw�J�a]�("��C�J�'��?r&N������X9ܶYPd�*�#�	��c�W�G��򬫠):���qR}N�j�W�v<~{��e]Ik��%�uJ+��'��HqC%�@�XsX
*	<�_�;�MM�[�8!|��"�݀��AxȸA�}��������I�0��6�������(k���LM'#\�O'�R���O��|�0g���:/����_)4U}�P
�����%�x�gI�CÓW��C2������f���pY�\Oi� ��	Z4�Z݋ˇ�j��+|{��T�����E��ZU��$�V���W9w"�P�tB��Rn��X~+#u�[XOOu,Px���eOJ��mG�Gj�ɃqP�.4hu�c�q��ӽd�>���%�t�G�S'���hX]�su<�8��J3nH%��FSco\����m;S�e0Ӥ,�6�����1�lp�Yhr�W�+݉P���I;��:*����!4�Ȕ��qG�#=�z�b�'H�UӞd�^V��2�A���i�s̆n���~���yy����و1�m��~�A��n�:�o���D*��oy��5n�WI�؃�^n��V�Xj�no�'��md�e����./[� +�K�S	*�?s��'@�����r��*�ݰS��Ǡd��KZp%�{E�]8�J�>�<��+��u��薵���� g�=v�3(8�fJ���c�{�`�w�Tav�!�]��������]:}�i�t$o��O�ⳤS�!x+dE�Ri�]AG�#�h���թ��P(�UN�h�t�iT�v�+��U��Z��0N�~H�+R����^��<�C��!S0����O{�~�ؗ�6�I��hn� ͮ9��9�K�h����!G�9��Gf�-,��Υ���w$�$ ű�a�X��S����[bpa2bW�X�$���qx[�� ����n�ln��§e0Y��)'񸫝x��-���~�q~+����w
�d��Ú��O�=�Z�]P�.Lb�^w�O�����[��:�,1�)Ƌ	�c���6PB�ߚ�@&�?�+���G(����C}�p11=�!�g<gH2�G
��3M�5��l ��m�:�Z�x0�H�N.f?�
��Q����e����DՒ���
��]��F�̒=O
��g�F�Og������u�tƘ(��\�s�Rc։Ǆ��M��^^א	|��F��?� �q�:���� `PC;Y��Xj1��/v><g2�݂�v�����#�\��@&�7�a�SD�IQA
ܦ�ah�Ց�H~�(�	
l9	��[����4u�
"�q@���Mf��!H��P�d��-�Tp����3��2�l��7��л��2�FO�լi*K.�M�f�u�1~D�Xr�F`'����<<�۷=�^��>��ţc�BEb7Ke��}�w�FS��,��\8\J�|El��8�,�{�NxCv����/�ܛC(�߫���;'o�"#�NAB���:U�Z�G���/)�B�r�R�qb����_&[�Z���drh�a#�� (_Gd0Sx6U��P}4�w��`"��6>,�w�t�f��s�9z:!�f����{xy����D�H+�����P� a��\סq��e�v`�yVV�	,@�í���̴QܨnP(4�#.iEi~S�@ͅ^ˮ�'���8���i��|7����R�Wܚo ��$���l_���`O�d�Sde�kIV�|(S��k�Y�8"q|fP��U�jk���iĀ{�\8o!�mh�'�0/��a�;
�ef�����- ��^�Pa�^�@(��tc��3��y�DNx{��!��d��d��k.�e�Dȯo>��F�!�c��OVz�{aw��Ju�� ��C��y�|�3�oَ~'^ �N#6E�X:���٭bA	t��w�Ȯ�h�� Y�K8gp�oXu��D�����qI�>aѧ�Gw,̮H�)IS�8>"t(�E��[���$��y�.�Ґ�P�h��dk���bU�\��=�`�V�P�?1�B�H��s�I/���#3w�A���Ҙ�)j��-�2s��:Y��_ᙝ�"��[\��lbaS4�_��k���%S�\�2ڔi�^'����'���͙��()�
 �︯�A�E�.��x�U��x�bO	�)�:�le-ƃNB��Bye�Nצ�Q���g� K%�0kU����1���:��]�&/�	�g�L�g�ՋZ5�u������j,��&+�B���	�H�<i�l7��W=E�!��3>*^B"f�מ��g.)��m�b��:�1fV�����7�X�r�z���3�Yv�(T�;2K�فXo�&��{&�	����S;��%r��#	z}���5�Q����gVԱ d�������=S�N's�#'�)M�q�'U�^�k3�l���:م�!���7r�&�x�BX�&�>	��9��X�Z<��,�bRǷ� �K�\�[����̑�S���7 mO� �L@��w@�&Y�|�L�96d@��ABn2=ӱ[J� \�)�����Z��^���،p_��c�"���`� � m����h����d�EZ��7z ���ΉI>E(��0QaѦC����D:z�[L�z� ��3�Yg�C;�a���B�����w�vd9�ŗ����<��G���*�M�T����Tz�)��k����C���c�s�L�S� ���az�hKԓ�rJi����g�
���n>#�;��%�k�*S~>�ՠ�y�Pu����fvۇ$��H&��{o����]�u�:�1F���fs�{m�/aoPǲ���G����G��"�Ge��`�N��+��V;�M��PrP���l�X�|l�P��@C�~�;�ٟ��gz.�pB=��UeZ����H�NF���B��k|3��\3M���º,�7di*�k/e�@32�bZ��ݓ�B��UsG�u��d��ְ�{��%3�D\�a�'[��|)xT!2K/�	�\{�ūvy���S`c�q�?��V4�:����	D�`@��o��ZA[�P���b��Y�7߉%��Dm��I[1mc�W�o]�����4�R�o	c�(;���8�����j��i��[_Ȱ�X��
y���ŷZ���Z�ܕ��6@X�\���ZE���V�1�=/��R_�9s�)ڤ�p[*.�����mЎ�^z��1�q
��J͎�_O�WE��w���a쪌�6��,�"�cafzs�D�D�~ظzv2�C���.�U���G�J̐FL�6�!���W�=�ZTlZN"@���L@�Z��tCt�ƱNc�%�{& �LW��W4��XF�@m���V��	k�
��p � �`.:��U�SZn�^H�7@UmG�e�vI:��#��@uu
?#GO�QV�����4��]����}��ؠ�{�9ل%����Bw�4gJǰÒ{L��<�ǏM��G9y��h\?��V*m��n�G�~��H{�YO�g6����B@{�MȲ!�R��2�,*?3U��5�dAj^PKF~���^����&h�Ȅ�DY����N�A���b�#��� ����\_�;�.� I���"����'�_1��+gP�J���l8����(礞)TYDv�J��g�k������!��H�A�	�����b����C�.s�q�V���/ʹ��b�gٙm�/�a8�ޠ-5\/jot���>�U���G�]Tzl�p˹F
BD:=&
�y? hnY�ä��s��<9��z���7ԩ�̅���мi#�Hh�ʋ�=I�1���G^��`���$c�Ol(d�_L�����g~OV�|&�PY�`Ηw��<G���A�e��vN;�&��m0렀��^�1�9����2n��G�J�����,mg��j,/tT(W'm���m(��N��%����#�M�h�U��ﺫ���X��2xc�U���y����#�N�U��uO.��Jh�(�S�@`(m9 )�]<2����5l�:&���?�|F��$���6AY��E5���\����ɇ_�1j	� ɧ���BB����@i�任���>¸[5)���B�����2�H(��&������ ��~!D-���ɴs�b�՗4�t�GPӊ߭�,1EzC�ϛ���"q�`����t�����id���,��F�l����� �83����&f76�����dCը��0!aQZ�J�'H�L��t�Gˈ�[���6��xmIw͵�Q�2��p��'�M��	C&��YjQy���1�v������}Do�̵��w�'���8W{͟������v6��Ź0��� �.^�t��SzW�&_1�98"9+e9�@���(G���ʲ�*�+��>���-&�L0j�)�R����`.ß����@��8w���)4@7�²b=��\�5g*yz�wmw ���i�j����xj�[��d���ʄ�3U�P�@=�+瑭�����&X�Ò��pW����C�	J7�M���Ӊd��y�9�j^e��X*��v��;�"�/2�gh��L�S���ݰ9Q7�m�z�Y��^�fǴ���g��6z`J��)� 01�|�1'�]������.��6�7�a�E�o4߲5_���s+FG=h6�y��rJ�IY:���K�E���L�Y_G�cl�=#�yO�1��,:1<W��M2"X�\N��Y�|�;��&I��ir~�*
����^ݖ\�\�n�jܠ-"�}t�B"�rf��/: �7�|�H�J,-�w�j�g���C�j9<�c΅zD��I��,�9Q���:���o)ik��ߠ��ξ
��1o"W`c��QCj��3�	Zb]�@ZrrQ���C�`U�ah�-����2�$�>K��q�?��k�>��~�袓�����t��V�?�È�mٸ02���܋���e���R���\�q[_���
�/ �5�-C��b�eu=�9G�(ϐ	��2���V��g�\�]�a�	�^ťG�s��3u,��04�CkЈ��:�K��q��������	T?Ԓ�x5��?�p�Z)�U���9�!o�Ƭ�]�-�rE�b7Ϧ)>�L.ה��ؗ���	��9����k/M����R�h�3��e��q��'��ټ��8�G�������.�U�r�|{�����lX9V5�	I+X'}q��v��p�t�ox-�7b�xJ/�*kE2N�2lw����[#IoZ���U�?;�s���K��CxW�F����NEh1R���X���w���0a��]�Iw���Y= ��E����w3�;����j V��:i�c2Q��������X=�!1��mGH
� ��jB�i���.N�IT��@��\ �8�q������~'"x�4��7���r�k��>�#��;�k���P�nv��o�X��ᷳA��v_������c�\���E�L*�-a��JQ��8��[~hD1&{�Ey�۬���ġ�l�m�3eoç#��V#*0��;I2T�2��f)���y�M���B�(����a0�^�P��h�4���6^i��	��Kb �~㈆0<r�g1&�#77&�e�@�����1�<��`%�:�g�Y���+s"����߼�7�K���t��H�E�ҊpI�q�{.h��GQK����``�ҟų���6q�@���H�\����e��ҍ�1��8�#�.���Ob���&����Z�\�#KG����k�Ї��!� ���[���bP�)�x}�]e<��M?�Z�.�ъ�[vES &�9Ӓ-�J��%�E���^>�l�7NJ��s�L�1z;��kc7�����鱪�	���\x^�1B;�t)�& �����C��T^��Xa|�x�M��ZM��t��E�ڰ��B'>调ܪ���Ǣ���Y�-��t��c�Ga\|P(��<;޼�*8I\3��!�+�������h��*	g$J���L��>U���(�δAܨ�Ԇ���mw���?��
0'ѫ`��Rc�\�Ah`�a����w�Bvo"q�N&��Q����~,j���(n�|��o�9L��9�O�2 Ʋgf�Ym��y���&�;�~RNñ��rP-o�}$+~@c]��#\��#O�>�&�]�*�����Y6,8�c߉c�
Є��S_.�	�l�h�hm����\�.���u� N��T�T섄 ����G�>��[�z�B�v�&�sL&�����x��<�D|w�!w����/|&}�?�\U?�������4X����f�g�=NUօ�{t6����)ZQ�af���+!-�2Z�L�K�Gjt�w�`i$���!�����wi^K/[@�����*�s��,��������m�M�D�F�L�p��N���㕻���ػ�H�i��wp�O��X�ى�yѭ`P�$�����O�h7A��ۑ0Vcq�������,OL�����j���km� ����Uij醃_��� u�7�B�drZ��_i,n�k7"�oɯ�;�8�R
���kΥFg���������s�%Q 5ގ��[ժ���4�u�=� f��k:���#E���W���3�9�H�l�βR����9%p��̢�1� ��̛���;���6c�(H��a-!×��&����"���6��Շ�5��`����9nN9���%�X�=�tʸ�0&��ëH������c0xؙ�i�r�}�W�RP$G�^qX#�$��`s,#�M�,q_������������4�u��C6��
ȑQ������Ŝ���������īSu6�q.Hˊt�a;"����	��@�O�T��~�[c��	^�$~�8�B��Ŗ!����=fx4�1A�(�e������b��A`r�L��ՙ��B,�׃C$8�f�,}�%�)��⵼j�_rU�%����l/�l��Ⱥ�I ʵs���G����uO]7`�w�P�3~Z�m��l���%ֱ�};R.;O���T-����=�⪚��-�ͼ0�&�PI4�p�1{9C�r�� ��aP���MA0�c���&�3�Hd=y�����ZR�y鹍�(-q/a��px��v��UV2<���
{�[��HY��6@tH�r� |a��T3�4�Vd4 ��#�G�V\��ԣ���#�y�I�����:�HP���!�ۼ�Q�_��l�z�Q�~"�'}�8�kDq��1Ν%x�^�뷙O�x�Y~?H��ҥ!���g������@���o���7�M�d�}�0���TP[I��T4ȩG3q!���O����ԏ������h��p}L�ͤ�Sw��(�!��sC�F��.G�bh�R���+ �GIZ�Ш�<>��ro�=���}ߩ�x�G���S�L�~0F�u2��,����J�,�U�S5&H��z߷�3*?�qvX��KC�G<�~�h���
�-�s�(��cgsx�7�DE1;nBho��T�]h�A�`�璝�a"AB��̢��jH������u�����������6��\�S�,DJ���-� `�"��ܘ��r�h�؍D�����_��JcIr������U�Q�O����.����!L;}<U�/G5�4�I̪�Ɂ��p�Q�lњ|6����+�&D	y،�Rt��O��F��	�;�����H��2���c�Ѻ�Z�eZ���v�XΟ�Qd�?�$��(b@���01��szP'�^Wh鲼%�`T�$A�cqj]�îO�ʹ:�赬��z�(�w{�5�OPJ���n��+a�L1�c�l�e��T��PP� &��X���e�ʓ���_R��n8�`4�:��@q	���=�o���N6l/7Q���vwr�lS8v��<l��Ǌ����&O�r?Ю7��HDy~S� �ԝ'��������U�׃l�w�k`)���[y�@R��2�Ae��O�̉�[t�0�8�� х�Z���x��|L5�J��&Ť�u����qJ�tj[Ҿk�� x����i �i�C����o����4���t.���%}XqK����D|����9z�|���(>ȴa�M�j���1V\h�;�~�üI������@�ز�Ӈ�6/?4r�!��~$�!*yb�:;L^���W�<�O�V�*�,�G|�6׀;Qol5�ZQ������R����^n$;z����I(�܄��%k!��+w�K���Z1&M	����#��ۻ�,���&�$T����Sٟ�n~ג��9#P�-���,\��Ԇ�']��;��������9d^�L($ޭ� ,<F0_Y��I�[��_�4ymt�p򉆳kp���ʶ�U���M^u��-���y�C�����WY� 4�z�P���Z��R�cH�JK����wp�}�-}�<^�|���{�2�**�%8�ekȭz�)�W����ǋ�D���2*r͉<ZE���6K���uo�'�Қ�'G_ļY��C,f�̲�g'Et�F �ʪ��,`��?�t\����[�����xϧZ�1�&�ޑ�׆$��1��^s�� ��T���A�1,(;�\�o�٪���au�O�V��y�- �i��q�k^�]���gL	o:C��IK��gW�j�<�L0���+Ez��u���Wn�Xc&m��̴)<��'��Q9��?#%&)g�wE��V*H�˘���Z�tU������ceo0����LR �j�N�w���>J�j�
�"�c����Ofo;�3��`F'������ \����ol8HN���3#�6S*T��ls�e����5���P�����MOʕxf�v�9�q�-S�.�Ge�a��$�	Ya���튕$�@���LeIa��s�&������3�Y��{p�U�iE8���p͘�:���8LmC8L��n��M�#|��t�s"#tVJYq���a��N[&��1 ����_�ŧ0P0��54/ID�H��#jf��1l���ǘ4}(��`u�b�oe�
=œN�0J�vc��!ߦ �6�aH����B��#��ܒXN���g�Zp�$����o,����lP���T(�I�_�:��� Ӈ色�Ic:)��Y��qN��ܼ��L�$�W�V2�-�\{�|!N���I_��'>N�3���F�S��8#�}��)S�\?�lOp�,�"�-���V������tE6̌�ڀ	%�"Ċ��D�+���
�e����lL�aCS�I��@'�C=Q����\�P�3������i��Н���
9�Zt=�[ۤ�-lA)X�P�����&X&Ӿ�s��s����5_�U'w}`�@ :l!�F�f�~��t�^y���n ���ʓ��-�l�I�� �V*��A�Z��Qo��5jM�}4�ϩ$�0�Z��h�$)~�EX�W}�P�>I���`OC��$�'��ρR��(f
����8�h�ģ�3+�D��cM� .S�xv���@^[�/�x�.D�,��)�Q��k*+�y��n�����le/�e��97�x�,u�kDjڞ�RP{�)=!�MkY�Hn)!>OH0<���H�-N��H�愲��#S�N�s�t1`�H^��^NIv|#o�6�L�Vד�YA�х�Ś�w*T�a�l|��+�<�$ji�Y���Ô0���S�m�9�[�%�B�M�L[�S�]sƋ�u�Aڷ�ӡ�wzTMI����Q�h2�B���>�n.������<���LÜ[K�b�+3��V��,���q�^
߄��;���d�yv�jh*/؈�gA^�S�/�ͽ��&�4��t����Z��s���:�DӴ�D3Y�@��v��.���Ңl�A���i,��TG��0��د� ���j��x肱(9_�����
r���:S�+XE�~�����}�;��ָ0��,�CO�]��}JQ�K�l͑(�ɚ�^?d�"¤ n��>'s�
Г�_(��X;������"�H�/������K��'<���QL�6y��A�ͲX6��ô���UI�9��8-�SΕu�Xmzc��l$�of=# �1$5�B�.��r�r'�BR������Z�g����L�-�4OD��}	_e�P8�S���k���#�����C�Ƴ�ұJL��{����\��;�S���/8�?%zՄ���}��^c��4XĞ�p��U�Or�A%�y�?�ߨ_����"a�B����yjF�ڢ�Tnóv;�P��h	�F�Y�����$q=`�b^ɤ�I�ΰ|������C�O��g�^o�}LD�M%��yk��K���A��
 č��Fz��Dq+^)	��I�4�3�����2��+���?��B��~p��s�?�ʘ6獏�Qwܩ��1�>M~ (�<�'�0V�V�b�����C��p�F��:K���P���`>!�p�$�<��{9�$=d��v�{*�N�K\��[���Ƀ� Mǖ޺5�?"�N��?.o�Ȫ�<�7�0�C'l�N���J��'��藃PF�X�����Id|�f���A��������S�-�j�R��:��F62u)��r�:G��%c*��N�$u�z�KU �dc�z,P��)�gC�bi~z����U�bc �2
3�����C@����3I����iT)�&P�wtF��Ygld��3|ҋG���x���i[x)a��׿��6,Z�j'g��:�<�����/`2nf�5�ws�ֈk��R�6yF���pT�/��srѾ�,x�0%%����/(
j�vDS{��\ߔjr��.��H,E�;;�ؾwO�ܮEH*FJM�$B����_���vǗ�P�k�]R.�L�Wͥ�G��w�;�M�G��G��[&�3��]L��D� ��}$X�*Ӥ��_��S��\Nb����L���w^2�Dj[�������I}K��������,l��ˌ���b鸦1讹��9)���.��UP���_�H��R�ݗ��9"-d�m����m1��������DM����40R�)�۫��6z�"������֕�O3q?{�3,�~�{���I��DZ�$<� ��띘��! 7w?�QtA��c��oh6�R��Sa	c�-������9c �%6ޒJЋ|U4tz�w�a�p���h�Z�l����}�ʯ���y�|hW��V��/Вb R0��F��˟D�=Uh;0i�Uǥ��q���$�,�Q��IEq)���$�2�x;v��#(���5��g�]mfTX����g����_+~��"�����r�;��r���/Q�68���ey��a��*�H�J<<���@A�xR����f�/�4����9��rlE�n��2v���2�$����S�Q�����$�'B.���:>�?�{2�~g����o�´�9A�v�æ�_�:�W��@/T��R�G��8=�=hV;E8^/�󍥑�G��5�?m�zb���<r0�J�<�D4����"f%7Zˁ&�Ue�,`:�ji7W�h#z$�\�r=������7㏯�kǂ�݁*~+7��kʽl�ս��y����=�2�b�Q���zK]�N���{kvԹ�G�8(:�@?�ZW��X �;����f��>�LK�I��1%i� �·��ObAQ7=�(�D�%<ɻG���Q�	���Rz����Qap	 ��j]��\!�wժ�������I�!l"��\п-�L�:$�ֆD�<���iN�!��=���J��U���')1��"���&m��=��omܔ�ƝSsP~�I��K�~G0m&A�b!�Ѭ���ݡ��h"��0~��
ہ$�@���w0
p��N��R����m�0_g���(<M�B"���J!��5�YQW��қ� �l0SN�$f�s��%�M��Ճ�ɡz�rK��~
�:�}�E�l��5��N5�0TQz��nnG$e.�B�/tҺ�����[a��5j��f�����^MT��<Tl���X�5.�H���z��&�@GD��m���>��j,�{
�1��H�	q) ����:�7Pڳ����$�@8^�tv��>���`�:E���V���L1��R2[��M/�w�T���x>X�ߵ%C���J��Yn���h���!�8A��aڟ�%�e��Q9@u*väNo��E� �}<�l�ӫ�L�P��o1& v0�QaE�n��	�O�a�HyT�Rf���*a�}�t�A螒�k#���A��~K�wk�6���y�� ��c���5h�v��	��W,;z����NFt���#"g,"��8�u���OF�`|����v��y2�%�1��b>tVWR©��a�,���Td��騵Kۨ�"˟�ÇH��Z�S[K��R`�:�(�iGM,<pe9�t�|(��e�]q�8$�n�u���}�vx �����1����ƥ!N����I
I�%�x�DyUA'�E�D��ȯ��t�N���C����@��%���<���i�vi6O(�����1�0�m��Rm�YdV�X���h愰�a�5]�;�U��<�{����z&>�X�D�Me͹n'^^����h�7�IλH��bS�a>�i�I�`Ld�����D�LAuv��D-[ Y�&��v���I�]ㄓ4��ϓ���ͩ"n7;��<Z���vb��N���C���K�M����ϭ�o�V6�*�$AY�~~��*�S�ȗ?#�u;��E�o߀)��m��2��p���WTX�h�7D��<��!*At��>*��2�+g@%0���%Zp�Y'�,������A�"���s�I��E�`&%$��\�7��߳�Рj�T�˘��&���S4�����E�t�YW
e?��:ڱ��#����d�(� �`�6�����7�!f� X�*����g����Oג$�f[;��|��i�n�v�ߪd�+:��L��`���%Vp�C�i�(�q
Za�j��9Hf��U�2��Xa6�f!᷺��Qh�KÒ@���:J$������!�4S���Z�������p�E��2��6dA&�2�5�@�H"1,W)
�����6�)�'����W���~�f4��u3i)M��d�K�y>�oG	>y�(�����T�u���A;�J�^fi��B�W��#TI@�	�����<j��a
R_e�4/\>ú�kl��@��� ��I���|��-�{b��9/ʆ>�"���w�B�����>��×T�A��X1��	�������i[��#��6��U�>s��ÿc�)]�a~�&I�X!;���#��K����o���l���q1-'��ix��2�	kAu?��vF�H���k�����5NWm�uJU�V���4I�eS"���#ُ�
�`.�b�)���0�8��vyY!|p����f�Ù	����$���E�p�����o8ڱ3�EW3�ä�}��fM��iI�/s^�gD��]3��/�6�)WMK��'j��F32�]Q�����K5����A��d5o7/�φ|m��¸��(�oGMJ���*�;�U=�����r6'ڸ��4�k�V�4�,��/[�G:����q�
��'���^+V�Hџ$�C�4�������������ւ��D����l��&�]�>�"_r���N,dqa[�UX���ۇ�{˷!W3 �J� 		��gtԁ0GNм^ƸS��2�ݣI$��te)W+�bj��I+j"oA�+�є狓v�ޘ��\��e7{�U�2�ZP3������UmҾu�K�w�R
N���j_�Z�.U&��]2$�L�xiP�#�i`�i��&�ZMj��{e�����=���-[{�j��;�`C}EM��N�-h������rUKQ���@@��΃`rç��ҝ�p�F�nk���}ߊ)��,�i���O�`f���$r���]+r�e�5���l Y����eλ�@a
벀,٠:84n}%�M3)�ru�]�2D[\�ب����CFq�'�4�KgVz�.-��#��Y�N<j?�{��z3�rVٸA[tp����!���R�5������4J��#��7�H�D��E�B(�vu�V)	@��a���rz�����AqΎ�n�`/��l�'�(�&ɧ�&�B/�!�:�7V$*.� ʟ=B����e�S��EW��L/�+\��������֝0w8<s�n��a3.��4��f��?�M
����?k�}��}!@�4&zk-|j+�et���^̲)��q g?a��|M�kD�������٥M�	@��3v��%b��b���0���*=�W�-��7$�M����W��0�T���,,�ذ��N~
u�U�g�*�6�+	Z5�r�j�b�"��k"<��p����ib�7N�p�&���ᲅ�ҋ=�&#,(n=Q�.��b�k��x��*v�O]F��X�G�a%2Ȣ���tБ�Ӹ�EÍ���67(�>� �^#Q-Я9�1�˖4��D�糰�>�H*��#�q=`9Q��,�/�}֭r�s}	��z/j������s�6��hu��S�J蠚������2�0)繗�H����5�2�	T�#dj �˼DH7�� G �%\^��]=AmJ�fo"�+��a�hN?�V���f�p��C�>l(��q�8��v3����(X';e�M���~�57�Y@��s��x-��ڂ��'p]R9��j�/i�X�S*b��H����YC��0��F�t=^�_P�X�Ӵނ��L{��)�c��T���R(��!hn����3��Y��_c�s�փ�䷡�� <]�mF¹�w�i���L�Q���� ���e`h�ҭ)��[�����L4E��E Ν7�`��z�4K�0�#�u!���2j�,��Q�=ҍ���؜C{�8�����Uŷ�~�?h4]�O�9�d��j�z瓲o�������xj��3G�¹Dj����T�V��U��[�˰�)G�4C��P-]��P���+��RƸ��6�!
�꫗�\�Ȑ�\��t����I�����{iv?�]�Lz:�Q��z�e0M������5	=��ࡓ����1��6Y� ǎ}�_�VT��S���$g���hN;m�z�s�G�D�9�$B�7��8[�1�(�e���33t˄��w�cK��61g�$��޶-�:��a�9ܞkw�L�]���C�E�8ę^���Q����0��5u;�e7�nR|RZ��������a��C�I�̀$��1(�N~�(N��a�r߽�q���Θ�]�մ��Lk�;�[����r J�ϔ�P�e�Jh�^��x�oԸ�_!�	�j�6#��J ��I�$8�DaNl�`�/	򗙉ʱb��T���N<�g�KC�.9C�k �0{��/���023�1a��ϵ����]ܿ��U��J�F��|)�/����De�a4@�6r��c�E�S���c椢�V��|;C��M(v k�C����B�h��E�Ag�IU[�� "�G?]k�aZ�����(.bw�^��Q��X%z�K���,y���=���/���k�`f�f/�B�bM
��K7ְ�i/dy̰�i+ܡ�#*��XUo'q�Q��� N;E)��~8<H��N��S͘S��/}Wܶ�����x�|�v�G)!��V�P�_�l���	rSd��6t���@",�EU}���R��ӟX��_$�b̀7���)	E��6��
h���!W�QgG#��{=���ƌ�ï�32V��e�����$s��n���:�\OI���E�A.2W��֕�HmT?Yg�*]EBTgn'+h",x\B'ߒ!�}  mo�����v �D����1B���k�}��.����7� P04ޏZ)%�V=awA�l��{1�J�%氘`.��_�e|s��Z������}�����T�C�&�9�� r>���^c�,�$����P2\��4��_��r���m+A٨&���|��)�jw*�80"�"�}UH�ލ_\�7իdjȤc��K	��Q���2�F o��j���]��Cax#iW���J��{��B��zO���Ҷqr�j�@[�y�s1�F>,�@/�_5���n��;���:
����v��
�xJ6F�L1��7s;R��X�Vz�&BgR]ȭ��^�%��<8�ݎ���"�"�2/� rϡ��?���6w��KX��]��42NL}��,���5_qza�,b�BzH���1�-PE�@G/��*�
�~/�������h:j`�iŀ�{�a�c1�Y�F���$+��g�]���+�*ށ�t��#�����L^'��e�Q:� -(0ar�#U�s�O �v/M����c�!�=��J�,r�/k���	��m?l�zN�1;�	v�>ē�ϮҨ�t��%R�!ͦ>�^:��$��LX��(w��C  �9,(��F�R1��W��c->ݥ0zi�5<�Z/�>U)�.E9�$c�90��-��gķ�e��>x���>Ms��E&�ؚL/#��Ie{�9l"����S�?T���3�������[�%Y�^�����7q�j4���MU���{�w�}q�&]�t�1�m�mp:�,�T|�O�u9�K��SS�V����Fv��1��-�3�j+7��&��aD;{ ���
��ȝI�Λ�)�J�dY���ҧ�|Ů�'�T�wg�4�
�=D�E�FmG���=�T���8LY�&ӿ���O�,SƇ�;�B3�����8t�����e���L�aE��l�\�@>�>�X���S���B;�f�׀�g�/�F�{�f�"q��yz�q�AEd`m(!#�]X��G�(	�-T���\�S>~o�۳��6��Ozm�1<�|0�Gf�_q
�n��%1"%i��b�t޹��w�7 V�)t[Z>K�A�ӏ~�T�+BV
�����W|�e'���H�"|E��N���ݿZc�U��0����#e<���௬ҏr�gwbj��0=�i��b�j���-�B�C%��C*�W+Ɉ�m���ԊH��S�a��R��N�j_p�����#��m�^�7�����r�~�1?���Γ�C[���]�o���?d �Jj��O��4����������=���e�$4�-�(�l��dY�
m�`����b�R����<��B.@Ax���t=�0.���y����66wS��h��hZh=.�/���H֥Q�#A6��zyx2�4D1�dk�>���k�T�r��h���ψ5)�b���a^��s3�G)a��������(/-zVu�������LŐ��
u$�7�n,Jm�}�G�u���'��Ȉβ�������p���x[��jw�M�0�s,��3�u$��b}2�?�b�F��/,n�ۦ�}T�2q����ߗ+{����o�wKm�SfH�
W�^���/�A��ݡ>���kz�8�M�֬}'�(E�"�i��v>���ޝ+=�cu~�:�<e�ƻ]��]V���PL%�""<w���eq�F>Š�mN�#�s��Ƶ2���%�=���$x�%�s'i�RM�<��щ��"�fw ����?������40��i��F�I+l��<�ϵ�$lWv\):ҍ�I���S�{�q:��I��'��S���LB�!�<1l[<��s|'�ı#�0�.�]��g�.������
B�R(�D���VP���*��,r_ `*rld���u�/� D�f$'�$�_G��"�m�5��	����34
~Vx��{�dY���?��<�F����Æu�?��B�> TrX��'��2�4w�p���iӼo_Y2��3�w��ǃ|8�8�^|�����)��̊��&[����K��LS^���&TI���)��d���G�7���`�OX���M�6ً��I.7ӄ���a�^�;0�BL���ɸ�=[��g**1{����W��j`˧O��~G2�YR{�ԭ@BR�,�Ǵ�:��ʃ�5@p�� ��eͅ���/�����r-�w2�����0��"����g'	�+
ke%��O�hBD�Y�ΟY�#�;h�XX��t�����;���|V�ӪP�m0ׅ�`0��;��Rv�QB�?1E�>z��͘<\���fQ��Ǫp�#���3�tH��qaY�)��ɵ>�c]-ό/�0E�3RZ�"�ԙ��_�7��M���,h7�ұī>���uCvs��5C���	�_m\�� �7�����j�t�����!��P};
�39N����L���!�c0��	��c�y� �)A����fC"Ո��Q���m�>�8���L8�ߏMf�����#��;-���$��2Y$&�(�Хʕ�]�(:
~�#Q޽V@� Ya���o�j��k�M)�l��}0磇�z�$0; ��
^i+��(����O搰� Z1A�Dp����^�tQ��OD]r�� ���;���8 �@g�6	�V칺�|?^~��s{�574Ӆ��%�PK�'4���g��_�-�6�1�ǈ���ܜ��O�M�,��8\�U��ౙ�)�0��$�Q�$��=�=��8޿�ƫ�e�1�F-����;�v��<�f�1�&ca'�`�y��ह��Ƕ�0�o�a�V��(S�ۍ���PT��&�f�d�V:�>P��"����u�^T���ʇi`���)��	xQ?�خ�֍d����/c~��n�\��r�V�њy��G��y���������5u��[�¡m|;��*Ш�:V��(7���4r�4��B�� *B�C���X����s ኺ���e�H�?�h�<6���Yò��/���	r��q.p LԽ�H��.���Z�N՛h�G�..]��1[$�q��- �i��U������N��W�t�J��+?�eu��Ǳ�#���-�9ޘc;)bS�6�şם
���(C�q��
�I���X�~r��	y�]@?�Ί����w5�������V��=�+(,�?���n��lɠ�9�K��띝[��
�}rSRK�N�wJX���ga,Th����Zd(��D�����, b+����������K��${_h��w���h�?bKЋ0ʛz�6�y�nV�ߜl����$�'UnQW��1W�H�D򍾏յ��E�����ƘɌ�Q�9ФY������nQ�J����/��^�A���Y@��m&�\xP-㙁�j����WE�P~����
�b�ݯKA�ǂ+�g��G>x�2O��^[��@A��a�}�%el9g�G�tp��>��/2�����_���P$�UsUsisk��Qs�v���0�|�Ω>d��y�y֘Xd�C9��0��C�RfZhE_��̝���.� ^W0��qU���Q�B���`C�8���nz�)A��..E��[w�M������X�Q�Y07=�b
10v0'm]��u~1.q����XV>A&�jk`e�o���J������m=DH����V~�6CW�fP��(f�`�@�^: #;=똀J��S���e�vmO��w��Ad�6 ��.� �K�����޳;�[����y/��7��t�M�����ө��F�����N{& ��{�S�8�{��"��&�����Wڟ��<�b�.+����h]�.2�N~�Z����G���>� ���c%_��*J,�o��F6Rt�)d���\)[ |l�����%���;��v*�L5���5��Dݵ��PO��h��
B҇�s5�됻�Փz8���n�졗:�-�~��uԶڗ�g�G:ů��,�w��a��,M��z���Z�3����� H�:`�e��"�ݢZ,{VXs��:�|�03t$}�'Հb��oUE�8I�0�@Q]�8�+��}H�p�)����Ի���b�{��ϻ,"d3QlӴ�>5���ܮ%��"	���)�^��QO���:J����dZ������\���cK$o~�?��Z
�I,�d �X5"��0���#�����	>J��[#Q���q�`��Eq;�R^��.\�/�mD/
>fʢĦ_�Z{��bc�1m��_z����쑡CJ~��J;H�|A�'���@7�Or��!�4ɳcE�P(�Z��!]m7TB����e���Q�|�!]�6P�:5�Kb�/>^��WS���0҇]5pvՇ�K����`E}˽�)�{0���<�/�g#@�^9�|���t3�'�?7���\�/�c�j�pj�E�R��?�ݬ<+�`�r{k�\�=�6RB�oo5�vP�s��H�H7T�1+P�����2�K�#�������T
�����ǟ=0�<��ry����#�m-�d&"â�C��M�?П�&�y^Υ��}R	��):hQ�X�9y�ь��B�-:JW��L.Uu��(���φl>l�<�I�奨�ts����&��HEeD)����y�kg� �oyX�wŅ��)��
.��;,1X+�!�TlD�0�Ɏ(�!��@���7Й��*����	&�y4}�!̅Cϖ!dN:J���Z4�Z*��M��4�/l���(��V��#��Y�&@#��ܺ,69(�.F�@�f�k���I/��K�<mlN�t�>�\t�o�8>�2�/-`��RM����}m��a�PR���� $��
�u�X�4 o�1[��t�x����Gw���*�%�:iK�S��9���l����e���9p.��<�S�v6yƅ�|i�^?ܽP�x�����h�$:���}�0'WLhV������~��Ф (Sm)���1��F�(���_�E�H��,��崸"C�k�M���o�4���D�1d�n�j�I�:��#�I��~Y��L��5�y�a��K!û@j䄻�w;N�g\h?�[�nߒ}�Q\o]
��h̸���	�􀦡�԰u,�G�g��;�nxO��痂�a��g����\]�G��D������ǋ�!����>b1������������?C�(J���gbe����l����ܲ<,��Alb5���vn��Kt(˗��*K-ݺ��_�F]�7UR3<�gO�fq�m9��6/U[��nY�y�&��)|�ӿ�zY-�?�x[��+0G��M��9Lb2r<2R�-oF����dT���̑�\!r՚���[��������腞�~��t����cd!'m ��� ;�F������ӘXN���*q�ӧ����I���Bh嫌47]����`�V�~8��!��R�;�h����gkh�R�lS�'}�`����I0-���7u~	��6�G�$nAĽ{�J�s4� ��%�.�,ICt`��ˋ�^L>_j���5y�!�y������y"����#�'�� �"���B��M;Rc�P�ji�ھa�5*��O��G��|�.P!�F~M�����v^���l��Hu��{ɕ������̮�<�/X����I�z��!�$�3�8��~��ګ���D��%8�����la��O�Z�05��4���?��|��46�U*K��h�$�(�]kx�Ř�hG�E}���XS��c�S^3&�Y�&ߡ��dʟ\gd�����;��S����5N�t�j���2E�ن��#^v1���_/�A�k�����蚖#\l�\X�N͕:�� ��	�ԥw��;&�ل��Q�c�5Sn����(T���@²�{�)�}r-_�+y��־�o +�����5���<5`	�_������L�3�����]X�ف�<�f�-a��ZH{�
�=H�kQP[�������IQi�"�J�1Փ�J���[��Ї�ք��4���c�"�v�P�G�K��������rOYY����mIn^�9��)�"q_�~�{mI���k(c���t����db�UR6�Dmm��%$�vJ����U�ӷsG��Y\�K�SQ��-?�|��%�G�@�7��+H��c��ʣ���.�����*���
�����?�Vř��p�2a6��Z13��e���KZ��ȡ�h�}c���[?e}�x����&��C�m ��:?��zs B�������V�D�>�B��#�B.\����˺����r�%7�e�%�$�c@�_�Ժ�v-�W��@|����Q��>��!#���Gb��L�p��\K.�V^��r��,���T|ֻ�d�/>�D$�^�B� O��#�K���nl��w��bo��?�1ʻK7��t�����u�Wq4iģWY� 9�d}���S�(ox,�<�c��[y��&�E���A,��Ód%��
�ܖv!ƾ��v(b8jrR��=�"���D[j���C"�;agt���@Y��|&�ϟG��*H�Z��� r���DHv��O�^.��NLi�!�L�k裈\�.Ř����^���%�$�P�Z��v|�O�;��S�T�@2S��#��t[�6�!k�� x�����xE/.�r�2/�<y�f-���@B��؃����5\}݋��>|���>�W5�Җ�u������z�����/ɵ�\�z/̚��2��+P<]��W�<�o��U(q�+w��gfcO���pz`�ׯ�8����>ߚ��<��V�\�Ġ$�e������)�([N�J�~j�;��/�q�2����<O6*�1��3���/���<g� Kc���#���d�LB�ݴ���0����9�*�{�U��L�)�x�+.��)$I�X���d�j�{Cb�� ?Ńc��6���m��G7t��_�H��.�)�`�v[ms�-���|�PM�{{^.����/)��9�AW���81��XAk��+�M��c�5a���Gj^�6�e��;�#���$���Qd�(*��ks�1��i�!%�M������7���"���ʙ{�d�1��h��^����Nn>�A��i���w�F�`ڞ���q���ʮ��Ƿ�⁯�W<~�6�?a7<�gqki�O=3�	a��E,[8�56��"�Ԓ�{���W��S�	�P�7||�(���z�v�M�TtZCm|Rh*�7?#����EW�ܷVǇ:��������W�h�������mE�^]e}nK܎�r�����N^a'1M�?�|tى�bu=��A{��f�e�Ǒ�=��f:���~%4�nh��O7�o�(�[q1(Q	_��|H��Ӥ�7�P����q�<#��Y.���kx�@�鬕���A��'&�h�K���aZ�"\8%��~vmNv�x�S����?:=������?\N��m�a������Q��4q�.��Y4m���>�?,|Y_��%��!�e긡S�1�2G�QN����:Kq��9��aPf��==����a����e�Ӡ6#^
��'Fp�cw ]�l�.{5�U�k�i���a7%�+	i���Ju[<��d�nEVR���\���t�����O��*��2��Ϥ�8	[�*�TsV��6PB�٥F,h�xs��ژӲ��]_����F�3V#���+��鿫�;@E�V�Y5�0Q^�pUON��D��vF��q���9���}쾜L���7���f�EB$Z� �Y|@�݂8f����^���o3;���@�*e�����C�Y�2 7cNI�=w��5-��K�܋nH�70��)�gD��(M�[���B������c�+~qObPa�߯�k�3������ä�)�¾.�zZ��N������:�D�ۻM8�W��-S
�����؁��µ1^���x�<GX�4�)ᕯ���Rp�?�K����vxs��}/#��8y��}����AF����ex���Rm���cÓ0S� �W���`-��Fz�R�\������LMF��ni)��V���z��v��=u`d�𯰉�~]:D�K
 ۛ��}'�<�}*� ##���c�*�~0�R�A�bO���<I��ϧ�U�ry;w%T_2�C�)<�5��9����q5�D�(q���Ͱa({6��n�c�����.���y��c�ZP�N�D���F���&�)���se���"Q&�kؐa��̝�:�@�;���I���I8��(���3�DP{U�#m멍�X��1W�!�$�i$}_p,;���BKM�y��V�Jc&Utz�rc	����n�`<[I������5�����8���J�<.뫣4�������d3=a������q��8�x���uR͸�"l���%��C%�髸���P�D��/�}��'P�Y�4�HA>ãaԠx��y��|�
���NHٴB�\8~��\�aW��^�J�U1�(�Υ�/��il�4@<g�0�Zʵ��T��o�=Lw�y�`����v�fR��&tl$���}5k,&p]���w�*taN��	F\E��r�ލ���V-I�*�Rf�,c>�M;������]	���a�Yy�*���Ofw�$X |�7�8m<�"�	,zRl������3/S�������fp���y5�de�����yQ��'��A����D���X�S������-ښZG���ΰ�/F	h�L�K�n�螒�"�a�9�4n�B�-}hI��q78-���.��:8�
_¾Y޳ɮ�L�1��o�K1L=z��A��Aa?>/T�E,���m��y��形���=[$ǫ�g�T�l�<��G���2��V{�h���K����|���h-뗕J��KgC�ᜍ4���F�p�+b BO���Z��7�t�-R�����M���&{�rC�`�H,���<��곔��)h&CO݊8���nr��-�qص
������{�~�i!�#��gDA*5ٸL�a�$��\Oį���ϦF={������V�܏\�ֈu��}�?�Z�y�Zȓ�h��*�� �)1�:�'�TX�	U�T��Z8�U�I��l���3���#�_�0����x㌞ n�\"T��]iW�Μ�\C9s�{�{Y����K����&���l�$Ӟ*XJagA`�佔�����+�8'�$�N�}�K_w�J���u��.=�L�3��a����s�.!�������dX�y�h��5��h�	�#�Z��d�d��*�d��q ��Ć��ɁL�llθx�V����^&���:�*z�ŭ���G�_㗮Nw�0D���JJxk_��9j���=X3�����{��?g�<WM�:?�c���M��O�^"��4b���ʠbo�?�q_�|$^����$�/��)���w��5e� b�,* EΛ��Ciq���j�_\�!�J
��Tr�t��"�FLփ!Ǝ�p�1�,��1�@�6ba1�٠�����ǨR#�~o��f�.�bQ�gC\�ӫƎv)ǐ"i�A-�D��>��P�NE�������ʠ���2au�c�+6wu��ūLkQ]�m���*��G����T�VrV"A�����`-҈	��RhJ��o�LՋ��)��5=w�I���[�ZDt� ��ލ#�iN]�tMhF�����r���PpqK3$Ϻ�`�@�O�M���k���CU��V�rM#��SH�JØ!�ZhKqE�V��Q˛=!)R�&�&`I))wU.���BˌM=��	�憆a��'���W����zn���ain� ,|�;&m��[0zdb�$�A3�3A%95UcڌH�XqLd�
���-l��؛J:��S�ó��[!�P���Z���5�*�>~�)�y,,[�BQ�o�Li;a��d9��]}�_�F����ƃ�W	1ێ�'�����$mF��nxS�	;&^�	�So�َId��D��mjP`2�G�;w��c��*��4�|����X	U�r�k���� ��h�������K�����z��xpI�"�ST2"A��;�A��O��ҽ&5�h�9RFHIA�y�j�xVQbVP���"b�v��~n���
T���fȖ%�\zYޮ�L�y�f���jz���P��ʹ8�Q\�.P��gP�D/b`�@�#)lMS��m������dƊ�c	�����K�f�
tuw�OMZ~�cv,�}|�l]}��b�� g軂���[�M`J�!��x��"��h1D���Kf�1a��F��Pض�V��o������]G��Q :�Țq0p�F�p z����h��z��+��&�Ү�(�))PɮZ>w�������S��ަ	�䅢����P��[ :S�)���#
��}|�k΢M�+�1�?s�����7�%ꐯ�K�Yq�h$ʑ�-�D©� EN�?=���.���~�=��V��
�=��ke��Ntڍ
E0r�Ӳd��{��>pSeA�m#9�}\�D����&jLU?�*���BM��Y��V0��b�>���%x`w��STP{a�gk1_`�m~ ��ۂ��@Av h�Ө �e�����IP���$/?��1��E(��[�̵!g��[�O����՝m��
������n��͒��EZ�J�����}]VHT�N�[�nRaFTd�$�p,���^����T<ݵAm{8�]#9�u�4X���~��C�Q��~��ٰp�.����;��c�m _��}f[�1���V��x�9�'�n�㑩y����y�t�S�8�pX���=]�<�N��b�+����V���dV��5�6�d�RZ��@2���2<�3'A#,V#C읶��6%&�h⤇"S�͖̎t hd��%h�������\P��R�GBe, �.���~�X%gNPn9��@���Ǹ۷�5{��!�H>�R&�T8���s\�����2��,��#�����6�r�hRJ��< 樳��)�jo|=�f�?X��T�ս�#D��/�X {ix@ܲb8�p�d���8����*�|:��������̜S�Q�
�D��Ħ��[ۮv]f\��j���HD��b�2�O�΅���Suo�(?�Uq����6��8	ɱ�]�H��B��
-$����;��ָ���C*�j�H�1�hw��r5ۃ�r�]��	nq�!E7X}��.Ʒ����n��w'�E!��v�>x�Ҕ�(䋍���lX���T,{XG[�PZ��u��틩��q�Ul�{���釖aq,��)���1L�zH⃉B�_=��=?��~?t:	r���9��ڮܫ��:y�S��d��2|	����s��{�O�m;.^� ���C��,�S��j׎����~Γ�H&K�7��&�����o��~G7������Ȳܹ�@�c;�+V�m����1�w�Jc8�����,bb��EDks#�<4ln|m�88��>P��e�rF��7�Ɉ��K�{�쒍	����fÒHUl�I��]hVT���
�b�!;.�
�ZS�ID���!�fơ��/�ht9��?� 0L�h&d�A��ݫ,#}u�$�r`F��������cv����J#z���rb_U���F�%�W`�-�I�B���PΏY,��-�S�3� ����>�P_�>#7"��<��܈���\D"�rG�*,J�����A�E��E������ ����|�ϊ��̔�8U.�/��3�bճD"g�ȼ�D*�}/9Գ�R��N;K5�켵�����<Q�Q{�""�Pʦ%�N�����f�@���fۀZ[`LR|ބ-Jz,a B�u��1W�ǡK��!+�G������|0�3��5��UV�-pJ�|��%�/ �@
�����n���r񢔺����{�$�!��Ja��9"q�S��HU��X(�~:��	�e?	FC�8�
�O"�,�p����UP���3f�ГI]�b��켇u=�9��A$#.��ޟty_�[�oY�Xz߅[�h{w����TІ3��у@U���ʦ7���hA�x	Ãs~zHĔ��L����L��i[���]fR[�(U�5d@3Y�$��qB�j}�&i�N�$��5��a"���`��r5Q,]m�WҮI�t��G�{AQ�g�^��læ��'����wk��I��R{4��&�S5�f�Q�T���Ԗm�*A0��I����{ҠP����:tg�`��YZ���?�2�k*֚l��_ܧ� ��ŕ���z�5��S��A�JzM�IP=Ũ#zu,�K�;��u�?O�U�����q���&�Q�����u3�.��69���St��B
iJ�P�x���[t·@	�DHd�h�z�N.'%�
fi	��D9��
��������--t.:E%w�:����'d�>>�Y�w)*����
�Δ�C��M�H0��Y.)[�.c��9�Q��\��/U��2�i3�����)J�ؑ�g��Β�}�)��EX��p�'Q(39�0�����Y�6�-9F,�k���)��܇�T�� j�;��	�>I���[�) ��F����^Q��	�[��6�5BN��A*\���9�u��W��d��E�)BL�ZL0��Y>TN��ے�N �p�����&�l�����
$�R��zz������/�C��xd�e�vC0ϯ�r�>��"%F-/y�dC�� ����xD�g뎓�J���e�M�a����+q�	>~��C�h�v	�]/杲,�f��y��'�%�6����)"Λ�.��.D����؆�����@$[�a9�"�sf�IY��Ym����{�XB�㬯��S5܊c���X�0	3�7Oix�d�h�%$��S���7=�]Y���C�f�vy���\�̠&�zR�.Q[�=3�4�f�$�G{�penp�3<u����i�j;�u�1z1G*�� �I�������K>���@b����'�l�������Q�e"�voS��gs���S�}�4=�}U�'�>�fM;�j���(䲢$�Ɯ��ſw)ӛ-ʤDJkv@`���a�N,i��Jf�4��}��_kum����a7*��d�,�S�T��m�Z�{�(�!f��tu{��(�?<����9Nw���Xt��1䝘��R���b�NR��Q�Z¬1���q+f�+�^y�\��c1�ב����>�ZM��h�;{p��z%��BV!?'>W��bjaX��uWK�02�I�=�K�i�ץ�,�&�qw�a�b�����'���S�*,%��a�� :�;�@���ez���d��)�U��fR&E��}�_�.k��@}I�j����^�6�cH���k���Ë����`}����q[� �Mw�}US*.����?��8���,��=4L�9�]B�6`c�~	:��Ṟ*7.-ˬw���h'���3̺*�z�D���F���pҋI�=��4���4�v!��ͰM�S�%�=���y9C^�%��o�K�9O��L"$@8u��t�C!9�:Ǟ��vSoS1�,syʎ������J� �]��c�Y>�i=:4dl7�:ϩv:��z�}_��b����t
?I��%�����BԄ}�9�慿��~v�����YHr�w��ґn�9��pqvN�����T�l77:�����S��u�r��:��:�i=`D��5H��!�_	������?������Ld �;�����"��?,�t������p�U��9�ZD�
�������z��"�@bd}팎bf�}1�\S7�`g���A6]"���Rf;uçO���H��ՠf[Elʽ�yke�d-�9{��'R*���@�Yj�)�sT\I�
4��ę���Ԍ�D���74�/��	�5������챹��v%� �@Ӳ���a�y���b6��|j�0�l�Q98�?��
I3��������@���K�h��N�[b9�4��J1��-N��qQ����!�f6�.�t~c������Z��S�X���D0�ֲ�h����&*C���l���&l+y�,���_ �4�iےL<���H�^M�*D��c �E�Y�"��QK$�XӲ{�ܢ�/���� �	�"u�S�dF�͎z���o�Váh����OS���S�v2~ߓ�D���4Q-��`J��ew5'X�zီXh����ԶO0=�?I�5��f�6b��)�s/���;*��FB�Զ^����	K?�*�}d�@	���K.0EB�ɵɛ`���W��\yI��V1�ej>̹�������Vm+���8��r�}������j�T�/�Yx7�_�T�m��:���EL��h��\������A>�B?����h4"��/e���H�w0�n�� m9�7B�謡W#��rU&[���ψ~q9�MS��~5�bO�r��$Qq�1�R#ھ(+�}�a�~���u�f_Z��c�NI����9]��w N�6� %QUV7�$ޫ������S�(W�z}�-��n�s��߽�LD�R��
	v+�w׮��7�<F�c�R�"��_��i��d�V߄��\(��*�kʯ�s�Ύ�L$�@��j�ֈ�8����y��ԗ>��T����1��m�h,��԰��l�s�������H-O"��}Y�<"�{�_�Ht��	K8��Qc���\�+V�ߠ/&����'�G��$���VDQUUgoX䒁��������&xYP���,kͱF���|"��jGaTd�!N͕�eN2�o������Π�J\�j�J~���]��a�*�ǰֿU-ʟ`V�7�s��"�N5�������b�W���TA��Y��K��}�bl���mfl~�p��v�j�z�.S;��A�|=d�(@2eO����.�h+���:��u�v~�Z�H���˿���Թ�f�����(���je��{ڡG;َ���Y�a��~QH1����6D���γ�%���3gDF& �,r������]'��uDT�������ao&p	���@��eq8�A7�	�����/3M�/����ı*�1�B���-��M���c�QQÙ����j�������&'�G�XB�N���M�|s$��mon�3ʋsA�R�ͨ�%�|��g��P���"��uŉb��zʡƦn@Л��x1 ��q�W����G�)V����=����6"I�m2����2�[�b���F��'�6\��S"AB�)X��Bif�k��V������N�-sK-�>o�(�)wU����{�v��5�@�:�{�o�D�uv�	 �<B10��v��3���
r�Y�/��o�㶅���j͖����ĕ����|@��A����&V��n��|2�r� ��,
��#�QM���s~���z�p��2��n@2+���CW�ޭ�%��m�]e�A3���O�$}7��}w��̍G�%���l&��n�>�P'����W����-t�A���b|)�u�Js�l�y�rPQ�^�6��� a�i�1��O�=q�y���1NJf��+�Q.8�k	�#���0^�g>.yP�F��W�찂���m��9�&(��M=ʺ�܋�k'�L�/*%��/�4�kd!��Ú�GBN��׹g����(t���ݍA%�.�[c �R���Q��湊��#tfA�c
����e��;}s���(Ѧ'�)��_�3,�t�v�G��@�E�e�s�>/t�]��YѮ��C�x&�J.f�<�Vd=d��a����=nD�	�5�m����ם��V}�wV�I[�*ò�A;���eW,��VJ��IR	���DHb�s���ȓ!ϭW�
G[�</�A��f��&R����3Gȯ�gf� �94��P��m���m�-�u�}z���$<�z�;���9HY�|&����IU�pWAV8�b���ЪIŤ#�ޭ�����N�����r����h�r�uT�;�'1]uWu� 	;͵��}A"8`�%Ri��z��5�`�n��P���?]8�e������Yݭ����f𠻿��e�4)]�C?͙f���c& �o߯����G�R���EDd�Z� ��aV)�r^ce��fԄ��Y�"�n��b!�b@�� ��.�8?�����Gb���"N6 ���,��F��=�> Q� �L��o�z`�RI�������n�{zX�c[ֹ=�u?W��:�&�"t���?���
5�2+��3P���e����i�`�4���7�� ,/�������L��װʐf�%��.���,mIFqWhܰ�ե͏���q��}�o����#�\�C>у�X��ԌW�Ѭg �09=�'���h��̓��-�~���\�IϲZWD.n�:X2魮M�Յy6?rY��u@Q'�i��F҂̡�҃�� �PM�ǘH�T2�XL�R(
sz�(�DTv�%��xவ�𴖙'�X<\��g�5�=�9�?�|�����ZQubŷ)z��bY��[e�/�lx|�f��.@ww;?���!L��وԐ@Ԇ�d9�_m7�^��=��x�K����{�@ ���~���Q ����t���8Er�2��YI��|�WcP�={�T�<�_��l3��w�E��':D(�Ĭ\r`z��ٚm� c�'�*i�5�cV�W���I���G%��0�G��m��[<h%v�{����/:�5�/�����IA�g(bW��^>��!$�R���b��V!����W�|��*�`x痮ܞ]�=V!X&��y�����YDAPcB�7=�E�����0��j㸰֓���io�6�kF0:�WCjFo*�����ߗO��E1�p�� ����kW�oH-������n�g�V,�ܫ�T�-��o�087��Ȕ�P�G��r��}�݁��s�F�1:�G���������M�2��*ݬ)7*:mL�Wh��Rl)o\+	TC��"���ϺZ�K��f�=���J)�U����|� ;O�T�b���)$�ܯ	&Yq�2�Q����F\*=LұZ�
U�I;�3S�AY��e$ތ��q!���F����楇6�Y�8BtW���~�� �-�.]M��{�������V��ՙ��Iw5�ƒ\d0���<.���V�lӲ�n�#��� ��^x/�{��G�@�}�/���L�������3l���"��zn��Й_��	RV`�2w��" ;av��vXr�
�.��O(��Ѐ� �&jV�&,	���\�?j���K�$���1�$���1�k+�z�����3���z9����ނĺ}}0�ѣ�I�5�D����ö�fz�@Z}��TVX��7�{Z�wΜ=���(Sт9S����.���5�*{���,jޘh�E�a���o�|;z8�P}�9o \<AMY�)�'��m��/a�F9H��+H'�T~��-`����jI#��Q����\"��.�ǒ>���[ #ٵQ�+Q���W�0�F$���@1k� �)�L�� p4.ɫ�6L�<�/�hvKӠ�;��}N��NFs����ut�8_!�DhcD��N.l#V�W'*�٩�fn�OɆļ�3�*C����s3�S=��W`���9�B�t�f�	%㣏�ϲFo! um�)c��H*C���x����c��h%{k\μ|��]D�l�����/���!�w',��֗�a}� ����	IH�c��)%(@���>��bq�,�0zL�/����"G�y4�^�UC����i2�5ДU���܃��-��:l�E��9�VV�n���d*�#���gMD�[�9B�/����2ʻ~S͔�m�p$�
�Ǘ��PZ��sP�kf�|��~�QҴT�����ҝ`"����l�({kYy�1ͅm�mg�.?7*��|��n�יĳX�o��y� �9j�;~�A%��3� ��ܴSl�g�U4�Z@��@��!y�MZ�8t&L��
hw�p�ޝ}�F�}��.r��T�����q8�T�p:]��5���ub�N�P]Q�X++���r�j�N_Q)jn����s٫�S��ߤƹ�&���� f9Y�f��Q���Rtۧ�c�(�$��q�iV�ìuS5g8^���}�;�
�-D��e*�F�μ�@�k�9x�Cp0P�;�2�L�B�=uc�%7R�g	�V��
�J@�[yM\-��U㌑���4�SF!]q��)���7��?�4�*���GP�Vww�&�b	d���;��:�����{�leӮZ��$@�^M��O#�]-G� �F�v+�-Q�9C&k�S���BuF4��������%���qZ3и\��!M�[�۠��b ���,�+���=D�uqPܒ�W��ٟ0�yx3+��O
5os?Z��fkz�cu]�w]_{�ߖ��� ���*�ƺ6����V_ �R��5	VI-���B���X]9����I��R@��MzP�S��c���d��h �U2g�#�&\��p�h�~'d�gc@"�&1���M�_ ���+O���UO2����;����S8(N����ڠM�<���P�L�6��(1Z׍�?�@M�&�R��,�sl*D{2�! ��f���O���ޏ�n��1�b��a�7j�(��Wk��p�i�)�����2��,6����91�6t`��]�:��k��@FH�]Q;���ƺ�����m� amnM|w/�u������Y��H���,��Q�i(B/�㊥TR���p���b��U\�b��9�ݭ��&�D��s!4��ԙ�C�͗���ݷ���M���\ d+l����5���@\�>��UC �?{�1i��f�u.ER�D_Aw�
P�s����:��,�m(��k�����n2�L�y����5�%�Ԥ�����]rS���G�6d0����$�\r\��u@�tw��J�W9D�Gl椗���{&J_���3���Jʳ-D���V#�L��pq7��ӳ3�1m۳ �~ �]�mp��EI[ŷ� 3��R��J���<���<���7�M���RF���8�Τ<�hq��y�VP�����M�:���p�)0���UW�.�W| �\ܓC��ʹ��Ԥ�&VC#W���)�u��e<�e�{+�;��%�9�%��ϊ��vq�e٬����3"K�c��ö�C=<�~nK���@dV�\+J�2y��S@�1eB轲�4��J�$�S�SZgsp��g�o	*F�L}h��Jʩ>�Z�$��#�J��f֒��L'j�#\��+v̡�@ d1WN���S�,�Dv�g�P���U
`�#)�uGM�p�^{Z^�� ���&�=�u7��U/���%�� �y�J����<�7�P�ܚ��U�Äf��K3���E����J2D�d(˲~�x��̍�,.��$�����)x�9Z~vfܜ V[Bq��Qx9e	�O�a`>bj����*@����H��\T�[�ۊtE����3�$!���ɢ��%����a����?���������A��2hk;�(��S&+�j��p{1�f|`PS�����N��"�"'��r	���f)G���*�s� ���~��%}f�D�vk|���z���(Ǝ%�v�&@����#h�5����h70� ���n&A�, q_���蟺��a
(N�-���q�ϖ]��.��<�x�L�m���Y�>��zVo�#���n�n�Q��MIC>>u_�}��3i����<� u�L�߱/��`�EЭ��ּ����Az3NC�GS�^��uĩ�zn�,���Z�q~���&�V��c�y�l}�$�����2++�TG��x�HD��6AP��<[���^BU�_�%l��|��Ms<�1���m��O��LM������7�Y~�|B���)ȑ����D3b�D ގ�t����'\4`�-9.«_�$���,�L��w#�Q�Ix\H�!�����A�C�������@����H���|H�v�=�ʂ�����F�Ԫ9��^�9�5�s�k�&�n1�C�ɂI�~V���!���pVEi�E{_K���<�t�$��y؜r���`뾾����]��w�=��:��ѓ��{"��
������c	�ŵY-W��$+FJ���-M����\���Y�]j������9��3� ��紳�ۙ�(���v&(.�f`>�0ܥ�m���ZG ���RD���3�V,$��tZ�x7�A^��#p�~��zٹz�S�:O}_��|l�2&��eL��)�Y�f�� 
���G���H�Ã�e���t��.	�����8�Z�h�g����=��QE0	��<y ��[9�8:*�]��-��e<ydҡ��	���P�BX����A3����ZC�����}?�l �� df˭;i�����@��tR��U�qܻ���^��v��ף̦�7+�7G�^�S�)c}��v�7l���~z���$�!4�=l�O�����Z�X�8���o���Nq��zC鲤
(P�[^ڞR�e�FB��;Qxv?��������1kf {���/Y o~U��A�W�£�w�81�zLb�S�6H�$?��n�ӂ,1JJ'�H��ŝ���)�Ak�q�w*ͯ�|�g[sffPs,j�#��[7�T1!�<���17���`�8U��A���{'�]( cB��T����s\z�3pK����TD}���a(�ޟj<jmId�q_@���@�,�ґa~�8���U����X��f�C*���Ғ��nܶh��fq���=h�JIU��W��+�2�/K��Jyy�o�!��?�+|�3���4MR�����M}{׸������s����J@ڣ;�i�u�;�n��oj�|҂��A��Ϸ�+*ɫJ��ˠ�C��՝��_���lD��!�Q�zx�9u��my��7y�}�r�t?���3���ZC6�k;{�g�c���#ϟ��	�'��vO,�菸?F���̕C)��M�a���д�I���$W��E�vq�
�DU�l��*f_���ԋ�~���Y�\fR�n��_-Y��G��x�Oŧ
��SG3�>�y��N�@O��y���̔!)����٤���F�_ٌ����V|d�I�"$}���3>f���Ң�/ �s�!���D�������͐���N�Okk�7K�ן��L\*ω<j�M� ����Q���T�>M��fC&N��b� ��x��/܂��C�FB�P݉�7*b�K�����}�Oݎ�s� J;��"�ݳ�xC�\x�r�U�3x2�s�NR�[U����*sǌLi���,�;�\'���^�Z�a����E�U2qq�-�����Ÿy���>`��n~H���w�V��O���+��̸/�uj�9��P>]�0	d����O��ސO�ƛc�Snl�*h�϶oQ����C`&<��Y1�G���ɝF����������F����M߻�aR+cK��U��dYN�̻�lGkiG��F����~��+F�6�P���1�XbHb���A��-?W��8$w�!s��1/�R����8>��E�z<
@�|;�Ee�:��[�G2�?��P[�F3��,@o"O�}�\�Q�ܡT<fv�Di�ZWe��:�{�q��x2�#�v���zZ�ȉ�J+�p�С��6�����6;Ȗ�U���0Nm����5�7��Ð�Âx�7�5�kj.+�t(�,�s+�2.��$�}��|wdj˾����"r�T �Ut���lwd�O)>�D����(��8����\Q��')Z)�҉d*���JM�_p0�=����98������3�!,VЅ)E�s��p��`���1�F���r�!��&��B�ʚ����vs���� a�CT@�ٴ�d��L��d�+0�t�U�(��D�jr!�������E����O�%��)�GD��lpʷg ̔7�֠הC�TH�vc��o��]-��x��ƣ%+͢
<���4��J� V�SHb�4� �ﲬ�w�B���c������Y�&����BᒦR��wB�r+�ȕjN��lQ���w~�ڢ�^t$�����Pܷ��X��pf�`��Ζ-�h���=ɍ�o��Ք�� �yi���L����OH��DL�Q2N�%�.r�e�|u����� -�D#�V���>}���h��R&5ΉaZ����������'����jVE���y�x�,�9���J��$&��,?.K�HX-��4B�N���˫-/fo�d����a4�L�)��#r5��̩�t+����V�^��'��~�VM�����}+&Z�;�~B����,�g�C��?0͡-��$Z�slc�`�Y�4�p���M;=�{� y#X�/[GL_���Q!t֬��<reLF���L���1
�� �H��.�$B��P`_��-�r�6��nr��1�
]���'^!ꥴ���f�p�ҵ��f��P 4�ԝ�תU!����D"�raP�e�BF�s����%9�kD�\�y�Rd��9ly��&�T�9t`1�����%��c��d�x�eM�'�%}sG��o�	'��V/v(����f���i;�b�_��c����@1�$��y�e�N���;G�b=�]��D�G�2?.�-"�?�$�Q�<���N��L�RdE&��Yp���o�C��s ��񳛬�{�\0�r�yi�aub�Í�������_ ����#��B�����[�"JGԪ�X�B�`��6;0	��ܖ�&��8�	a�����W;����	�%s�0�&�)�����T~���Z��Y���@���3��	��=x���42�C�A�zT�Y�I;�����	"{�M�'������f�Rf�p�+��x*�v�C�$�ҳ������߫Biۅ�s�]�$�S��+/Ȩh��¬M�n}�?_�-�!0�?�g�*Z�_Z#���Vz�[�y��#W~_�2&�'G;�(�b[���`����"���CF�Tq�׀Vx��)��e�ѝ�ڞo7f�Ѽ�P��[��mF%夨�q�T��-*6`*���[J��R	A�x4�
����Ts��2p�)�{U3<�V^��������8��D��ȧۏ?mF�a����mu�d����D���Ea;��gW3
�4���˿�G([������������~��C�֞0�4q)+J�޹���17�G��eE�C1�y�!1"�i�7�� ��,�Od��2J|�	�Tn|"��+�X���W^o����"�?�U]2������+""���V��w��]��{h��@hen��[�I)ϫ7N��ǕCF�Z��N��n���Ut1�&
CA[u:��6E�bB��s�*�]t�K�Q�h��� ��>->E	{f���s!��:�x�Z,�WP4f��>ցd�P-�
����ڼT�R���G&x6ؓ��a���rw{0��	�6�zަJelv�	 <z�E�?��zE��U��7h�=�ﰋ����Z��U��$��ԋ�Qh0IOHۚ!1�)��o2��]��c܀7t;�"���	���v��I��vA�s#���Н��3k��@�t�&�V�0��0� �g�Z���ҡ¦��n�;�O��˛��ߟ˴���aJ2�g!���r�^�C���U�<� ��J�Q��p�M$�r�9^y��*�o��2z�N��"�N���@�5voPem���=q=	��-O��P�on9��C=}U ��c�T�"�P��z��,-�k�������G�*2�. ��ބ�.v���O����
i���$M!�ڡ�ߢ#쑕y�/��ޅU��s[AC�l(��x��/4�>��wDA���=8�Q��28��W}��$��e�uR�5'p¥VQ���mF��X�Wt@�y%W4ӈ:��G0WM]�u|�M��d�HPU>�L&|����p�6�&�)|�D�}ȏ���dR�ׯ]Թ',��pܚȩ�si�7�~(ү2�p���Q�x��A��pc+1_N��us��1\!B)��	�S���.�q��Ć;�Q 8>��)�7�=�Z�Ҵj3/ќY�Ǹ/�"�.�ƂK�JRbL.����h�>#�`��)7�"�B!fe������a�;�����1X��aY����0�?pF4�S�J�F6٪�Z#�����#���|v�^����+��0|V2�m�����h� Z~Ed�DhtG^���+����1����{|^���d˗��U�_T�� �+{8_�W��1āS�-

��B�Ө�M-`��^Kj!��ic����䐩�6��>0��ڵl ��B'0O�m���y�3'��P4v�s}΂��1ݲ��.�B��I>�c�jt}ܨ�^�+�˥�A�A�#EH�zm���������u�W��� �7���a���.�IE��������]$nZ������O���$�_l�I���2�xj_P��H<V�a�P)]�� '��,'�!��x\X�G�;Q�e��SU���8�1������u����Y���:PΣ�  �Tl4�Zț�e|��i��/W���m) ��{�a�-B�ٺ�b�B�A�1�6�z{<�4�y��j�j��A�\bQ�6����#�����+�(a9�R\�kV��)�/�U�,�ϗ��0�o��iK� ���z�������a��M)��Qa��:������`������M�N#h%3�e	�>U�p]�H,��t���S���f$`>��$3�s��.���Ut��=!=��rgR1��S�I�7�z��
,܂N<�c(�լ���M�/�̈́J}Q�KȉY �.��T.����Pb�K�M��Z�K��)��~��H�`�Q˞L���x`�8��!�z|��s,F��|��X�z�9l��dZ"]�i�&m��+�����R��{6ɪ���&��KI2��²�h|C��׼����{	��1��'7�S>�S�����'[U��P���C��*�1Go!(�����9�$-�a��.T�p	���+5]: �~���ف�RoR�W��\߃�e��%���&�M�
���?ZE�-<�fx�zYK{�!u�<�
��K$@"K�b�n�"����ΕV�����]~&�J�~�⚏��u�/~���-��Û-g�W�^UɯJ�R.-��W@�Zh�7�E�`W��.��}�a1,@�V�Gp���9�I	���'���GBt=�!�X��Q�\ĉ��h���c��t�X�7���O��r�JDz���$��`�WG	�n/��wO� ��Z�Б5�ė�h%ރ��tr:���A�.�� g����&Ft;�/�v�<�-��i�빂j��j�JnA����{fg7��/��T3K�УWH)�Ѡ�.���zCb�(�Iwt�5�08��բ"t�������G��e��U�C�%�8�4��6/\C��O:����vÆ��6��D��
����a�&U�.-���_E�	��XQO��Ƚ?��d�v~n�����j+�2
��?�©>ďM�î��R+�8�]u	{��r}�2�CQ��n����7K0�>d�sψ�L�<���Pw�v��|��6�+1��L���_�5q��L�� ގ(�*qߤggc�1�~(`��+��:�#h`�@���x���}PO|��9k�� ����2iKZ�^EU< H��s�v�y�I�I��*�(��-FU��Y2xptmh�UM�
�`���Z�[����$�%=Jmf�\��_�7҃ʹ_���l$0 � �����B������P.A7
h�m�+\N@��k>�xI{��o����-����&8�𐮸��	uFڷTF�R��>�'��R,�Yl& �Ɇ
�J�J�P�	� >|_��[mM.�IP֡ij����x�â}�0�w��қ���Z
Mn�й�-`�7s%�$n�<z�0/h+I�Gk��K:�Ez(߰C}"�^��n+�ZYW���ͮ�Ѐ����mp�fi��7��q������S򖶕E;�Ȓw�QD��(|����U��Y�Qo��}:�k���v��v�e����H0D�i�����i�3s�cl*̋F��a��<	����ٰ2�ut�g��z&v3u�d��ܖi.F��cz$t��LEB��.�-��T�E��c?幙5���R葎�����I���$dxXBae�/��y�� !C!�K�9��K����E���C�������������f�`(y��\�����WR�q/Y�`�-Bw���%����'p|�	Z���>M�:'Wg�1@;��y�nq
���L:
����I/�������5YV��hz�y��
��ݯ����/[�����X��`�
���Xa�,@"�oc�==�����J�U�UC�a���1M�.�\Q��x6�af��h��G�^n���>(1r��9�	�F����;˹4�I}�0����y���F�Wd׫�{֢q����\C>�;7�5�-�3/6��$����3������{4OX���p<����8�܋��T�D�L��{
[�bn�����ܷwt���:���C��E���s��ϐ� ����Zy�.+܉T?�&�<�J)��dKo���¿3|�5��e���g�k��;Rt{�+��5c@Ӆ#���q�.Q~�h
�� )���fQb���,a����G^���m7���)ᡏ$�|�(�+�?ŗ;�7���E�~d;�q0��M��B	������k�?�<>Xy��1��1F`�.�FW�����M�� VV�Yd����½�1s5q&a"����h���lr$U�"���C�����ͳP��.Y$����2?&n� F_D��&V�V�iH �Z)K�<��,x��9)�[��.P��!���\�[{>Q�:G��k�ҽ�jS���J;�&w.���� ��]�Nd� ıٹ��� ���Q�b��)�9Y��h���szA3�o�׮��
�w�q�>�ܟơ�,f	2����*��H�^�v#��b���ƹ���~�������
����I>H��ӛ�s�خw����׺.�7;Rqh��*u�4�8����4�73 �f��9iW�ùȁen>�)�0�:8�
H���}�k�r��D����)�|�'����5��疛�Fa2����3�
�ɐ��}��8v?
�'Q"�j�79g.l�îA�ܮy%>��δ��嘖7����~<��A{�k���C�WK�V�N���h�W�_ģ��J;����[Y ���a��Erg%���<U�SU�!�W��W��E$4u��	�i�J	xP���oެ%!�;X@>l?�)�lS	R��b#���93+}�
1��x�����:�ܢ�.�!�����Rn֪�p��t2�KN�M�B�ra6N���R)�v�c����_��	
���2W/��(�[��cc�UM� ��!����/;�)��l������W�U�| T�����GL��V�&z��57�N�L�k�Y@�vP�b_0b(����P�
��_�Ȫ$��<�0^ޗ��?f��d�a��mM�l�d�7n��R��9I��u✽d${s?����!A���al/_�8�o�i]BzGgV�Z�3��VS�?
9&y����
��E�/���o(�i�]�Zk)a�*�.ʕ�i$�i�s_ ���r�H2iq�*3�}y1��e-�s�0?�rB��Q��0�D��1�ȼ�$�ﭶCϪ[б'n船�ڿ�7�u[G�2-%�.����X�raH��	�z�,ޗ�7��z�`���亘�}�<��҆�s�oD+��d��p�O8��6씏�y)���D��'������*wR%�g�}�d�?�E���V�;��w�P��c�cg:�*ki-��+�ڷ{�O6��!�G��u�������8��EZь֜~�v�d��=Ft�dG&��<%2(vQy�<#��F�ISn���W}5��X;됺Cq=ז�Ȕ��?ѯ�	"����7��-z�l�Va��Qh�Ӛ�Įv���e�
j�_��f��%˱���?���@p^��g���Jݎ�@��i��+4��	\���f�![�J�l�*7#�(�����>"A���?7��ܺ��/��o�5�#F|�1:�jq�(��+���.@¤���cc ���N.��i�}SC�Iz|�oݬC��Vdr��®�)��]�>]����|'E�U׽�hu��L�6�٭�X=�b3���&>��(4fӸ�*��V:Q5b�X��W�uZ�B�JB��Ǭ���Yhc�VbG���~L-ڤ �K�<x/E$�T�ΟY��(���xT�s@9e��}Ղ�%�I�GQ���)5H$�$-C�fr����]&>Β��e66��f�I;sR�P�C��^>5�h������rxmH�>9�jBIڞ��Z��^�割����#f��OX�Qf`��4�ٟ&
<��@��L7��/�k�w�S�x��L[�ݯ&b�~�pC�С_M!s������KWh e�Q5�ڜ��A��}/C|���es��io�:�z��)�O�m��k�&Ve��5�f�0c�3*�؞�f���J�72�hr�2���ף�et֓��iO��c��2�h[b�U����El���l��ݤ�Ο����G'n-Gzuf|]�P�~�ӂ�T�M8ܖҝd�� �,�C�(����4`��_?H-��qw�5��_���Kn���'k��iþ��N�{0�C����/�'����EI�ސ$��`Aq=3'ֲ���/R{�EV��Ή�9Y^���p3L���	Q�0��%�D�P�u�2G,��u�0�3ٳ6f��E,S�2��ǼNʠ�5>ɱ����G���<8&O��g6��^���V߾�Ƶ�֨Y����)�|�y��^�ը��s���e���;o�_���]�x��.�ĭ'E`�A"��[p�m�d"wo��C0?�B�Q��V%�#̊%���(��?r
Y
�C+���b1s���-_5)[Z}��|����=��U��,��M�3q�W�O2H�0/�Sf��W7��������7��R�,Dy�r1��z���ټ�zk�9��t�{���F��J���� �1�����u�6��,W�qϦ�ч,_����\&��(��� Yi>/C�b|�����a)|�� 4�^�a֡W�&7��ʖG�i����Ay1�P�����ٲA	����hSR9��*���l�yH ��%�z?�p��j)�T6��L�&��k!s�FQ�'����r�A�����l*u�'��B:\V�������~R��s���!��j�����e9�=xӛ�]�!�A4�����!Ǯ���A��m���%̒��:�9MI�z%����C��"��y̤�B}�9�[ T�)�������.��$�l�<�:���(g71��]�zE�����	L���C�_M�8`�5�N���
6z�aR���rn����W'����I�+#k��6���m�������pU��wTl:����~�I��tn��(�#�u���8|���[��4�NzʈT��y ��:���*�&Kf�d�.�F�Lh"$ڣ��sk���q�P�"�nB39Y���Ob�ڤٳ�Z�Y>�ʝI�kt�d⁠Zb�VP���"�����,�h�)B8F��p���H����L�y�1���νG�p�P;�p8��J�˕�P����Ǧ=q}d�+�@=���-0Y����	�&�}F�4ɣ�9>2 ��� �z�e[�e��� ���B�,Մ�v/�4Wr��mM��=^����GQ�)��"���ķ4����v��	�n�ͷ�z��HDb ��k��۬�rp]3�~��"��w�.:����v,<@g�U�����.�ꅇ���i�5IoJ-��-3��	'�L�����~XN;�:�;����ƳP���.F���!�)bڃ/��ޤ��r?�!�_��S8w���6��XHym�.����-�4���=GA����`,�նO�9���4p;H��������}−S���yz�ԓg�N� ��"���:�Z�j��L=Na�@{��d�;ߓ��������*����=ɇ�����x��Q�61(I��b��N��Q��5Ao��)J#	�t��v�����]���4e�n8��E�Ժ���W�i�Kl���˻g��a� L:GxM����}�UU��0���H���o!5�wp8�M,B��ҿw�X��?�|�*e�^��<�e�C.9��ܐ}�z'�/R"�1�#Y�.rn�&���$�e���/���,M���1��/�0���x4 ���!l	��J\��x��^�v Y1�y�{��N�걋f����-�MIA��򪼮��o�t�����Y��	NmV�]��c̻D�ܧ�1�$isG�-Y���[�Z����]W�7�ٳ�S$��;�wt|f��H�=�o]<�Z[�U��opU@��E�����$Xy3�tm\�t�4���%�����n�Ö�����Qa��皆�k��w���f�l��C�療iuI��V��0ߤTE�ޝ4pvڃրI�C�O��3Wv��=�A�W�S`s���8���Q!�����(����V�K�A�xC�|���/ 1����NV.�<_Rz�	bge�7�2x^����������,a/�oNe����O7���>Zm�}֘�%T3/�cU��d�ĸ񔎥zJ�����@�c^��U��g�~p����g��&��+�u_D�B�/F��,�Q)*7���H'��J�)@S]?�j$�!�:V�<pZ��׭9g~8��O����k��3��}0��d��h��߉��,�	Z�^���L��(Ui� C�Eqp4���ԏ�·Yz��We�H�o���=�S�R0��I<bh��w1R�˓��Q�j7 Elj�\���j>5���F��[d;殍	%~��2U�O�����yʂ�a�ێ���Yi������_��k`�ۧ0
`�*o�GB2�o������kY+�����P��Ȼ�:���XH���}_fH�kr�Ѯ�V�u���֛�?$_�E�������G �ؤg�BED��(�-nQΗ�!ғ+�ŪA�И����	�x�2�B9@X$��Q�^�F}R���B��g観ޅ�\bف*�"��F�̞������Ѽ\�d�m�9֐n��5�^�v�K��9���@����וb��ȏ�p�,��kKM�(:�L!�5+X�y�A�uf��o���p9����>�-�N����XK�%G�-��u�e�]u����Y0�Lf�Q���7K��g�԰n)Fz$\��_K�{�{8[�>6S*���OlDJ��m�9�H��
"}��3�h��ŴQ͎�;Vk�m�^� 1Z҆�saN�Dj����O	`Qt���E�9\L#g�.Ν�K�;fZ�/�F7����ӹ��`1�ی<��Ĭ�G�/��?c�jTI���k�+LqK�x�nNOq���)��Pz��hS/���E�Іt�ǚ$8�`����i%�'���Tt��t��=M*"���k ��y�g:�;>�m]t��y_���JQ��V(`�mv�SzZB�1R�;��s� �B,�V�_ƕ5!q��f��h)lPX~I��c-�ui��]J���	t��;E��&��Wd2$�
�A�~f�P,��"4������X2d���x���C�b�~O�����Tu����f�ViQ:��Ɣœc�&�h�L�l}ۧj����W:���I;�'Fn[�n��Ko&�L��y=&��hAjL�)ʶDk�\�i�Q���zV������z�� l�Ri��w�8����p�	I0`Կ��(��Ǵf$C�É�M�N����`p|C�Y���l����ݶ�ǧ���5�����ނu�L	��QW��>� ��q�J^�gL�'Y��s��f� I�:�9p�����ȎG��� ;����9��ת�!';-C�=�W�_:T�8��:eEJ>�� ��y���;x�Lb0�r5�r�6�c���ʤlj ��ǃ^4h�>ċ�T;�C��:h�MC��W'jD?ƪ� PN�V�����']�+�r.���e��ճ�2ɚ䉨�'Ɏ�m6�G%���k�?��썒��y^�=�N;n#R�l� {�/�?��N����l��Q��[��l�� >qh�jqf��3K���f�.����l[0�����?mhL��ȀE�9�mbѣu�/�R���]K����zۘ$���B��}9��ӽF�*/+g�s�^q?ܧ;G�?;/��'5�㼘��vf	�i�m��6E��j� ؗ,�a�hxy¢t�V)��<�+'r/+#�5#�X�0-.	����3�o��1��A�~�-T�x�8�xϦ�e}$�]cX0�]lr�Nk�:��+!�i\q��X���!��ڭ�?���dvk�D5d�J��/Я�YՌ�m_�ƒϫ�� 2Yd4��Y�Y�z{�PdƵB����!7����W_�yRhFAT�x�u٧C���#����3AP�>VՕ���a�!��i�o\C��$� _�����%b�Pi`;
!6��5��_U�j1y�������ͤ��-��8ƨ7���u8%���������_���#�U��iw�Th��OH��?j�}$���5�n}��V�Wze���e��S�2��5n���J_�l?�W���O�~����BmZ�����#�d����a&Ի�Vu�a(|�����w�S@O���o�| L3nC��d Ԩ�;���ЙM��SR�!E�m���F�sP
eU�d�+�{���Q[�^�Q@�`�����������cP��B�b?�7E1�� ���g�$�"��k���˒q�����u�1�W�3�(�|vбJ���K�ںרi�{Di�.��n�ɥ0�������+��*E8ʩ�r�+�'�Wq-��}mYT٘F�A(3�A���RLx�a�ۇ��ݽܙk�;fYs�b;��0�8^j����˭��5�	1�j�����|�XC�P됔�i�aߵƆ��h^T�ޜ����:����)W�0�P���ݖ������y�㾶Z��8L�P�����i%��b�p��z�^;�z�F	��λ,��ϘE�^voD��T�����U�h��֮S�гG�:]��U(m1��H�"���V�+;��nЖ%S�K����t�����.��-��ά��h4�9�vw����Z,C�7�
�*+��<Dd=�T��`(Ah~D�DV����"�{���'��;�����M��h(G�h����@'ߴQ��|fP����ʌ�I�7<G���=��ޏ���J@WZ��e�q�K_h+��)v�]�����������ʠ ��q���9cs�����.&��C@gp-������m���lֽ�*hW�O������^����N�qWu�K��B"��ݺ鸶�	���߆6<v��!���=a �/� ����N-����|{������>����M�\�J��Z��9 ڨ*�KҒYdS��(|f��f�v���,Z8�g�� ωG�h혃PM�Ҙ�>����0|�GWy��3<o�1�`.�����8�FJ��ć�5ϰ�]CTm8DK|Hy�|��;oշ҃��Y��Pɺ�j>X��IE�j��PJ$�FL���>EI����H�yF6(�|BtD��D���Zt�x��iu��Ⱥ�HL����yl��ˡ�T�`�@d2���~��|qB=pw�9��0h��]жɴ=��R� t�u�0�[�*mHC��$��yPn��<N�7�{ڤag��/e ��
/s�˟���U��%�����ȇr����[�����~�p�wI�`��<&�P{*&�{��J���A%(R�4���5����w�qkD�{�p;�y��畇�?EpEk��a����6v��T"J�nu��a�SS4�y�o+G������V�҄�ƶ��k�Z�~X6��:����XR�)��FO�A���O=w�#8d�1����ş�P:�-O8��&��Rd��]�� �S�
>-)zy�8���
���s{����x�y��Q�u0����0��QT�=N'ً@��鴈m��}6�����]�7�[W�+q�[�_�(�[0S 1�����%����դ�'
�S��,yf�eͳ���)�#�g��H*�>�`�����"~�j�\Ig�|�"���U�%�@u`!����D����FJ0`3x�Gϱ��q�=�8>�o[mѝ�q`�R<�Ms,�	�v����4�b6�a��t�ڠ�{�"^b�	�8q�A�E4�b@�)���t�dG1�hiXX�a����z
~1�DR|gQo�(����/C���y}��tܡ��}u��ߺ�mRD�j�y-2�t�+����9�?����J6���1h
�����!!�N	�p�~�!}z8���ڨ�~��Me��ZS��ǌ�E4>R�.<���D~\�Ij����m�ن�����XGz�d�C>�&␰a����8D ���R�;4q࠽L9��·)�5��}O�70\CmDx�{����$▍I�+���j�i�AQ����V�1�ywS+��,����>��T��f��0�0��j�4�4��sZ�ץs3u�Z����K#C�k�(r�FC����$WKY�+���Wq9;@��5w��2y��0��|��T����gs��I���Lvx��$��J=�X����sL�S�K�¾Y\����O���F�@�����\=J<�\��U�?�:Iưh���L +Rw��4՟b���CT#��Ӻ�%�M�~�z����P{�Rp�%VcO��>Q�r#X�y�K8��yl�v��qE#�
ȉJ(�m��xl�V�d�h�����l���Ƹ�V���R��l8O���	����{��t����/�*����5>&��d(������k��'C o1M����M����c ,�HlU�k�(��y��U�%�(�F5����b^��V<����siIg-u��)VsGV1�d?nq�Z��傸���5�+�
?�c��Lx�%t�h���:�.'�dQ�4�~{������/��xث7@�+!�T��9�P�Z4I�|��VϽw5�h���y�G� eU+"���hV��2�P��T+/��$�1O4f�Q�`�6������S�b'axsHQV�T|7��Ie��[{=I%��~�YɄ[0o�凈&���/��^���^��E{�����Z�z���u��|=�e45,W·��� ��j���5&���y����ާ���ʔ֝��ߖ��W8U�)����(	���6yzQ��������K�6��>_}�����[3�uc�Kd�?�����J�+�d�ܥ�ͫ�!�-� i�����>��z��@�`P�]�b�+2=,t�0��%�q���D��z��|"�)�` �mI�SP��l��sv���5y�=�Ep⍂6gz�'���'#<�ܧ�Q�1A`��d�QFt�G����i�|ZYO��d�X#�6^٘��}ሮ���d���ǩ�����o7<G���#�\ֶ�AI<��5*d��$f2����k>���ž����,��Ew��ڿ��8�iU/�OHX��0#��h���ҽ�- �$���.��� ��MJ4%�3M�
�>P��f��D-x@��g���������ZC�����*:�^%�&'�"��$#Bl���Hw�38�T�.`0�5D����`4�r�o�a�x�Ġ�R�R/�6���,�_�*/����?]IY/(�Mqv��N۾Y9 tn7m��7)^\�F}�hJ�}��nS�0[�&e z��âp��������g]�|�2�<����v�S�E��KP��IU��g'a��XxQJ���ۇ��(g���]���˛�]�d0N�M�6�䆖ML%���ߩ-S���25� ���&�?�yR�K�'��S4���(zb��w*$��jL������H��v��Z�i��OSd�0��|(w���K���A<s\/�kJEX������F�L@��@L�h�H����#�p&NL� �C (:Ϣp��3���sA�g�ӱf_��9�3�Q�4�fx&䭠>��(��'�n%�q�)�U@VAM�����a2 ���m�lB���,y�N!������Q��_C#A�~�&9�ve���BL�J	�p����'�:v���C�+먻���u��,�)d�=�H'˶%��A_���M���؄��3j��J�H��}$��Y���<�4�����!�Ea���O���D*����s2����!�sz�_fك>��I��б�EL8{�``n�IP�����Őj;�P�?ı�����.	g�>�� �9G@�����^4��>
GevY&sX��%/baN�}_lBl�J\)l��M���L�,��^���]<d����Mj�� ^s2U�d�p�=+V80�$G�-�śSj�vH�r����qx�T���x_��mU����)�-�,o39S
t�dT���ًdk�Z��>�1�B������W�p<T�D�*��5��vs�U�}a������~᝽����������1���~N+ ����٫��fP��|�G�/J��!�m=;�W��io"�f����g*�6�H��}��n�����7(��� {5�W1�K���E[�X�}r��I���a�x� �"�e�7W{�9J�C*茈.�_��2p�[���N�r4nٶy��lstһ^�w�s5 �.V��V��#ǩ���<�Ί�H4��nV�p20=��ޛ��?�LP�feX���d���Rz�×���]�Po٫e����b���d��e5����㮹ؾG	�%�c<XQ��V��M	�F���ک�M���3r�5�1�;HF��#��*�M~w�XEJ��9���!a|��𼘆�G�����6�3J�Jz\�D���݁(�~� �	/��$g����6��5�<S��g֚�)��4��E�����<is
�`-�?�Z�#V�B�n���ʼ�zt�H0���� 3���?e~�& ���G�#4i3��ǌ/�a.�,x�q���b��%0\��N�'�g�0	��NbNL�����hޥ�����_Ym���hѷ泳�����nT��`	L^�ڳ*���w
o�y��	��7j�,rje��y�pm-�NKoy5�g
��M�TZ�$Ajn�<Rs1�/���l�<����;,GU�PA�3gM'=���0�]E�!LG�g+_\���(�[��֜��D���蹣��g��3�*c�T'>�ܻ�i�Ӟ%<�}6@�q�YV	�g=hMв]�K�πDs�Z�8h#��-F?o)��b�&�8 ��SmX.�[��ɧ�\9ɔ(v^g����:8����T�~�(�ܕ6ީ����"�,��u�0����a}�3�3#�Ğ��!>�L ���u<��y�ۏ{��!Ñ�!���/ˇ�L2�o��
5g���qݺw�^�H�>�f#���ʉ�~R'Q��#��5��Y�M�uhk/Y��Ҵ�?�j�%��'���P�@��G� ����<��Ʉ��G���M�N3�yp�}�k�Ժ��,ЫuO�n��[�@an3�KZdx�cAۂ�m��)�#�(���/~��m���)Z�|���?L��$y_~�pyƜS#�?�"�j��c�������9�z���nʀ˸Q[�|�G|OT$FC�?n>�A#N�E���'~h�߀np���L��G���u�H���p���Y�9���������u~�������"����^�^Z�s�Y*� �nf�zVi�]�ssˬsфy��#�$8����e�YǏ�a>�D�ܶȭ��o�̶PϹg>g�;S���f��lcf�x�L���#eT�ej��o�A��4���9'I/WC(q��;��2%��OJy���?��e )tH<���6a��Dc�ߧ������o�UI���"�D',���Q�7�'ѻ�N4�<?^㴶���<��N�	�a7��?�b ��h�0�[��G@k��Y�Vi]�K���D�W��#r��?ܽu c�_K	��h~d�S����5#>���bd������n
�*3&*S���l@ ��0�jL���X�z"�{&�,�!�����J����a���9�P�v�<��z�>=P`p�mS	�=f�<�0�֚r��H=���ϙ �~���c�#
#l�ok�`���8[uEj|pԋ^�tya���`|<aY��y��H��E��S?����зkwM�`#�8T����D�۰��ӻ]JG=�D�g�0��e=΁N�Q����؜�˝3k���X̙}�TI0<��yf��B�J�Vς|�n�]�;�G��5��"3��CBM�[��n�֋B�y.��["��]g!R�*7���?�uL���O>��e2"I�ew���`d��%�w�kKW�5����T��9s0�O��;��-�Y�Xf&���5jL�9�]C��`���U����g�V�@���6)��xg?v�ӵ�F�N?�y��7�tm���(r��؆ݲ��������# �U���yQ�����,h���`ś��0y"}T~���8�#:���|�Z����5��u��/��+�.r�y'v:���/���^���ڭp^�&�?ұ�T1$xa�%-SK�l�M�Y��kN$�B������|��I��ͭ��77p�䒞{v�1��l�j2�Ȳ-ҏ�!�Du�G
�5�pC���.z���k�K?n�9�μ������N{ȧk9u��ܸ�2C�3�t��$�&�A��\��Q�g�P�z��s8�N�>�^L�)�:^�Os�\�=����o��M��L���Gb�H���Б�P�P���D^�%�����;Ъl�PTu�bm�J����}�մN�U}�ZVh|��M���p�&��G# ��2�l��̥D���r���ۍ+n�w��ͅ�ͻ�X�R1�Ac!SȽ��{W���)a|I�߱\�!�!'����D�3d�����{��3`M4�؈7<��wk�!��ɷ�P��c����yT�s�}̫�GG<�n���"�a��o\��u�����f��Z���{��c��D��"��&���K�tg#٪:���:A�W�d��\7�t���/��� D�WlWo���:��/A���tan׍�������j2X\�V/��U�mf�%郞�]q���0㩏�?-�$�k@��,����#�y��7ً~�$�qX�����&)j�ؚ� �N�C�Z����w�"�P��O&ںB=?�0=U��i�fUt�Dƾ*��f.<Vg�c�c��?���׭[t��z]�<�quH�ݿ=8;���}T� �4�U�E��������B�ޒ�A�@;�dc�t����7HM�?�Cok�xv��½��'#]��y"����p}�g&��a@ ���7hx��:�J��ʯ��C!7�2@E������L��CiZՏ���K���̴��m)��B*�N��$��4Y)��f��o����n�X1�9��7��0G~��n�8��������E'�nRWA�9O���+<;Q�DV&(�P���8'��l���p��WJ.�;\A!������9�n�a�yGD�`����~����/���Hs��_(~��I� 3�������$ �(q9e��f�!O�Ty�?FCLj̽�(L�ü�h�ݔ�C�^t�bW}�LES�W�=V%�J������PI@Y��g�G�0�t4��>��|��
�kU�;� ��J�_g_�~n���߱�Թ 	0�[ӳ��xO 2���x8)�4��ǘ�. ��2�BR莫�k���~��I�@���X:��O#��6��	I�CНэ�*�����櫥P�c���@�)������L��*����m�8~�W��
#���˳���Q@a������@q�� �;��f"��o3������m�@�A˲[���Iق�V�]��l>q㉒�#^�OP)t��9.<�>	8�l��i|RA3�Xwx���$_�9��v��\u����4���Ϛ:��;�����a(�|�bI<�θ����ΏV!����֊��U��PX	�$ }x�z���-�����'��d���y��ҟX��Q�o�I�M��v	�h�t�8��S��^mV�yյ�K!��P��^�A[��xu  ��v�o7�RV+�"��x�c�n�2ž�N7�h�|Z�ǰ����٦�N�C�x���딳��)N�$5O>��%$�2I�N�s��2��*d�gBҤ���&^�%J�d\���PCf��"䃑7�� �W�e;^/���oO4�Ѥ�}(k���Y07˱�K��y�_�Zx�J|���������ʳ2P���֏�}��՜m�i�Ǩ gX���jW�o4���Qn��
����u�����o�aKH�.g�ĖX)]�.�f	g�h����<F��{%4q�kuh5��M6��&�E
[�z@����'��H�������].e{� pi;�`�|�wd����c3ۦv�,B�{�o�M���	!��R^�/�e٤XFQP��%�Ջ�өYyH�@�hL"�3��؀gW�C�(�;��>a*c����P��,D� ��dAE�@� 4DM3�ռ��x8P�S������X��'f�j�+�id�CI
���������(��wwxɪ��'-���`�Fo^��wڀQ�� �����8�A�ν9rW� ��i-'�������A�n�#����H�O噬�D�ux����Z��Ȑw��e�Yb�w��Rࢨ�ON"-��R#���B嫎�L�:������\��1T�E�^c�$[�G0�5�W%��v�Nt�]A1�M��1��i�������L���=�AWw�/7��(��[|�/[~)T�ZY9��S�-��'��P�/�]��ڇ��P�U�NE=K�	Q7��0����AP�$����!�qI�7xrA p�	I���*�(wu�XY�B%�	
PT��F%"���`/*��ų&�q�[�\��uD^z�%�1��a+�M����6B�b���a�Փ�K���;�a��!��T�G��Dy�;0�1Sb�!�6�c�mڷ��%ǹ�\5�⣑{�2@5�xBO&��Dc�\�V�J@�?���5i�J�N�k�7?߳+�Y���Uu����A��vv#:��/���ە�(��>4&��1L��!�\V����he'�B:jv����Q3�G�'������J>%�uS�7�Eb+�]*%Z.������`��j�QGbVտʖɢN�% �:&�r�Q2���uu�v��~�����p�,�OQ�)�A�k�ծb#�Q��m������|;	�w�V��X7����'�IR�yv|/�=Bahۣ]f��] Q��Ln��u����/\�?:�sF����?J�ihrhP)d$��s�7����v���|�)�����Z�z�]���=f�V�l4G`���e��ANTo;����鈕k'�:B�K�&��Ӧ
�k�����ZCl�5;��&�NWVx|�(�H�����vU$$<>S���lOt�xO�w���ުv���w(\ԛ����P�TtMhU��ۤ�E-5�oC�Xӣ�JqI�A���(e��H7G���ʖWv.�x�c.��N�_τV%�`k%c'�f�`D�z@�&K���J��īH�S�l��\��=)�g������n�;�����X�Qrvj�a��U�2��Y-�E�I0k��ǡ��Z=�p�t�so-�����S�H��h��*S��R���eʴ�z�j-�֭�S���+�&GQ��hp#���:kS�Q6K�A����v])+ܓ��4��qQ�;�����2Oz\D�e�9�a��"������m}����:��B�o7�s��C��R���4'��>��Ƞ;#Du��O���0� �K���m�?�fA�Q؂�o�	��l��Uߊ�;l�s�,f1���P��l//�4�����Hj�0˯��fӑ�#+ɑ`��E�N��k�2.���m�˿\����u%��+��{	k�vH�#��6��Y�T��H�0����x"��[�	��p��<�S��w�'�n�k?��*"&s}8��?��?^ڌ~D�S�B�%M�[��uu�./[�����"�5��ɏ����!��$�7w+8`,:EY�_0\���<s�09|��$�:de0@������R��x԰���{����X�>־}{��mW���K��i�
y�H�PJ=�1�{�ݍ��Wq��"R���{�����7{�����Fa�r��!"^p�ː����怣NA�{��+�U?w�
���ɚ���:@Wb�-fD�����Qk˹X+I�N�Q�m�N-"��3��Dy�0�@)������wJ�{���P#3$7�O�MG"z�(,�	r�N��o�M�

�ڴB����s��1Amo��*�w�o�Z����+ j�I	N����׷c��a �3r�7�C1��jVyʗY����b_W[b�Y$wt�w����8�З���Ep}	^�u�����O<�z����iL�.�I�K>���S�f�AܤHÜ���:3� 	��Un�)U�?�.�
��ud'O����'XP�-�Q� �2����_g@�e'M�P�G��M��4yX?��c�F �$h(�<�dz}� %uR����[��7x�	�x�}[k����`:�G���7KC�
Q� �s�t;#��j�+�� �G+��߆ys����'zU������!�ߖ1U���n8}~i��kw��6���P�;k�/�Z#���a�c�0Ӻ�������`���F��e�} E��rQy�HzU< g��r�8ru.�"p�ߍ_n�Rw�ٚy��Zxw�in�L�����a�p��&9�`��C[ͫՁ�ǩo��u�	"��[;�y�v�34�ѱ����Dy�P�إ=�(x}/��kH�õ��Mn��f�5�smbf�9��ߠ��@Iz�
��8�@Y+�fT�z\9@�X�؟������Hu�P��4����K?��O��Ճ���ٹ��DGj������OKSG%�.���?^g�������4�����/3k8 +Z�������W�I�kl��1x'%��p<g3�n�$Ë�O�C�+}�����!q!��@�9Ñ#J���9���{8��)g(�L�0�~�z����m|���K��1f5XQ O��>�o�쫊Y���h�q�~�i���_���O:@4m���A�˦�u�^�f!/��.>Ix*j�=�d��.:�*�T���l�D�
7Tm����o�e������@x#vѳƧC����Җa5����Ñ�iI�\��|,�a�����&y�JxrP����K��r��SPFK��4Xd���⶞w����R��;K+w.P�0f��ʓ�Ã�.F�B'L)��ΡXˌ���~�����'�;��6P��_p��LSd$�ʡ�LS<)�\)޸#T�lH���%+s�@Y��;���Ry[�,*ՠC�*���ZJM������\$��a������b�n��X[2�L[�H~Eơ��}:���d��cwK�%�'AA��7V
!�B��B���IX�k���荥N�\#"",l
�J��m���)���gHez�S1�H(�Qj�g���ڋ�4yI���]���'��L9�6��ئ<�7�j�	��IAc�'D�ZsX1�4?yv}U���Qa��痾��A*�s��E�aGuQ]�1�QA6���ѳ�t[������|`� J�L���L�j�_Ky�����o��kn�)�
hd,esI���(Kk�(P���Y��f�,��\�f-����pz�T�O;Q���}�R��;��*�C	��
:>�F?��M�I{S#g�"��EN[K�`?<s~��}Z��X�st� �q�(]�}��}Q%��q�<�
��YUI��T��D�@�:%��E!�`�{�H�Aڲ3J(�4�Vd�hA�^�(-�cG��o���2	��[T�q��vWwӮ5y���F#��I\��.�r
R��3/�.�ĄH=5Sm��uxz�GzW�.��0�h�:X8�'����i.��u$�
���~����GߣG?	�#�FIw��[���-�89'�����~��AB��#nj�ԥ�$uw��:i5�#���A
 ��:w
��+ "h�}g�GB=C���OM���Xc2���-܉��C����ٰ�j��yZ�k�� H���諩>����ܮT�E����r�'/4�c�X�oUm"�?� d�ׅ���˿���𞯨��!K�R������^ �W'b��d�9I�Ku�u�R���R�c�����(�u����z��0�k�C����ZE�{z��0�N��f���ax�Vk�2����d<<��?7��K��H2V�r��,�5���W��~�d%���]��JG���.�sW悚���B�q�������n�>+�l��c[�V!+Л��+m` :%�Ԕ��w�%�}bs5�S9t܃vJ���T}	��¼�_��2��m�Xa�u���L��e�u�\�nи��J\�Ά��u��^;������������E��Tq�����/Pa�r�ɿj�ꕱ�,grK���u�}�u�H"	o�+�VFeDU�/�S"��coW�o���{G-[\�͙X���̈^���2fL�ǌԝ���4�|4��d�$s��S2�;
<	r� �ήr����KB��g����+��MISS�*S�힖�ZY�uh����� y�2� WI�qO�Iq��H'�7W�,��noB̦[ ���}�cD���/PiH��w�T�Ⱦ{\'C	f	8������n��K�ݰ����~� XW9��EI��z��5x�ȟ�d��c&d�I*]��[���<��NHe}4M��P���o�J �?<XP��v(��SA��fr��Q��mc`}	k�@����T�dt���o$ϒ��#!Ja�"��*�6��KPPVv�	?����,��*v7��o�M
��Q��
��Iz�ٝ���A�^�\/D,]���I��Н[��4�i���D�����y?��w�����T,���t<�d}L[M���,9`�oF�Ɲ�XxhPz�};X�?����c2Q�8F-zqY��I�k�T!��te����YOU�PbTj��_�G�ү?"n8�=C���_z�ŕ��;5�6ɻ0��!�q��j�:%����R#��T�(c^�����y�Rh�_dQB�MA/�_"ꪂ���{��6�fX9֑�z��g*7�k��f��x�{��%��!lb�q�����L��x�; e�L��>���$KW�]fN��|ڑ�0w�.p��xT�BT�=T�"d2Ϥ��/�6���և��?��{����ίa�_���_6s���pgE��7WpP�?{ģC��q�)�/�U�ir|Sh�rmE��2�@���涽�2t�$�����"���U�hڼ�&�Ӄ�6����-�6�[�\�S�#�Mkk�hԒ ͅ��'`�Y�U��;�#yް�4��Dtb2�kS�/{���]�̍���y�UM̵�A_v柷d��K��T�b�"O%��w��Tn�<�$ƴ�2?���U%;B$�
7U��H���h���N�Лcp�sJu��� K1��o�럝����ߒ�.O�h-쌁��Ji�E����b;d��gm��m<��D� <zj	xV���MĉY��\ߚ�yET���M՟E�fk�޻�(�)|����"V��RfA/��'��D�?0k�h7�#�����'긜��$�u��� O�uu�Q���i�g�$�TvW>��ܫ>�EB&py͟	\K��,��P��`�y�����t�K�ဂ�޿�5r~��O��u�Y��.�g7F�O�vi�C{/��B�a��s��B��0�x�^�4&`Ԕ���+�%�����f&Ro����;K2� J�66e��<S��:��c��dKq�"w/ZF���]��q	�I2�1����~��a���6+��D((ZS+y�9E$��1+���*L;��1�=w���v��� ���?�"����|Y�N���R;�grL���?��xr�ԣ��T$;�O���������ňhyZ�T�ұKb��П"099�����U��%3d�/�d�q�׎D�F@~�~ݜ .�v++���Yg.�N�yC�_S=��6�A캥f���(����J5�������dHg����b3<�� ������;��Һ~��9O�}O�*8|�� �6�J�8A{΍>�"AĢm!DD<�.0���Wu,FV�B�\S�k�~�͸Er���o�e�s����ȸGX�Y�ߥ���'�XY�_x�K�w��c��X`��x��[����*OF�ø��{�.E*r�{������?MjqG��H��@��I��>3���2�"�V���Ą�����˾�3?�}�A�v���(�0Sq��?P��y��~9�ᕙy��`I�<�t��|�
�_c���"@?��pa��!�����O�����6=�����@����S�0�'���
_��|�����ڈ*Af��%�Ca� jmY��֐ά������� ��J�n$���vϨ���� ��:c�1�#�eS��.90H�iĈ*Ok���N��pǟ�R��Į��1&V��Z�6��<�̉R�2t���@�����˄ �̅",�	��q[�2��?i�q�j�EN+m�UN�
�N��-E��j��du�%��|Y��,p�0=�J戋���JL�TǓ�$[��-���.�w�A��v�a�C�{LKb[~��7�f����k0���K��7!Sb\/����I�4�b3�&��q��:� ��r�f�0�<���k�"���<e�I��!�	Ub���F���������	���<�N��{�G��m��4:b��'���'Dܕ��� v+�5?�l�ѵ*�'l�ѱ P ��|�>�X��i��t����7�喘#��A3[R�����<��4��n?���83�"^JͺF��"�����	�\1���D�G�DE��NW'��Cl���/�aĎڂ��@hJ��k����k�S�G}LM����M�X2�!��h(~�ƑC8�p�f��M���m�ڥ?�<2���1k{شX���;�j޹9�@�*�L�����T�O��� �P�w�(��i�n��*���B�*�AP�E�_,��T�,�랯5�d��0����z@�{"'G&4^(	PǨ�&��n������[�a����Fg��	����x� ��ʁ�G�4�(�����[�A�9#�fP�+k����>��U�'��h��o5�/8l�>p|q��.�޴�,5�_��U�lvӫ
r2�w"���d��e��u�/�7���EvD-&�Xp���d�$ֹFI�'��ޗ$)اgFyHֿf5�����;�P]�LુRi�Ys��`��6�FM����؋��������]����~���1"����������Z�졉C�����E~ֺ�/���ƾ�; V�6}z�,�0��~��M�YS�HA?���̬�f����ƷBI=}�p(�����*j�[G�jz��� �{u�96��2&�r>���_CWk�^	[쓬��W9+1���IZ5Ǖ�Vi���8��r��.�T���|��({P�HQ>��˨8�w6�t*Gt���gZ�[ŉ����6 ELM������g�i�����6(#������H�t>ތ9fD�d�C�x��^��P
K��6����3G��,ᴱ���:u��;��|P��G���W�?#wUJ`�+�{i������j��
ܡ(��Ŵ�b��jF�>Bu��x�؆���Yj�F,,��������yP_{t���
h�@��A���cR:G�jA�o����������D�\q�&�H��	�v鑈q�
����ۭ�1ŗ`׹g� }�*���O��_��K0��4%LK�"�dog�f�&|�T����K�xjj'6�ϗ���S����M�-��U�ȌT����zb��5��@h-���h�K�VT���&ɛ�"6.�{�3��yF�`"�6��'7�/T/Fz�����)�쭗+�Zi�𤯸F*͚yʹ�Ўͮz]6��ܪ��4>����;_������e�;���`��|�ڎ<��X�H=mɕ@i�A@/2�1�l��vU�]�*Zӎ�^Y��hl�S�u%�� �i�D����l�Զ%��]�"�1�RPɉ�R�ws����������c�O��.�xc�7���-�Ȉ���]�1XG5يp��0L�3sf��
�ق5fJ��J�SXc�F��^vud�xZETG�_!���itY�R�Og���P�ܜ�!� j�mz��j�v"{��
b^�{���!" )_v���|,��R,G��ԕ�������|���՜Ph
o��������h����U�y���	���S=im<�纖1�;N%���,/p��]�ԥ�pjw(�%kZ�T?���vG]�b8-v/�ջHpߠ��9����=2����vYؑ�1m���K�ʸw<<��2
h�9Z�U|s�Uo�Y� �5��8��36����%S�{���,�LqVq^S��f�3�pτ������8}L������B(�
�Ζ1	�*�;,�i,]���˻Q���^��=Se�#��Մ�>m���DسSџDP���4�+��I���.�Ä��j!�������-������
�Ț�����M�1�2�,nY鎊JZ��cwDb��H+�D`)�)�`�l�TZ7C�TV�pb/<I�l\C%���E�}��0�x'��v��j����q.�N��~a����q1���I�l���E�q�-�|碒!� 1�!BD�@���~�B�i�@�\�|��]7M����=���ĺ�BZ��
P�3
���!���� ���N�u��M���<Y��0��G2�L��c�P��e��W��$NF���p���ptw�@?��;�R�����5?PY�t<2Lf�GU��1�礙8�Z|�%�vj�B��6��[�>�b�l�M$�3Іo� 0�RI%�=�J�烳I�m3	��3u.>��ki��<#W�*O���K��gK.�,ri
w�g6���?��K��(����WhwS@3հg�η1��W�1�;�]7[�?ռ���z*��rF�_P��8ҙZ��q�,m���_Q?��7}��/���i+��9R�o�9��Q@��?pX��B� �N���LP��%6��c�A/3̡=Ẹa/��Z�-Ey�:@a/B��HA��K���Aꈄ�D��"s�٠g���!D�i��$�4��N�4a��/�ciu���(���o�g<��{�-���1��G�زi�n��AV���9 ����S�- �g��C�uyQ�h�~��K
�?�����|�a�p"}6]ߢ��+&v]/OF(\-WD .���xb�^;���[�Ǯ����n]tN菤�:������(؏��*=�q����6��-��\�H:���

�SC@@���C�&�U�9�/3;��.ڤD&L�
���](��Nճ��T���w�#l��[ћl��)�;Mdg��2��8�+5��������"Ru��F��&A��d,,`$�i��kN��f��7��J&D}yl��Y5��;��_���ёY�dG��n��ŔC�X�mϤT!-.���^ o7>���ΑE���{h'�z):&4/���)��*; �d����1'\��]Fl���=D�n"KDWǮؽ�wZ���ԕ�:��H����z���(���Q��L��p
�%UB����E"��W�Q�҃g� �$��4��U��{�}�6�)O>�e�AJ��	$|����h�ǅ㌺��w���1�x�p<o����*#!y=�y�FF��l�֑������Xi�S2�W+�~�W����~�h.P��z�8��{MC���*���-� ����<�%�5�����d*N�v��p�o�$�OP�o�k��������ݹ[�"A�'5O���Q�Yl�f�.���� �����<��a���ʐ~��R��M�ƍ�DU4�����]~z��<8����\kc��l7D������v�}*�D#Aa�Fy=g,�tH;ɭݠ|��}���7�L�M@'�ы�fi�y�+��U����Z��_ ��S4Ы+H�����f��/��ۣ�?�%쵷��0�yd����U�:M�US�5�y�<���	��a�/G��s�!�&�B�3#(��}����2����ĐDY��L*۫�����G�����bx`Ex2��sU+�8+���S����q�U�n��
�i<�~5s͕��/�!����V���y,�\���h(�����壉QV�f삠��_D�fRF����dPy����Y}�D�g��yf{iݜ�g,~�5\r�S"�!�'W2{�>�m*S��S^�V�t�>}� ZD\�_;��+I�g�[��y�Wbh�W�Sm���tge�t�T�}II*�9�9���t�0&�@��t�����*(�Z�J�a	ds��ن��e �d�7��F�f E�(�E��D��җ4!nj�b�37�jC����=�.`aF�*t�Ҭ��~씪�O8j�G��4�-��l ۆej4)�_oav��Ay���8�Ln���$(�9�=9aI��$����HD���5� �yD�_�rNѰ��r��T	�A�?f=�	���m!I�Lm�]-]%�E�껣��K�$�����F)n�Md4������5��5-MW9��y�����QlL�,��c��;֜����>0Ӏ��uWu
Э�g4ȓk�i�
�]<��Kf�P�$���=�T�Q'}���V8 d�:�Yh�w��B�6���F��s���5_$���[	U_�Z���0y0a2t���b��,�R����� ;Ȩ��o��6��	�A�c�lM������`933'1`���#��������}gaɳل��Py�x�dUH86if�}S�f�c��l�=��ɓl<n��;IqK������&����
��e�SYB�D��H{I5�	;<Sq��OL֍:�j������q�K�F����R���a>~c�=����_^-����~v;��wi� ��/�
��3��N���7�3kqF�h�k��\ox������Z�����j6. 	�\�#���I����th�ԁ?*,%�w ���,�_W�p~� ƌ,�Y|��,]��,�������y�@'L�C�kkR��M�J��}������Z�������c��V%!�ve7Fan��giu���n��H��.E| �����dJc�}�A8��N�Tn�Z���v�O�>,��b8?'b .�Dk�x\Y��qƘ���x&�͈sf�Թ����w�R�\�z�HM��A��uyφ�E�Nm|ȱ�L�}ߩ0��Qj6���#F��fH"�ݻ��J:K��tK��U��,Ư��}��0O���loe�|�͸i�6���w���o�Z��G*�b��VH��K��6��"�4ȋ���섒�
��%�$"R� �_�z߾A��P��{�!�զA	��ؠ+�XϤ�y�)��ZC�v/� ��	��IX��'({dv�<��4��0��"����T�����ISTF���ռ��W�t�w53�v�E���b3{�Y�I�)IO����6+�~���S���[Tu�5I�_�L�}���i/�}~�F8m��c�T��/B�梁���y�5�^��:�T��e сg����o����w���'����Ei.���W���lJb����b�
,�54(hŒ���Ƙ��������.t���-n2G������˚����(_�M�ѥ�L֛���
��Ǹ��̔�͊t�������&��p��[��D���W��'Y8��u:���ǖ��� ��<]��5~�*��ٲU��é#���a�Q
�(��U���nL�<�D�	k���HX�x�m�L�,n&�x)����*�U���NuQt�����Tuo���f�1��T͍T<��~��ټ#Ou�h3���4�
�qO8^@c ez��󬖃�L @�R�>ձkβ�AA�����$gЈ���?�� I�LVDh���Ѩ�v�"'|��kub'��0��.�4�����.�����¯0���5y���/�����c� C��ٍE5E�������d�ΐ�!J���a�C������؝
�[c��͹(,�����Qq�v�_D��PUي�D��rȋHз��l�Z[^�-�f��C!�Ƨ�Lh [��I�i�?�7��a�ͽ����M�h�9��� *���mT�l����E[��ʼ��|��檿����U&��D�|�&�2�X���5pv��0�h	�{[kק� ���\ѳ�Ӣ���7pF�|���{��ZP?�O0���ܨ�#1f籕��&R���s�[=���5��ʓ�=Az9&G[xC����Ե w�h�3p���h*���?����3���<Ӷ�S��M1rkj���*��T��LC�0:�l��}B]���"�������ڥ�k�n��%�ޅ�9�50���{4\1f�`_�_����v��3��v!F#��Xv��t�q��S�2nPm� �h� �'�z$Vs|���/.�I�6��<��D��*>1*�2S{ّLދU S�?Y2�}E�>k8UcW�w >��
�1�U�Jq���8%�%V�>�Ok��:!WGX����I'��[�K�f�?��>t�~[H����A��Sǡ"�MsL9����D�{����:4o�i4S�0�d�0q�נ_�˝ʒ+<>�H�-S;����(���w��M;��^P�d���#�Nw�rhGN㊎�5��p0�=�!*$���a�c���`<Hz���ۥk?��{��`G���pu�S��0�MiK=o2��\�t3��ۓ5)�F�	�<�ۍ+gnk�I���o$Y�^�e�g���Ru،.���7�7nϵ1!l� ���Q��'���b�/��Q��������<����%��W�<�Y_�a&�
z;�_f��	�Muώ�O��n��̹A�c^E��94�����CK-�W؛�V���=��_�1���V�m�%a<+I��0�A��\o�X��pm�Fd���S�c�r!Ǽ�&��Յ��/�,Ҋ5�~V��^x��!nh-,:�M�	[��	�F�����[��*���8˛�5L���ܸ�Oh��g��&M�b2'!�7씑�\q�/���K�H�g��� ��YnV�Oj,�]��g�G�����-6䏨��psjEu슊RTN=�?��é��I�2m4�"Z9��Dn (>��p���M�%��ݘ��
�`f	�se�,%��w��s��$�����T�Fi��G��C�|K���_�
�E�*��� U�V��M�wo���f�d�-B�_�2%���,�hv���ܓ;րa��ӛ
�j�=�<��!4���t,��JO�h#�j��;}���J���� �5�d��7�������WAx�(��󯔊���d:���Qd��X;"���@�d���ڞ8��g�ܱ��M=1�h����յG��%�k�9 ���]��z�_t�&uB�'=��&�|�u�Umj�?z%�bU�,��x����j�1�$U})%Q!�N]�����l�jg�r�uy�{(없�{{�d7�S��ؔR\�3>!���g?D�H��u��.SZ���?J��5��l��$�G���^������Em��e���^\��E Q�U�n�	[bI��_R�_����䮷��Fs��Kv9����������j%�o�2>e \(b!��.����o����ͮ4�"�~��\��u�A�@k9߰�
'6��M%̿�Iƫ��/�Vg��j��B�;���Ҧ��L�c ����^�qOc>��,fkJ��JZ}�I$	����7[�k�X]���P�y��Ҁ�D���=FM7�Xh�%C���#�v��� >v��G��t�L�A���`:�ӥ���,�-�C�R�i����m�C��8��N{���Yry�1&��m�k� !ko�͢����d�y��_�Ɋ�>ĵ^rA�x�C���_D��m7��7���.��<��݋y*�.���+�)�NJ�K�Hy�=�g�*xz�b=E����|���D��*-{�[w�6�P�WY>�3�0_�x����P�����ya�*���^����Ot9��t5�O�I�M$�G=3d�T��n���o��������8��N
�mr/䠰��q>h�y�x�;�J�J:D�oG	�Q�ǧ�'HF��u��_
���z��q���+�_��Q0��dESp����\QP������ra"G�ǞNN;gC�Mf����0���,v�Z�Xi`�6=�*�rg��4�;Ffg�"$5�����������h��P��Y�n�P�*�j`��A������
^i ��vKg�ѱ}�m��Ց� �{�����`N�F����6���y��x�y��<	��YǓ�) �V�w1Md5Yc�eƉ�Ƶ�](�88i�!�P�&i']h��B���Eφ�W�U�3n3,r�' d<-�#��@bWw��?������M�7s����n>�w�Z�d����0h�$�T\�Դv�ød�N����@����╈|���{�4b�,��aib@\��{��vs�l��}fٔ�3k�*����rE�9/��i<����9!x��a�B{�?t���7�����e��F:hF4������/���� 6=4�Vp6S7��D�i��h�,�΍����`�P��T����E�3��Z�?�3D�}���]�W�e��/D"�G�:��,k�S �f�9c��O)� Mu�@��u�!q��0o��ֶi�_�x��B�MdW���A�&����'�Y��2T��e�B&PѓMc;�o�qXt@��]H��h�D �Zl���@v� �^Z��ʨ�A�-'�u��V�$+�X�u7��$1�C�5^��_�c˗��(�p�$pR�ަ��R���Y3�N��*1��	r�����,}ܛһ�����)Z�RC�x3'&�ݖߚL+=���|wD� ��
2�\�8?h�����&&�C�߉��"�3$���<��t�̊+�=h���~�cml�*��š2����+MC�t�Zwc�� $�xB7 P*,���N�c�������K��}�&��	E��W�'&�-�+y0��ݩ�L�	��p�`g�:��o;o�;�A�[O���$O� M`��0|��bߢ�xb"�'=3;�Ow�o���Z���?�J�P̬I���	�AP�����P��I^���������{�r�x����i�L]�W�f����ck`�����*��n9Bg�&�q�־ܔ������l���*0F�d�:���Fi�!+��6��x	qJ�����x����4��6���������i�}p���ؕ�^�76�k^?Blڧ7��]k�Z��lG �/S�����N!�辱����M�2�s��=��z�#hrh����'M@3@k�w���u�X[Ex��Q ���}����Ѩ/K�ie��N�4@�p���f΃5�,{����Ip��g��`j�Y^�(Hn��E���o�AKڄ��{��n���t��=Uq�k�{�R��}�Y��W�0���j�:���{V/�
�V���9e�HOj�����{9�ox�1ggr��ޔ.B���2�џ\3��ze�g2+O����Z�LhΑL�JҰg��1S�-�x��`�g?��s��d�9F���Ʒ	��`yAM^��!Z��D��a��/d�f
�ծ�?o>���x�w���O��	���W���f�A��n\Q�Cu_=�W�Y�3mn�_&�����)�HhQ�YL��U��"�;Ir��Y<Қ��K\�Z�Vۋׯߘ~�a����84�D`%=�6�*�B	KEv���6B�e;hjQ����Ŵc�����#����֝/�UĞ%�
�Mbm�Ԡ�����F�;K �t����Da��E]������A3��D������T0VKM�a
+�ʬ�I�3b�$XCm�=�p�Rc��Yq�u"B���������<�i��,o�'G�^�k����3/�a�g�$���`�ٻ)�D"�Pp�Z��$ё��'�h�iB� �b¼���!������K����13�.�q-�>���A�i��B*�ޥ�x<M��;��_&�ć&��e�l��-�b�)��;~���;���J���o�杇S j��S���� ���h�K�:�ĸ���/<4��UX��	��Ȃ��Ye����L�-'H/�5�2<��މ��z����'�Tu$C&�&������lѵ\|k�eA^�hG�9��7��)牨��h{�OE�Ba�� ��p���=�d?�\&�Jh��:��Q��� �ƾ~ڦ}���HE�uS���m"hT��ΔU�H�YdF�}����'�]�����U:�X�lq���m���1ci��s,�IY�PH������u�6�O�	�ʷ$?s�֯>���].Krsj�ƫ�[�^5kP��,C�V`?K���$�Q��c�{�삢{H����E��i��Z�{3u���R�aQe(�?X�r8�g��g�	�R���f �s6%��cl��������l�"�(���{��ɪ��_]�'[�=y�-��KO\�S����V���iY״�j��5��{pf��q���J����X���׳���E��K�u�=K�����m=��ƃB�	�y��|>���M��rq�B�*":=��|/>}�� \YX�/6X���Q`\P�?��A2�Ⴏ��%U
�\�U��u��y�p]�	�(&\�Y��0V�w�>Nh���1�J�����%O��v\m#��ePń���]Q�Q �S|R/��7.i��(�����f1 �JnE�O���d݉��M�]F�U\Ξ����8F���y�nd�7�9�ω5ZG8�w)���S��#ڤI���g�v���g7�O���������mOZY`�\�ܫ������ߟq�ɷz�%ٰ��:|���K�����KN�@�%'Xd�ӡ��9��ηiB�L��;˰vwe�x�dIj/	7��[�L�f����]^����a�z�<=n: ��BǥP�����>"1k��g�z&o��n����>�B�z���
�F[&�d���)��$[Њ�S�aN��ϟtE�̶a󻝵<�~���l�R���!2ZzX���_%�
� ��ݦ��Z��y��e[t�C��(��ڐǀ�����{�v��f�sÉ�
nW^�L:]�����8q+�V�K�1C�К�`b⻒�ܺD�L@k��R���&�[����ˤnW#�-���2`�Ma-[���3���Ķ�kO�Sm~�^a����2d�z�n����7<;P��F6v�Q���#S��w�RQa�R����u�]^,�W!��ä#i�|����	��a���t6�L|b�Nv����5�S��{sⱝF'M���MO��c��fs(��L���E. ��h�������Lø��3U�WI�ߧ��%7�f�Y�T�&��@w��bsۉt�Fy��V�;�����ć��j���x��*�E�}�smkږ��v]2�>3�?2�ŨU�fM`�E�ɲҹ�I&53��B b�x��&���X﷝����@��\����od5�n[��5�b�ѐ��hU�h�ޅ�(̡���g�GUt�9��QW�� ��k3��XR;�� o]%Ӥ8i�-������:a��"�P�,�1 P �1�n� ����+�W���aY_��.>#��������7M|3r�8��BVr��1z�F��.Ѳ(4����AQ���"�'�����)�A^�y�M�୏E�/��8�(F�s�I�!���rR���L��H^�ş�g�=�D������}n��0`g��1���k���(�ϳ�&�i���hz�+�*K��^�~��5.�ړA$,���m���;�kd������OwF�wW� ��Xo ���;�.��7��2�����E*(�p:z����o��o�QruD�E�M�iJ�{CEv����<"�..;:ma��m.-�tt�,���ߴ�U����t�2�D,�l�G]Yru���Ut�%R�>�TӍ�a����)'�����QA�L���>�W��7!�*a��<ic#�역�|*�0���^�����^���v-	(�Q��{�s��o!_o!!�����7X� �y�$
mw�c�"��5��O\8����|'�i����ҐM���D�mi����d�au(F�|����ϬH����at��.�k�tC�ZƗ��P�����s���f�c�2���jOG����)������tc������[څ�1K6+��F���Z1P'�-r�m1�E�j�����"�P�53�vz,��֊�� �� x�@˥P{V=9B׷H��:����N��E���ٻ���Í������a��K�V,�yN���H[j-�F��P7;�j+�EU�!�D�[�d:�{�|��]��v\���-����	9�s˃xw,
>T��fpK_�O�>��>h��/T^`篑t��,1��{xM�����̧���j�ު�h��a/�Lhl��Sj^?6=y��xDj�Yȹ������3r�
 m/�ϭ���Yƾ�k]P�tO�c� ���G*�Y��$�O��5U�
���㿞��Z�,[��q�~Ę5l����Gk�f$�X�Z(�j��+�j�Ĩ4�s���l��r����=;�V�ZDZ�������b_fs�m�!q�#s$&ٴ�4c}D� �a��L$_V�X��]��j�}�G��b�"���>�.���L�9H>f�`z��0=�S�ֈ=��#�d- 5;��D�*'�ֺ>R<<9�JI��It���0�n]�d_i]2[�T�˽����?Z��P�k/P@��S���Ʉ����~oM%}z�)��3!���
���U���
-]JMb�����]y8X(6-�sֹ�P��kS��#ښ�J!�J����5�2�4)>B�&Z��/�"�:��2�G�7��<G"�ʃ������tU�!ܹN���ep��}E{^�y��Xݬ��?��JY�/[��"9�s�-�����Kh���W}�.Qc��l�A3@Ѱ5/�% ɶk�`�|�d/s�������7D�l�
�]m�.�:�/�;�1�a���r�BP�X��_�m�q�D7@����3��T"�^`��v:L���@�qѮ�K1�D�~4�1��c��2xZ%��L�`y�,K�
��u��;ѿ����H��H\��$-�>;0:b,��Pͷ����5������~��1�/dh~�RG��k	�k_iJ�}���s.1JA��.���z}7n��{Ê�;J�M�����o�eּ��;&M'8˔ٴS����������s�r�8.���*�����S�@��a5> �
�	@�u���߶G2��ORMy+�߲��qh��N�O�m����ؒ��Ȕ���R���PǃeCk�����Y�υ�"���x�H>���?�s�˹gw�}��yh����ϸ*ض Xdz�Y����HS��\;ݖM�0FS����sr���.~�bS'��x�Q��Q]L����C݉��ژ�9�I�ns��+��:�g�N�'�/�t����5.H��P�<�a�YwR�mP�{���8�$��>"�����o�5ƧD3�}B�1��{w������츉��fU������ט��?�ǕJgh�m�S��d�\�$�@G�ԑF�T>��	9#%0Av��/h��l�s�<�a��A ګ7Z]�� �d�L�Ĕ?1�N�v"#|�*�G���A�T�k�T8��HA�Qϗ]�=v���*��룱�:��Lu�[�Ǻk�g��A��gz^;-��b��<�r�zDxqξF�Ҟgew6��Bo������n�0e+���Ȑӧ�_�����]���e5@�@V�T��
��2a�����=��z�(A�]�I
��$�ҳE7H���A��8Xi/��aFq���a(��BlL�9������������>&R�����E�%׫��ȱe�P���dC�^�f9�F�PV@5�CfAH��KwLe��mj�R�xγ���Q��(Y���n��vNU�*�K��6��j�8y�N���YC;�ȏ]B�п� ��3[��T��u[�̊㩕�}�\��t�\2�n������U��_&vI$��7:�L^	��V#�T��)]t���ú�
���8W��,Y,���/�AKb�3���mX�ݞ�m��F�{�a��g*~/D���na����n���HD`r"4��ju�A�z]f�(�#o���a��E�W3^��ү9�(蠲V�jL&�(Ӹz�������Kx���f�ɲ:'4�U��B�7�k���]T(	��]5:.��rE]������u����}�9����K?!�?,�1��a̯/+�C[����f�?�0=��������&s<�ҍT������$��-�X��� <��6���g� �!H b�ӛ�j�6z�<����D-��&lZ�_zy��u��RWl�M����9ÿ��n���7/N��/����$���ht�cy�l��7mV�5)ϝ��<ʦ�n٥���&���2��d�EIa��=ug�ɕ��WK��-r1�$vu�ڛ�#b{\*|Xd�c�9�5�2z��#N�0�eBo��m�_2�GF��2󿜧�vѳ,�z�D`lT���z�Gv�ƴ��]��^,�L��+闳U:�\���X�mi\7���+]����c�f^QGc�M$Y��!q'�U��ۧ���+2|Xl��bތ�?�m뙯�)�HlXA^�o�d9|(�SE4=K���Q��ID��Z�)9�oIY�1�AJ4�_tL���j{7��|�M��y����k�ю���Y ��5Y;	u���\DGn��9�	����f�m�{@���?��:(�]�ၴ�mG�6���b���+3F%����<$�d�j*���UJn���bF�j�I�){P�&�\Y�@԰}���H�*�r�%��+����'���\�0�5A/���v��[�P�%A(ɩɦ��ּ��)_eF���	��&��a���DzEav�{?oe�Z�BrX�
!H��dk!�X�4.�<l'S��\�շY��89>�_��j�yµ��a.4��ǻ����2���@%��
M�&D�ھ�#��ب���G�[_e#�W���+p��{�9���@�]����hl��[0�VΙ*=��`y�&Y�{ybE�$[MRT�;¨=��E^�`�� �a����C_�+])e~��<�(��
�u�]"A���8!���������ٞ�����/���@��߿ ������a���	��19I�T��m_�9Ƨ6�j�+�`�iE�7�@��>I7W#Ő�N�[&��J��
�_o��6����3��*��2]�ݸ"m"kc2��f�$Qb��G�6�m��[�Y,E��Q1WȣD���DNt�>���{lC%ʕ�9���g!2=�ZT����k[�ԈwyO(�t�O�>�j�9�Wמ�'�0�YTQ铜�Y1a�ȍ4M���D�������6�;����W'�R#�a$8�{g H$��&�^�&j����5)Ɋܗ�[t_PT���j�3Fɠؔ3i9��U�2�2�^���w�۵�f�G��u:�:�è���dqaQ��d��*�9�`����<N�U��ID��~�� {�.�HX� �GA4��ˍ'hf�ɾ��.�9K�!?�Hz�Wh��X�4��l��*�T��c)��t�"^�z̈́��
�$���u�9�r�̴�.R-�qR:v"���	�fIWL�J/�� �ߨ~N�~�A��9f�z�(׉x��ZԀ��v���@�R��k����;ce(���V�jP���'e^"x��ٞ����׃wq�Or�n��.�gC>�Nn��e?��_�����0k��C�I�OM.�̅
ׄOT�u�J�\��J/_#�_D4B����E�ԋ��KylmSJ+a�h�}��Gީz�*�~�rY�D_���>����Ly����/k������4<z�j���+��7m��ٕ����x{P*��"��5\�r5����ܡJӗ�!,kM����d>#�!��� �{��&%�����F�}>��sj�a�#����\�Cn��U�
:W��1,��Ӆ�0A��	��Fi�U�9�UW�K�\ɇ�(}̭sy�Ϟ�b�&��~��1��NI���q�^+�Tv��i��}0�/;@����%��;�"V4z	�[�a���f&3~���_�����[ڂ�woի����È%P�@���;�?�B~����eY8!�+���[�B�_��J�	�YW��۩�JN9���7��!	��\�v��V1�)������Nǣכv�GG	�0ԓ`?h���Ig-L��2}���w��t -����8����+\e����R	.�� ��LS	L�ҫw!F|y$<�%�\QW�f@�^�0�F�sB���i����4��r��
w��{��ln�&؁�7ΟOi���Yq��p�:B$��������2��3H8��RJ����=��\P�S��+��!1�]H �Q�ڑV.A
)P�mzM�d1@���]��0OI�e�'f��X{��w#�Ex]�wl��I�ߌ��Ȍ�L`�о���'m�2W����ϓk���aE�<A�b�l�x����<��cMs������Դ�#4B�?}��R��� $���֖˃����s>��-j�� �������F\ٚð�Sg<��i4�����,���j�Q(o�`��,Ǽ��G	�~��@�x�Q;'���|��у7Y���#g�"���+�{�54�9�r���ot#�XfU��R���WtS�k��7�^�ɎDQ�;H�@�]�]7j(��eh���-���9����8���qvl�g�����?di�T~>� �E�F�lJ�0p�Ȇ�6�	&=^�+7D`��M&P������+1��v!�.֢�5؀�7)�69�����)�oK�9^iT��J5�F���K�U7пc����~�e��� L5U�!�۬vZ~�.S�P\40}$V���y,a8
�G[�wa�R�g���yl̝�?h�%��`�h�B $`�ȥ��o���1��p~h YF?����ɴD�Y@-8�.�m�e��Yk���]�����������><���E�x����14�Or/V���с�2��ڈI�S����rT�����i]���a�1�|z{�R%�/5���I=�!�@��iV�w+X9��1K&~%B�u,���c( 6F�x��"��+������;�u�=�+>FtU�"�,Dz���;Y0}��	��c,Z�v�O8����N� �R��W���#4j�ҧM�*�4�o�K�ҖM����v�����|�f���Ai�g<�]G��'�ڏT�wV������G3	��֢W�c.��w�y�~6�;�HuH��Yε�:�1GR4q�ϴ7�a_�������~aq��U"'ГG��\0�δ�w�q����ց����yA��$�9�SJ-Ӣ����&��ȓ&v��Z�7o���g����\�F�9ԋOaҴ�Ex�Z�\ţ��m�h�G�������?��������B~Ѽ�9����d	��A }-���!J�܌$>M���1���1W�T������3 � �0xTly ��6��1n��hV�	ѣ�gs���?Վ�:������n!ߑ[�귁��Y"}U?�Eζ
@�E��nH=��E8�<�̔�s;����w�7�w������e�܁�AG�&��k�\�="���Mߐ�~��Y���H���#��e�������($� ]��
�tb��eF��!D��T�Wt�(sw��p[V��lW}�`e�^��R��"�Q��>rf�݉("����R "? f�|�$����+å��H���<C��[���9���f�\��U����g	���]��t]h�w}d9d���S_$�
��e��M��i)j�qz:��yge�Gvi*�\��B�)����rD�u��$3�N|��q�@�1{cj:;Ģ&�[;��	1��0=a��b��YJ"(X�l��@���k�9g�v*!_"�Oǻ�Hoe�C风 ��u�l�'�Nԉ#���C4�ʥ�����Ǔ:��zS�M��B�, ��������43����~��;�dU,�Қ�FF��O9{-��-l�S�D�)^O���'���@O$��unps_�<>2�wd�b��<����a+���	�ORESb���զXR�XYU���r
� WP�ݷ8�e�X���Ŝ�0=��|Q��ɕX���kJuN������[�ljF�5J��^작���>q��7#���a�ɏ�\Fi !�l�����ݷ��QG`�q����w���h*���xr-y������]�'v3M�>��i2�4^��t��%������p�'6�#��)Y�eO}t� l��O�~�����|V";W���ߛ��L��_����p��#����'�]pJ}��#��0br��5\4|e�p�O՟�/YH���?�#���@
O0�e����O�[q�gf�B���˓2&�� ���E�:x�|K�����-��|W�����ۍӷ5<�J�4�w4����8��:��	zd�N_��h?x`R����N��~4wF�:?��`CkR�U��;��|�m��W�Ennz�v���Y�"שʟe����n�!/�V�X������(2N� �u�dB!`��t��&�!"$��U7�;<��#i����<����	^�O����� c�.v�����y��!c�dQm��I�;����1gk��Ah�8�>l"H-�J9pN�v��=[�����T����ۤ��V���� ݗxH��6�՟�ʬ���5oü�y�a^��ԎA�[��D���Hj�<# �i���"�B�"���[��ĹA�и�x���˄_t,_&��><��:����1,�T��@:�0�9p�cRqx�|�{W��Z�$�Y�(��r0��t\g����a��i?2O�Q+�c��×yD�����^�<��U�J�Z�J��J�w���<t������OQ̲�ՅkȾ�j*�Y]�	�SJ�^^'�!ګ��M�hH�ys�7���U�}�����o'_��%�]d_g(G�@�B��$�R0�
����X���W>49�>�q����tv�pY���Uc�i��kn*�&x�7��F�]g�lN��V��@�nNO��O�����أ44����ȂJ縝���,�?5���u���Ʊ���m����?j� 2�����+e��>�e�̊��olі��0T�l�b��GVʙ��ou��r�f�2��;Y�[�~����0�]���%��	�* �a9�i�~�����"�f��_ZC���1jT�g|���x �m�kG	����Q�Xr���h`jDM�����YK�Q)�HA���e�to� ����r�HKaҔ���d��������u�<�<��X�W[-�<�|L}J��ň�C�����\C��۠����to�5>��?e��|1$Qa�B�
I�؝�3�
=Qt�x�{X~�(��VTڬ40kq>+�*P��Rb�0��SK�~C�sBzd)�������&�2�87�����*�:O��E���J}+���};�0��t̎��YR4:�7a���|Ni�����d�I�m���l�d���S&�	�z��WkJ������^���ϭ����ۼ�{�v�y�Q�B���[!0��rsV��mWd� Y�V^��j)r��E��̏C����c������m����ʩ��n�>�����A�اB���9�ݸ�)
3E����c��\�i�h^��J�gm�"v<^Q?y�S�R"'���! Z+O2�&�qd/�����3��Y���[qǟ��Fq�Vm&MY-����O�ꀌ,���H��'إ��Ӗ�d�̌�_͔A;�����&���vT���!D����G�}�)�>�?�k��Q��{�{ s�Fv!-IӠ� ��n6 O6�0m�${��j��t4�y�[��D���m]X+�y]��<M��#���@T�f��A| g�}�Q'�_��=�.Q�"#��Ԣ��������ho9S�����Ѵ����<��ܰg�j�(�����d�"{oX��&֥�Z��-��Ė >��� Ϡn7�C�-�x0���g�����U%�1Aն�-o<�i�T��i��#�{I)YY�u�0t��p����xr��gd�Z	�b��B�,�?`CBn�!%�vg�]�Ea����-���c!]Шզm!T�Ӽ��/�e|��V�����x���/�ؑ.��c |���q4�Dh�WN��S*Uy�&���*����o��sW���I:2�u/���9uuT��l���y�H1xra�E���/�q��]Fj~)���<��fße��;�}�zl��}��5��&B�"�n��������ӹ���-1{��P�a���T܅t�ᕑmz_�7%J5>�k)�P� G��|�͡42yq��&F���d͜�Z۟g�˳�HA�Ovˮ4�L�VЂ�P���M>��������g���0G���I�yLAB�y�=c#��d�&�䦰齰8�13So\��\>n:-��o�O �Aw.�y��9�]�t���<5�p'�R���(6�톽���D�59V�����FnQ�&��WS²��)Ԃ砩R.E�
�������F)5|OL(y�^+����\*��T+���6]]�R7���<���c�54��<ՖD��b_��_}{����*�Y�I�v6åQT>˅���?8�	�
�ȾȒ�A6�?�ۏ�3��q{z�7E��`�U̗�#�	��)�5g�0+��K�b��P�oT���ϊI�����f&Ji��F���S&�q�k���X�p��_��BXQ.DǓ�3EU=\YU��2�2��Y1g'o��������-�|��bh׷�����)���wu����V7�����.2�7A� \z��NQ��� �ĐL��1V�u\���PK���'/a���w��7:hΩ�}�I�wr}�"�1��