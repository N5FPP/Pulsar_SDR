��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@���$U[H_#�/8�y��,��F��`G�m6f�f�aiI`������tC����dl���=eZ��^�٭����B�FYĸX�G�����݁�]}~�s�cC�_�V?o6���p!��#��9~̢z�x	����M�8�DӅ>q 6��n��  �	���Oi����P�ª�ج�9���Q3��eS�&�ʟ۹����:�V�ۂZ/'m}�Dv�Cf��)B
�n�ݘ�I`���e,����i�����r���+=���%{��V�ݴ����{��L�����3,{���<�@�3��N�0X )b�t��~����=����y��(�l\�m\���?��B�*"Rߎ�R�ʃ��t�6
dw=y`j�2�e��J������^��ò��-ƀ˘��yqXy��1Ȓ��h*�׈��.�T	森�y% \PU�*AH��i����Q��w�YH�#�k:����db�s叢]����8�Q�
���d]�5�h�Vr�(��C�c���¸޽`f���Y���#�:D?��.Ĥ_��5c����D�Q�{\l�M3�r�������
n��b�������6AZ3���r���%���Ly����7?i4p@�tƛW "�o`α����n0��dv�qnh9!��П4��[� k:{��ERS4�ۇ1"5�E:ԄxDL��AFqDu ��b��e���6ϛn�?;$�=_�t�s�RL8��""#�Z=vv|�g�t�嗻CYY���m�n���
����|�E}������aS0"d��*�q��h��a�9��Xy��1uY-6��Af�����F_���Ԩ��|�Ч���_�y��\ g��H(����|�&�D��F���Vv��&Y�kP;T�7چ>�tH�w[���W|��5u�S�p��[
�>���B ��{�t� и~h�j,^@0��Ƙ���(6�ɉw�ި�Q�D�je������g�����M��i �+�[b�d�rV��q���-?�靋`�:��q�[�&5^���!ؿ�J�5�r��[�,2��y�����5�Ts���D}Ag'�(�'�z�m5Q�D��\��R�@-�=����3]�7�f�ރy��:n�֔�W̤�/7c�~�
��dK�a���+�92���M\ayޟ߬��M�2�k&�yt��7<��2)/5^�+��K质Dlҧi-/��^�~���_WR��Y���%R}d<-^$�����+�3R��׉e<NH6qB{*n=�hCOQ��ڣ������qqK��x>b�h&uy���|;(yH\������{bՐf�p�/q
AS|�uv�ځ݃����ƀJd(U�dv��k����)ΰ�(B��Z����L� kygde�klz[���� oK�n��\��0����8�H���3��j#�ᄉ=�0]d�T8.�@�o"he�q�B���(�ә׭+0�9�����[C��J���ʊ�AW@f@��Ǎ��~��O�t��xď6r���X��X�ޗ���(�K���u
6�n~��t�j葷2�C�+V����䢉�m}|���[e�r1��Y\Z��]庎w��?[̞<�	b#��?�YUxuX�.�^�aX�$�SVӫ�o�~U��cٞ[e��\lT*���b���x�>�+l�^��K��n��� �_����z��e	'Z���Q8�­<�>�Y�tZO;������� \
�Z8�Ȟ-k8��ի]y�m�n��5�fω��:��MX�B��BH�?��ư�<AE;��j,�F�<����6(\(�/�I�ɶBvZ&�"�}��ܱ�c�Fe�e=�}ѾC�#$��\F��@E���Ti�#���Y�H�Q�P��B�N4ݚ��5��J�1kJiE� ���?(�?��{���*�-J���bŢX��O�kgD3ٷ�w�s+�[c�+ڙK�EC��B���&�����$�p1�6�M���Q��8{$��G޶l�0���!���
bBq-!��R³ԋn�Ы @�Y�μ�yO��8m� �ݯ���m^���]$@VGd(0Hf�~[��B��YBOGX�!G����	ݱ�}R�L��@{����?�.���Wq��TVf��%�� *>I�an	XF�N���4���pt҂�9&����ئ��;�Eo�zn�}��<ye�J��;b�Z�IZJ/�D'KpKk1�l���@������Q�&�[�	r>���ZǬ9
���IF[N{�����ʄ�[3Q�z0R�f�0n� ��>Dq�Ц|>~��4���7�	V��,
���MK�P�-���]��p�2|;��Bs�Үφ����l	�E����>?����1��p)�5�c�T��(z\�2����kA�}�{@t�F��TË��d�H�~��	Y�n����f���Z���8�5=)Dq{��/4eۖ�P���a�<>��ڤ-�A�����-6�΅0b�(��)�C�g�3�����u?/xܺD����7is�sz�����+k{)n9����xAګf֣�pV�YE�u-~����n�W�A�P��g�D5��{�P���^ǉu�.�g��b�����ͦ��3U�͑p �OMlĴ�"���c���&M�W��,UZ����ɵ�:䎗;�}�[��82.lf�d@t�L���(z��-��:;y�a���|E8�}K���y�I&��)Ņ4}ҶD (�����|��"�I;?��*nu'/�W��,�����$�9_���-�{�Z�a�Jo�p�������H�`n����<�
��p%�X��եj��1M*>tR2c'��[�⇊`�P��2[���ߧ�ߠ$k��bFht1+�ȼ��C��׬��ҧ*�X�����Q�G�K��3�_f�i.
3�X���e_!Ḡ��&�4���;_/���ψz��
&�pS�k�_7��W�p�t�}�-Q(��%M�T���]���X0Z�e��i�N�6\��+:�v[���ɸ\;��*o��v���U�G��k�_�R��,+�����2�~#a�N�o��쓊@�M�nӧ�"���ϼNBd^Z4֩}�5(Pe�Y���U�z�@��~�n��n=룦ɻ�*Oi/������>�zƣϫ�P���5���kۗ��A	B������#�rk�CH0��~��5����(�EZ���,��'�&4@��H�cV{
yu�ު*��F���D(%�Y}@��3�4�F�z����Cm'`/�Z�Dj��K��fB��*��@�a�:	�K� �4����Z�.�\�o�6��8�*D:��7lb��eC�/�n���F<��&�\��|�9�_�i�� !@aAh�T�*Ճ;|҇�C��ew�|����]E�sw9�)��©��r�Р�p��9�;g�!,�i�����6Q�q9�s�Nj4�Mx�	-��R������(%��S��@ļ'�����j%nK1��$��5]�`� r �/I@뼢2C����J��Ҿ��Xƴ���zґ���:m�>98��>=c� �qz��'��1F�JzVb���z�'�r�X>o����vX���*6�S��%Bp���<���	+Fe}\J��]%����[ox��1�$��:t��\�i�m��ް����ix5!�&�7�C�"��Z	i��e�2�k�d��ώ����n�
'�l3ե��/�)�񧨻��Q��ADn��)���w�f� Aі� ��ʹ���O�qff֪����β}�gf̮�E!��[|'��S��h<��Y �k'���*���-�{-� K��:3�=7tC���i�#�����tbq-�� Z�i��?�c�U�������Ǧ� d�Ƭeq�ض4"s�{,������P��ň�l��ˎ�7G1�[��e_��m�&�Ș�Ӿ$�X�|`p���}"��`�.��L\�R�1���&n�BX@QJ�{�s���޵6��;M�K��Z�Whoz�YP�F�W���;,F