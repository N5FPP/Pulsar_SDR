��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>b��z�P�͕�[���O���,����9��SF�ĪZ{��A�jb�$�5!��^���4�G�hJq=`��@E��G�В�Al�E�Q�
E���'E����8�j.�V�*�.�Ҋ[�6K�Z��5�Ιjγ*�P7ۮf�������������n��J\�Lt�4�R|�{�P��������~�Lߦ6���)�9�L��
8�Fe��a0(![��0��M",T>i`�͙I�nz�rr��_�v7�.x��û��D,
�C��Y�j �'�lB���e�_���̪[ԛ���)e#��V�&� 5ǖ���y��`��v�%y&D�X"��(����1ثDgc%b�ۡN���k5��`�^8��S&kp�o�yO��N��$HW�!��M��Zr5p��<u�3̂heP:n����Д #�Ljk#�~z'�G���ʂ�]��VS��(3�ྂn<�/����,�t��̙S���$��
�������ej_���wc��6;o�%�
�MՔ�?,��KS�AW����T��a��"��X+���'۞)�D��<����mM��774ТMAͱ����`�i1g��FSS�1.�XU�W=Mꩭ}V��'g3����6k��-�|�/"Uc6���Z<�� �H�OE�A)UI��1��pd�{��9�����-���x�kI(�Ek������G#\9��5�	|�����J��)���X�G|6H��/�.@E����J��<FRkp�e�������c�����H�W�~B���)���p�
�s����Q�ƜȽ�h�{�uו��N>����Ϝ����P}0g>)Bqsc{J9�����p򘥀k^�ߡ�!]l=��L�ך>��S?ٺ����Y��~W��bT����i쏼�p;!:�d��%P�_�r,���s�ȗx�8��|�K���<!����x�
����=(n���DNx�GA&�p�Y�^$��ie��z�i��\]E���ߦpټ����P���ϒǢ��~̇��Y�D���L�l�Є*�"��5;/�������p6�hJ�y�r�W9�ZD�Ssĭ���dw0Ơφn��C��E�V�6�\�6q��Nڱ�PR|��5z��gQ�{��~n!!�aN7��zI����zD�t�#Q��R3����(jYֹ�n��Ӆ���*�å�R�0��ς�vk�D��!����녡g �f�Ydx���z�>6�"���4�5�!4���Mr򦶒�#ϭξ�E�vº�KY����wA�k�psצz�.Vx�;كy^;jZV�i�p��E���������7���P"�-�߷yׂ����gL��Ċ�3��Ue�Z�G�4�M�k�g�@B�F�[�E9��>�J��R�6a�@[9�ˢښ����K�� �3-)dߐ��Ӄ��#�瀴-n����VxNͨ1{e��#
�8��[$��,"��,��0`��G�ei�琏�&Fӎw�l
y����k%'j@W$�O�Co�F����\��[c?���u�C!�����j�o�IyWWY�}��������q��,�������HΛ;��_�X����O-����.���I@��L�����m�5�0�/��>��˟`\����УB9)�Q3	�Tu�#"�-���u䆁V�t�#���S�uw���CO�N\��V���k#b�vSs�1���E���^�e��]"Lv75.�{����\(<��wy+��=j�J�nې�MJL:|F̥0�F	{v����ǩ{9~���4J"A���o��}1��Ê�5Hgt�A�V}�9I#>���2�#�<ޛuZ��ɯ�24�"�;�"�E��n��?���Ы�Z�Ҕ弆�G�t�~���h��$g��7o
4�sN#�@�y�L��m�j��̆; .�6����ĥ�;m� W5FYpQmp��f�(�;�{�F�X��S�u�hI��+$����2{ߩ��pMe�QE�o�;�䆺tc>Q6�T�S=�����E\nWxՌ��<��Rt�1�X�Q��+4ץ�E.ݛa�&�7���
u_���V���_��A�j������4n�N�[J�˴Ol#n��:�箏r��L߮	���wxR�I{�naQz3Ö��a��K��"��ZW54#i���?	�"ʜ03F��z}	qD �ݻ޷6�0�sL���h�����Q&Pf����#		>��s��\=qi���P���������ޠ8����V�9%���2�W��D6�\7�E����D5���2Nt�$5�/T���s/'������S����h��Ys�D�&� ���#Q���8�(�c�����A�;�ȝ����8Py�;��ͯ�ϑ�%�F+Zd�����D�]�������4%�&���.)��C����{
#-��,z�y�]϶}�~V�?�
�	�#}.P�8���Gό�&��i�gI����RuT�r>v��I@$�D8�W��� ���P*�qcv'�]���q$��˻>�������vk�fI.�m �M��%o�V�4�Ϳ�|ܯ�\G����dĪ���2�wQn�e�C��$T~ȗh]�1gR�I)�)j��p�l:�b�l!��l0����n�\F���낃j����W�rv�G�\]]{7�ay?����MĦ��.�v�-Yܖ�GRx!�/u��Bd= ��:�	W�����-��t[`����5,��03�uaf�	 �g��C{UP���ϳ���dk�U ,"i�*�b5�)�8��2k�H�Q�NDp9#<p�6��È'�i4��7�����(K�'�İ�Iq��ʕ���8�-� q	�j��4(���G��k�`�J�I�ɦ�`�q�+7�PA|�&���m�5 �5�	�g���;)U��=i�U�����S�	��4=$�3��T��\�����x��{a#7�"��!���Jrzː�>�ԥ�	�3�N7B�:���$��v(+h�¼����?;�7�<�	$	�Z��������$��,���f	jxz��T��q|���UU�XbO(��!�I�Ѧ�_���Cm���}�ʌP��2���(l�S�(��2�2;S_|�Kd��NvIV>:E����m�����17gU_i��MJ�5���`5~6P�1��ՠ֨x�+<�����@�դ��d�5��=ܘ�g��Jh#bt�����vAPh�W�9��7,�4����>�<�Kl�@~
���J��&���q���C���J��-F�eu�a�Y �5
ۃ��Z�۞}�6{�T�C��"u{ے< 7�_W}
n%F�!U��V��2w->I��B�cK
;ۑ2`�Y �[���y����k���!��D��{���$�?��ch�շ����Z����\{xLj��?��
m��$�'����9*���x��Ui��U7�����0)v�ϡ׼�{�u8�G;��uRj1���*��K�e�~;&�mM%CP.���_d��,��	|0q�ۄ$����ߛ�5'�o�ҟِ�@��t�����Eռg�Q%R���s�\q���x��]X�=b����Y�����Ȯx;E�<�U4�@8��S �<��� �/�7��PW�\�_�"��jf��cX��[l��	JhG���vZ^���Kw�U�HV�VǞ�����gk�������&3|��K�6}�h�m��4�`�>1��o�O�Z�9�'�A��YS��9iT�
&�~�$>?�I$˞�5Q��Eϔ��yȽ�\��W��̐�蜊:�t9���ϐ�D�o||-����#�0�bo�|�A1k^nn�F ;�.�?TP�|�J�׹5�'�0g�*4� ��,z���+u��R��j7pv���N9u��&ي`? $���=���PB19���vUd����~�6�Ȝ����4Z 7�� �[���)n�S7e8��YX����?A����/){ƚn�L,�@�����b?D^�.��rnifi����(&�9VԶ�̍׿�ت����e�� 8#��@��(�ĨP�c��v�dc���D��������I�t��K��p�R��7��?�7�d���%
�
9�EM����3�xoM<Gm���ƟK��	�nv*��S��_��D��`�j�׊d�� ��w�p�JT��
�U��F�2Э���Ұb7Ŕx�<D���W���R�����D䪛\����㝕*9��k�X���1�f�6R��`'��Vd'a��w���0�4��S\JF~����U�	��a��1��q3�o� մ$�:�Dа�_��n��)pE��!3]-��bʰ݁/����(�yוY�`�L#Z�����^yg�6;�u�I��f���?]/0%7����LY�*�֭;7�;}p@��O�F!,���U�D��,��W�C��R(�PiB�v�9%���Ù�@��Z��~q䚿�0�/�p�=/)�a�����68�2:�a�K���5��֣�1�5��j��s���@�s�q�-7���ֻ�UN�嘝��� �a|����r���e�&86�?����j��rU��<�A(���sVT��W�p�*j3� ͹y �:Y-�X]t�1F��"�ʸ���{dRmx{g$i,�^s��z$�k!8��5�7ɥ%%��w/K��
�h/P�/�鷸��߾�x0��d� �8�MH������9�UG��tN4S=�ɼQYqV�e{ʒ�{s���m�T��э��
\�&&ȏ�_��?a��p8�B�~��FF'wKGK�(��NqcO^!�@�PQ׊TB���gݍ�W�x�K���J4������)�ά�9�:�Y�W�y�'��7�݄�������'�(o�;*�,�����! �קR����&ԇ%b8���U���)���I��`Z� �!GE�J��S+"�/�V�t�ܺ
y*�"~)@6�����g�/ʺ�����ad;s6��Z+l���N��O�A�e�A�B���'��&��p؁�s
�%�d�������2�:)t�pR2C
.�T)P<�M��}��8�D^tj�+���Be�.�o.'�_����I�-<����8M$�w�w�>1�n�0Ӑ�  |�+�`AW��|`�.�T���ac|ҫ�JE-L9�*��)͞�*`:"�,�ר'��.�ڊȦ��+@�"�ӻM>a�5	V��$�c �G�#��=�(�ٳ�!\pB�{�
׺�ީzUx<���������,;�hx��,/
ܘ�V�ɦjʮ�W���	��'����	!�4�);�w$���W"6n�����/O\���H��>/��u�#MK�|f��.�td����׷�⿣�	,+���ĝY��8&�6��?rF��(�\a�G�������R?����͝8�5�� ��(��Y4Co�w�V����	�"�oq��ڔ���=�P[���[/���7J�w�-j�ca��Q[Sa�^�䳥��V32��fAI��U:�7�![�W��)Y�xFL�Lbl�x��~8Ź&3���'��ҭ8nu2O#Uǭc"�l����� J�qF�%?{����2S�{���E��>o�7�@�ӈٗ<�R�$�fs��a����Ud����c�����Y٬J>ʥ��)���ZK^呐�=Ͷ�M�5͙
�y%���}ԉ��SmR���ɪ��@^p�x%��
��,�qdP�
�-]��������}��`^0%���(+����x�m�c7[U�nww�5�8�w���6+���י
�!���>T�r�ͤ�z�	.��Ll������j!D�<�x!S��ȱ���K}�0��2[k��pϸ��&�a�2=�%횵���U>$���Nm�+���`�ܡvʦxJ��w��b�\u2Ye�h� ����w\����wC1����B)Q�wV�G���dֵNuAP��z	b��tѣt�x��ٚ�L��ʀ�Q)�/˭0��KY,���?��LuX��y�~ST����PN��}�xF����az�aw��R;�3%*x����]��ř�v(�j��8{�\���=��0����x#}� -����U|v�攸#@v�5�SZpe�~k�h��f�k^Ƅφ,��P�I���.��^,��܆�#�����1�& kɪ��2�����KA|�_�.9�)˿��|��s��q�X�sk��e.��H��+�_]�H�ג]ؒ�0�_��[#� ��.>���q@�hgq����|���l+��_`����>`sd#����F���T&!��Tמ�]S�S�U��޵t!�o�}�H'r��2T��w�XQ2+:Ͼ�:�͍���>P����S��Z�kSP��\���u�b�":�:�64* �◳�*>���|�:6�u!��!���CL����