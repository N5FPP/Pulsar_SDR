��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��e�ik3�������w$����g|��J^]���i<�����Լ�C��U��*�yh�'ؙ�-椂s&9�
����ů2�v7��?��+��nx�	���L ��є�'�H�84<c9N�z��M����#���yA'������Z��\�����ʫ��j�A�=mr3��(�<8%*��‼�`��z�
;/w�x���e.ʴJ,�!F����_{���=p���Ҁ-S��c"�+ڭ���v<l�@�`����˅m@<�jݞ��P�p�/��Cj5�w�D�t_Cs���A'>Wr�^��K�}����&��={��=-G��b�/�,;�fX)i�}�x���&��O#�	_8]7��.Q�JӺ���P��9x�BL������7�'YV���%~����LVK��^ӝ�=\��'�����d����'$4q�u�h�?ys�m��2X��U�،�h{��IVR]܍۝�i������l�N7m\	�_�X0JV�aX�Q�Z'H�C�]���h����B��5	Sna?�=?x�U%�W$?�F�k:��OT@Q�+�a�3�p�:��A�0���7]v܅��O;y�	Nͣ��.��03��)fp�8��c;��-�.���I��;��6^�N��PM�hu��0�YV�`!~�d�0��L�o�� o�9�������Ϙ��;E��i�:,�G�O}��� ��
�NZ�`s�4\_� ��h�f��=&�*>�ZqP�7��p�=%����ͭ��#m][-=|��j��z�QUMO���@�݂+n���9a�"��9
�M��Haf�/�Y�k�" �����vP<��S`������VR������UOH���us�<T.�C��R����0?���/�F$W���W1hS��(͡�CQ�v�S¦����&+爞�f��6���·��Lw��nLy'�S��0����w{�ʪ����&�y�o�ԑΑ�`gc!˧W���&�xR�o�Д����#��Կ��c���>��!��fB��xl'�Bu�	��7�m�@�ZG�����k��V�>m&�F�7$�B%9R�Ս�+R	<�l~� ^9}PțGa`�->0g�f�۩9G�7�(�ˉ�}��4xF���_�'ah�~wR�e�O��,s��;,�	"eR��	%
���c��|W��&��߭���f��]S�/F�:�����\9g����kS3+YHiQh�N����h\����J�~��#Y�0�]�n���6�ѭP��(z��� x]�X��K�ꪝ�`�a����a6	��������dj�^�B]��+D�e:���A�Q��J=��"eH�����E}��!�&����}�)��^�_]���762�0rx���b� �P="X$�G�����GU
�>�s&W!�3�`�m,4ڔč��N��۹���W�����]��h�:�j$��w<�3FL�\ߚ����d�����c04z1s���.锹�\��V��]��� �4:-��S��:�~�qi!��z
Xŉ�驆��zP��fZ��Ƌ.={y����b#�¶t��k����7� �Հ��$�s�Sy}Ğ:�MVK���nU(b'�����t��,��{�m�{�nD%i��I1O	+'�`�h��ps��,�N?�;!��&�+�R����*�p��9��Rkкj.8�q��<���xPf��u���"�(��"��Ѐt ����!W���Tu��A>=Y͠�������W�N7��M���N�*Ta���L/��{m�c�R�Y��\4t�����`z��N��C�Xl�����.0�Zf0!efR�;�M�L]g�oX=p�Ӹ��C�IC�T7����$MEVq�"���������Qb!��J��{��'����݂1ȖB��͠�3!"�6˃����5Vz�q��P��l0rd
^:��W���	�+�N�v9tn�xJ),���2vsR ڙ{2�$&���a�r��0ji����x��2vh��+wB���/s�c�^t�0v����k9�-�iة�*m�_78�a)O�6��'�_�$W�0,-p�p!򸲱����.!%�.u3Ҽ��sN�#��$�CN�L����Q�.��Q�n�Z��B�_�c⥘(�J�g�-���%C5�J��v�+$�ۈ���	���\��i����t�dQ�̡�!1�0��JK���iQ�/[�@b78e�Y�R��3x�$
���fԑ@>L8i�o�L��a����ʹZ;/��x��
W�t���v?�_�j�yg��Cy%��d�O��Y_ԦO]a���逤�%���I��$�垙���:����O����ΰil����{-�ă'�&�$��������<Cty������}�t�'1g�nԐ1y��!�Ɨ�j�h�i>x@�W�^�-T�=rg���bO�?�����qu�8&m�7�j�
��W9y/�Ρ��-䆖W����q^2qxJ����:m����91��ʭ<N5U���X������*z����+:f����S)0֭�p-��-��ĸ�A���*�Ex၃�s�O����[ÆWǜ��^����}�2{Q����8-�μ05�Trt��6>��i�0�aI%��=���B�y]z>����
�u��Lm�v)�ՂD��/��5ں�'b_��*"_i8�H{L�+WY�:dh�����>sXd�v����k2�B�N\2��-����F�������[�A�WI
l��F3����s��JNmx��Ԥ��ͳ�X�7�9�,�yb�e�W���ׄ�=�ܹ9�1���e�w�#��?a4ﰑ%%�g�#����;?\�V��t4R�u���Q���!t�ߍ�vj,̷ݿ��=wJ�̶!,rLݒ�_ ��*Sy}V��:aR��ֹq��4}wt,�>�m�����3z�5F��g�|���c(���7L2R����nV�B�#a���L[=�a'U�d�N�ۂ/rP����"���]���z�W�~:���M+��ĽU��������T�d�qѸ!ʑ�U]�L��Ta��:B���������ym�D����A
]!�7/?�=�B�j<T��ղ��u�i�{�l�Y��.?����1U:W�����Z�Hk�1"��}n�1f笸늁�W>��͇�%c���{�A�M��. ��՟y����{��z��
��i_y+q�1��8͢?�7��A�P��]��X��|���k6�#��DW
���$��P�A�Ic����_e�;�"p ��UPjp���~��O}W����Q)޲�u�q^�+�S��P����N$��%_$��B�3��w@O;cgP�S���ri ���{o{2���#=���sIs��F�����"�3�Ǖ� R|�3%DwR��,���^V��O̶	\��~_W�����ZS��ACc#l���$���3�y~�R PW�e��HC��L$��|����Q�E�?�W�?]8�s��K����ݚ|�A)ف�Q����ˆ���w�F-揸�ҭ��
0-V��L����	����e�ٶ���q�Q!9�Ds��e�.����í�ؙ���M|5)��Jsj3V%��l����#�Ŝ�h~@v��Y;�����sٕ��}�w�� �zR���k6Q2\��!-��o?B�kC�F$|�h㛑�⚣��ƈ�$��(<�c�V�&��0OO��Qj�X WiJ���H��{��~�u���+u<Ñ�k
��&��s� y:�/j�
)T�A�?C���e�ʌZA��.�4	Z���D�L��]T���M3�M	Z	���H�0�mr���*����h-�nU�ۃ���(u�]��ا���4W'��t[���JK��"I�R��!��45s����
2h4�J��|��8�k���b��y��K��i���NF�L�B���Z7_�Q�88gv�S�s�
���@*�n�9���Y'�����2��M�H5�I=I)�ϱ����N!�M0@uF�ER���俿�ث]�8�2�Gڹ�x����Y{�g���p�$7��MU�%i�	.�:�J�	�o1��/0w�+���OoX�����Z���tL��2�*�����x�Z)�
P����)�����d#��:��(����8k��B�v�� �������N��Bi�gb���[l��g�ŪI�ؼM7TW8�y~X�R�",-�jLb�(��af��>�7�vz[A����l&-	#�@��А����%Ϭ�(	ח�;R ����~���F���$P�+ƣoK�n��Qaw�7�39�J�ĭ*�.J�z�u^��,b���@��` o~\/�Z��� {.N���\�e�M� ���}����06���#�[b� 0�U�����.�y���{�F���
��''�������vW�i{��5O9��9[Зw��b����'����䭪D8��/"!F�oӜ;��=��v��]fІ�M��M��~��[(��6�a��\ġ{��5|��v��I�L�*j����&�3�Ț���|�4���=��᝕`�]��2+��
���"�uQ��L����j 0q쿐.%���|�d0�O΃!y&
 �R����p11[*���*.ݮ
y�]?@�,l�?�=b�B�1�~,H�VWJ_�j���XY̰�g���(�筹z�j-�2Q�kyX@U���?k�1����o�M��`�7�m�b����l%�gig �7I�V��#�E	8�@�1(�߾q��XC(���ނd�C��n���� ��������,�*?.M��������Kǝ1T��Y8��#��i������g=�y����5B�)����6l�L�W�C�١�W�_d���J���Bz�P�����92,�z#�D�3z��Hb=��Iٓ�}(�K�l�, )�w��,P7-� z��n�ޒ�-�~�����;V�4a�x�oq�z�=U�HiP[��CO��^��s�y�m�?%��$��.n#lK��[$1�|\D1�`�;vj�v��6.<Ƌ��t�Z��#��V�ą�楨'��D:���v�K}C�]6��4r�K����\�O'�l��ٞ�I��jW��B����"��[-q?~�U j����dNr�}��v5H~�1���`L��[&R�P��:�7I�m_����z|T�'w%�|���͓v <ϰ;���!O��N��'5�1�OG��$�"��^�܅�F�(���l�X7���˹J��[��s�u^�����,��-����7���By�h�xV���q|��+}�*!P�sq�d������PC��	�����nX/�V�k+��{r�,��xF�_�� ���F^�B�|��f��)��,���`ne�ib�pM�(����Q��yK}�v�2,A����)ґ���ZO����;�`<�Չ	+� ߨ�5��RX�k��0�nH��%SE4*&�2���n�Dhz���8l�T�sE�y���"� LQN���(#��6�p�{Lڢe�iD
�4��,�ɩ�3�X�E�:�4û.J�|Y��b��8P�)�>�*��-;Qw�+v��kc��	r>�v���k���Z��*�w�w�;���
�u޿� ����̷�`�
�ޠC1�b6�}3�
�H�O�.�?_��X&3��m8�L��Uy���\+�1�8�d�ߛ�k��h�|�v �+~t�����}�'�|�o����>������'���2�b��cD9�
~���	@'R��Ѧ�쿈$<��N���u�gn��.�yq�2E�|�!ruzX������M��[R� ~*��`��Y%�`���a�|C��Q����Ct�wS"�5E."5�b,�b����o0
���yI5Y����En�-�9B���!�'��v�m!Bk���p�<mGp�:�i������F ���+u��;���$F��_O�	:3�����Pԋ>�'$�2�;7q��7ԇ5����̕ɩ� ���/a{T�	���,lm<۱�g���E���� ���ȸΗ�4~�i:\|l�	?P}ҿ>f�,���њMQW����6ŹR�����y�:����*M
;>g�&c�Bߦ�n}�N���^�����Dz$:) h�^]�����kb�,����b�+"���v�hK�L7��uEد��批�d�� �k�E|��;��HEu��h��]�:s*#��ƓK=?Zn���)�˘�֤���<���8i_����
�-��֍�hèU ��y�&�B��7LD_F^�0(�5����}C�&���.$��w�3k/\��A��M��5랗0�B��`5@��@9�x��e�>��%[�J�^{�B]� 
|?�	\��ŘH�"� kw�Sal�&5z�ޠ���*Z�H��d-Q�lq?0�m�$���]^C��&t���fյ';�_�n�	U��FR�t��V��Oc�^��JB�4��E�C/!��;���Z��]Ԍ*ٓ��;�O��M��[o��8,@"�w8<i���Cv1%rΗD��?�*�1�0�
��)�c�����ꄏ9ZE�Z�@�>Ơ���鬜�BQD���P6J�U�ʻ��F����*�|-��ٸ�!/3P�=aV�D�|	,=ceW�v�M"!��lX<�������3���푞�L�qaj$�YxFX�	����9�U�R�
��`�����)�ld\B���/���i^y>��r�X�[Zecbޥ�n���/u���/g���+��}�0�W�}�M`���ME�D���Cd�t�hIq�&���/���
U��&�H��pԿ��)��g��H�,�-ۖ}d�^�P����^�M���ǃ���:<z�Ģ�n7O�{�2�M��y�����nsg���&Pq#�,�8U+���k�ܗ�MtK��!��fW�}�a����D���v���hdw��5ϧz��5ӹ�J�P�r��h����wp�*���nW@`�����v}t4x���\��";ܠs �G݈�nK Z���$#'
3��F��l��T�P_0�Ԥt�����k���fJ�}���Ё�˪=�
����� k���#{�A>���D;g��UD�ڃ��"�SG�P�7�r-����N���p�B��I1����oLò��)���m�qH~6��mv�����5�'��!m������V~!
*Q"G�n���PD9&"Rb���B� �(�V�M��*�,Wb�Y�B��W�9i���d.h��W�
�n�fz2ro����?Hs���)�3I�\
���8�w���DFF�_XC�0�ЈXY
�#�31A�_��E�^Y�I8��F��06%�v�<�CYs x)��5��+I�V��3�䊒��OÒ:�VG�BF0����ܧ��UwyX�t}����h-ȍ lѮ劬�jW6��#Xpe��p1&]��"�F���ϊ(}�}�贪b���ꍾ7��D��D3ILNW���Yn�}�˼���O�x���G�O@ax��쇿��<��+�8��][-RA�bPk��-����S���f5��(�$��ϔ�|��������'_z��{T_��j܂o�P�֊�5Q�8ץ��
gC�	̖�E�5���j���c� ����X�V������P��k�nS>�)6z' ��У����k����M�Ǒ ����5����$VYr������t���;��G=-��Ez������e���Vc�t�s`�������5��;���Fp��S�VM[���V@��0���)KE�����Av�t
�wk�ȏ�iɑ�_�P���M]�'Vi��0]0����&V�_�P5�fO�TNH1�'W�G4�M�f9/ސ����N��(F�|mB�QBu�*iP6Dx�	� �����u����|?�F@��M�m�q�� \*��+*k��q@	&Zy���/���"StG�V-��&0�����߯��9�B���& �"2�'�k|�4��/_�3��9���:�[�-:��z Q�J;�<�Me�\8�5��dd�p��͗J��fJ?��z� �j��X`���|�ë᏾N��o����f��h����/!��l����VG�@8m��פ�s���8�@ʈg�w�IX�����-���	�����"`�'���B���6����'�֍ '���4�w՜�
+ARL?��ZV�}�p�n!5�^���Y����<.�E4w�4'[�UC�r��뼿n <�CK���R��1�,
=�h���j�W���2x")!�H���*2 5v�"�J��l�1���m�u�ix�I��q�(L*��6�!\53ٗ�S`�kP9���Vt���B[�&O��Y�䨒���f#�N�q]z��,T����ڑ:�#�[���L��-����1����<�=��[?k?@ֺ�h�e��0��vG,� Ԣ>����Y�G�i�V�[5���X��B�a�c�դ .��ܑ��5��O��%9�˸:�˛2dak��g ��-����i�ho��ֳL�?~'m��s+���Z�3�䅓�б8��rݰ�G��D��*�'�ZY�;��b�6Ε`;M���v ����g��5ߣ������	}v{+�ɀ��/�F�S�%�_^�1sj%��:�U}��E�l��c�;������������Кȯ1�=.Ō�em]�M�Lz�mu��G ̰p2�i������\�{kowFO�0�sl����?dWUD�W�c���.�'�𐂛},�%��/I�~ɮ���/��8�ڪ�O2���y*�0����3����u/r��q���Rٓ�ۛ��H�����QS�}n^�^#r`��I?��nO�g�k�-���~�G��7�QB�3�Q�=�yJ��K�	��6d�Ni�C�E���~��e!�{�F�2�U2��ݝ��㿮� ��(�s<��>��-ۈ�V�[;�$L�u��>��~�7���v0�֐��ֹg���3�9�E��w��VG}���e������a�5nW�Wmr��OO[�5�LoyPP>`N�����k9�#�u����&�c��.@��	9���NSW����L�t((ΆnC��O�;{+>�ʒ��C%�6��Nc|���!�-*a�4��[�.>ÜI���wƴ5\1�b��U��ߧdH#&�v�],2�ך���j�T�ec� `�-VdX����.���Im��n�����Z;.���MD���욻9t��;|YD������O�u�ž^jd���֬Gd�M�k/!��Ꮧ��b"�C�}����9FJ�B�0�5Ũ�w��X���X�Ԛݻ�M�y��!!`�5�X$�&@�_~�;�@���{Z1�����qE���i
��)�s��7gt�p+��= _V��O.A��%y2U����#_*m����ʬ׀R@��kN��
4�YT�������w<�cFN���c̝���&8jg��2�}���WQ�(�~�������������Nj H��(0�5w��f���\�1���%гT+l!�f 9���͸m-�����I�n�Y^7َ�d0�l�U$- ɂέV�ei��13����������?[b�W���ͧ6bMv������W����u�$�٧pŹ��O�����O��~����ϱ/Wj4�w��E`��FR�s�.`�Wj-~��0��[4�) ���;z�	� �ɶ�B�-�(/���ε�BI������n�3x���rvn�1����	�D��ta����"��0��H����̐=1����n���f��M$�f��v#J��e����i�.?�pKF&�z�vZU�� 3"�[��<Rş��o��Z��+��s^�(u��ן���^�Y����+ǽ�>�E�����X�$gc��F�$e(�@(��ސ:>(�"ϴ�2�y�~�/S�=9�?�����\-�+�����7/W��Ǿ��(d���r�b&�k���kHFK�R�i.!�6ؙ>�#/��u�L����k#� ��l��(u�7BX�AU�/����0JJ�۵�>�c]��� �x�J��I�S��]
�v?P�ZH`z��)R�&;1MDɡ��|~^r^��O�o�Ʌ�$$�D��Qt2o�~���P�w��c���ߍ�oI�W��̑
E�I]f��C�	����J��x�Tz���sTM�,�=p�1�gb�[��7Ą�=pu�q��[�n���
��2u'���i�y��]t/o�$'����гC�+���0eY�.#��~�*Dk�q���!�n ?1Mi�yd���D�4�������7ƃb��<�@��D"��x�П�[z��g�I0s�yƘ���q]����S����rΫ���D�O�]N2(s1�*B�a�=�OjS9D2�qg«L��dF�߰��� "M^#���+�l�j�����w�bϺ�y-��Uз2��Y�:g�rg�}g)��Y�7����U칫|����@��lOuh9��6�Ӳo �s����i;�ô�`q�j�F�Y�EXfm2��#D��,eg@��n',�����X����]#�)��:� �yE�Q7K(F�Wو��.�mz|׋-H����V�iS(�_��l�R��~�i'�&?ݖ��jaၫ��x���N��џ����w����a
�#o�Em�(h�*�j=�#Pf<m�K�u✢"�1Qx^��X�9�C[��P<�1(p-�� �Z&4�@;�Hk��Js�Q�Z%E�B,�RW�\�}���=���=ͬ=� �н����}��s
-u����o���s#nVNg��@Byۏ�u���]F��t�^PD�j�<�jr��1%���1��g���6�%��f���k���'��E���S"/%2���W˼���r�r���q�5���8�k~�Z�_[�"� 䌗Fc����J �D`���64E�N��?�F��A�ѱ$B��w8�0�R�K���v%��Rܲӏ�/R��c%W�LМ�m4H�9�J��/��2-th�>٢v�+Vu�,5�M0F6(;��ˮ8��[ �K�9�$��mTO��y��ۉ1#���"�����xK�X���Ĉf.���i[�R_:wf�;�PЕ�v�8(�`f&��y\^G����pp���M�I��b�����hıT~;��A�'�� '>���?r+���%7Š�=R�+�tm�� �<�DFɬ�`-AW�"����Fu-�wI��Y ��E��ߠ���8�-->�@0��P��5S�)m��~~ܫ%��a������X�v�M��j!w('F��`�ISD��cmUOL+�2��_�bQ�|�����]J����j⫤�2Ԫ��ͳ�*;���B��6#�{�����K��DQ)���c�-���
4��<?�6�8�w���X�C+��ڏ��c��`8��̷۬*�6Y�E�؇!Eq��x����@&�V�d���p��G�G��H�����o�$�/jL�M� P���p����t��~��L
��N���X{�O����Ln��G,�/%��v[&�f��%�����D�9~���z�fi^��%_���3¨��l�0����8N	tXM�))GT^�=Խb�<�e��Ȼ���Gۻ�ŪԶ	c�)�T���ǉ�e;�M�?A�]$a�╡��1��p;(5�{K��E��J�7L�1���>!Jqp-9�Y8�F�P�xou��Ў	�?�ky�x'���U_S�^��d�+%^eM�O[��g7���y)c����tR�@��o���һ�|�k+c0 �D�D��}���R��t��m�|��F��i4����tq�[�i�@P]MG����S��QR�~��� �l�}��'�%gXU�G��5{�DE!�l�4L�H���x;\�0�}J:��ׅ������4d��,$ef�N#-H�֝d!��[a���YT�||�AUD	2B�ހ�#x�$�7@���eZ��/;b��lqx@����)p��P-���9#��/��:��Tq$)�Un)��S/����/I�0��&_!��@
S�U���X�)4_�uU~����~YS�m�/���c`�"��yr~��3%�f���Hk&"[W�ofbL��F�c1�DRA�%����da���R{8�5�ݎ�du�)�M9��r�vp'+5���E֟�p��lb��1�8D.W�eDl�SOH˝h�� �L���GN�i�x��̮=)t�. ��[J��vK ݅�T01�Z��Q�Œ���c�չ�Z]iU?�p%9�A/��:�8=|席�-��ɀ���3^�#5��Q ���a0!���g1�����l|���W5E|������V=�@[��v���^-��p��IK$�n3z�c�R1i�Ӆ����_�zw�т���s�!��6�V��Z
��\x���n����u�°pM]�
[[w��1��U�x��&�E�"KzJ�P@�#M�7�w��PR;F��E�`ȂC��u��˷d���#��ޫq�!��1��YQVڐ����H���w1'��b�Gת�n�EUS��:Hc!(��L�#�̋�칧�(����YQ�~�jypV也C_�Bi�9�Kdf#�]|7,�x�qW3�a-%ˍ�ja�(�f��2*���+��;kiџ�	��j���lx����Tx�c���ͮa�d�3�d��U,
du 
5,�"ŉ�5ޗ�ϵ�+��m�����c(Xe�	��#Ȝ��PT��
l9X�ˬ" ��Sjj�1���ԪYQ�51Gk�t@sc�8����l�xA%ҝ����<�Y����-zp���<&4��p)��bV�/0؍x�I��զ�I�gWM�N�C]�f��>�Ǔ�UT<�ڿ E�cX(r��|	[E�y�2�����ί��U�i�tz��L���.[�=H��e���sKK�6���.c@�"'ug��8M'�� �;Ԟ���x�T+�Bm���M����؈T���4i ���(���̓���
���������qn���� �*)>��Z'"�̣��of܌Yϭ0��Zxl�%w-���I5`�����nF􁽝E��=u04��c��i���V����죦iI��k��u+��y�@��1H>������@�н}��U|�Tkf�^�|��-J��s���\!~�/��^@W��|C���eѰ�r;��D�/���u0������[ <ck#9�k��Y�����H�
�
����y�	G�W�f��F$&ɡ�\}�c�Mm. ̒e/��ӊHWI~$�A��p��DR=4�
��W�r�3�0�q��$�Z���)��	���@��d�;C�E��=�/���u!�q��#�Շ�(�  �&v7���o�i��4��NE��607�	�v��p� ){�W�ӒI�NI��@
G7׋4KC�9$Ѵ�{�pEؚ�$e�kb�|g	��V�d�76{�A��8�x&��7!��dl$`��x�V�M$���$J�k��Kp.{���G�
�Mu	�?R���R##e����W}�,�2�"{s�ӑ��s%-�U�:�$���˵Y�)'-���>{>�t����ɜ��F�5���f�˱����
��2�X��b�88T�;�d�?)ؽ#�d[Cp�c��N��6ģg�k�v�jv��jqV��.LLD
=к��Z���ʹ,N?ɹ�� MP��fSG�<z�� X��U�#�}��!�lq�<�
e⤔a@.+���.�W�j)M���
��/c�wM�s�J%� �ʀ~��tv͡�1'A��9��ܦX` LU�EFp����Je����;<MQs�n=ow����^���H6QǎnN�("�_Q��ل�~�q�ɌOH�l�̋��N�?D,�iN�rf��͍��N�y�\�s����&������-�!D��E�p�acƲ_�i^�NI�Z7�S̨�E��h'��d��3���
*2Òe�UH�8��������Qc�#��c�"�,>@r�B��<bw��g�*�b���LH:���M��s�N��D~���HXn��b}g�2���mOrG�m�,�Ͻ��7뀥`���T���|��p:��G�5G��Ɗ�_��ɴ�U�Mu��X%�<?��J����H\��˃6_�w�Ht�J]D@�i�!`�͹� Y�7�VF�[ٱ�D�S�����HlY�S؂��[����)2�}P�I��DT֚�	���J7�s��������	���6Q�(%M���W]X�Y
�q', PA?_=�ҩ�e+�B�h�6"�gv��ϸw��+��������~�,,'���Ou�i1����eWMRs�i�Nj�����,�o;�4Zd���(mӔ��@��%�D=��nVk��$�j(i�h��\��:����� ��4�0��4Y�`:3�'�Ż���S���В;�^4b���q�g+E�!F�n���Tzֵ�Q�1� Eg_���,��ʀF�Qԟ�J�K��,5x^~���@Dц�1s6�r��*!�4y�TΟ�7 |_��?p����F�&.��(={��Je���,�!��o�@A���^{-�%���7��'�6���IM.օ���%b'�? �Ηo�QxY����Fz��N�� c܃�7;����ϲXb��?<�d�;�K�)���t�� �nf�����	4e����=�!u�S�.ת���������b�P"aˠh��%�r���6 N�%����7m����#Z~�R?�H�P���%��m �0���i� #9J�P����)�rx+����4������G�Y�SG�˦��u��C��F>������v�fn��7Ó�� �\��_�=��HL d�)�<�Ȋ5��'��4i->�)�αC���B&�}ָ�s��t���2�=�	�!�l� �|g���v��H�YMe�TJ	���� ַ�PȾA`e��O��]8�E�ɷ0����x�$�`X�9���V�����/�3���v%7����Fm-|J��E��S�c��'�e��v`\8˪�2vn�=�K8��륈5t��\�bȌ�Ę�q��&Zƞ�Ql�ʣ�'�<ȥN8^��r��tkw�o�4�>�N�Ї��8�]��ܐ���@!E�������9&��Ó���D�BκU��C���̐$6*���_i���!�Y���}tG�b�S���S��jN����yg��T
QL-O�73�Y�O�5�ĥ1V��1!iԭ���|.s�9�!^=��d�8��eUr΂V
p������#I��dU O���=���բ, �ה���7�D���B�ԯ�I V�u�mPu���ŋ����UVx!"�����:���V~E>�������h� �Kc,�p{���5�4�|�g`5A�L�RhTQQ�����z4D�i����7���HX��HI2�����>)Ay��O��n�ҼHSԈF�U�bS"���Ξ״���z.����z�E㧇�5���a�x�y�Nq�ţG%L������{�#��9���%Pq�)��=�FX]�y��8����8���`�4C�8�q�����n�_���t�tm�ly��+g�E�?=C s��"�g��
"��3ͺ/�ꄶ����������Z�mr1�T���^h�+�[!6/I#h_<��"�n��A��C�$�������J}'
�6x)��veh�j�;��'�o<u*o�t��GSUK!_�S��S%g�y'ے����?����ZqoӼD���D���}��̓�k`�ց{1x� ^�c�1yN��8V� ��h��3��J�V��d
�zM��!�*]q�n�L�Rm���� ����5��rB;\�J��D���SP���1;�!�HS�ʩ�7m��_/S-'�E5���� _/�$�]Ṉ���\�Ԕ ����_�>!&y҇K~���b^�����sr��*��i��Q�%G�<�49���9%5�64yR}G��c��,��:���6�Ža��ޠ�J��Cg�!���z�6-�L5�!?���h������Ƅ<�o��zE�q�W(�.c��-g(����-i�g��$��f��/M]kq<~"�����Y���~\np6�-����i�(�������H&;���5i]XKߖ��W$���}�������c�õ�y��-W��_L~�W,g�G)�c�~�SJ}X)����1V�R�� ֦NUJ"�ݢE̮����M���B@\R0~���@����)u������0�e�P���,�F�1�����&��c	0tO�;�K�*�������*�:A������F�[��XA��Ƃ䒿ARTs-f��Q]\ច��9$��ȿ��L�����d�-���k嘂P�d�a�K	�(��uTA%K��r��zu!�Z�v`U ���S7_4C.y*!z�ݜ���+��(�{)��n�`C�-���]���~֣�z��s�K�4�M��$
�I3Op��Hb$ېb�fK�D{��ȱ!J�"�@0��z�u�;QK3�H��Z\t`&+yfZX��w��¤�!��;�GM3���F!�Ҭ�;���'kǠ�I��+�;��M\]�-s��#�xZK*:�q��.�讂���b���|/�~̜E��6�,ޚʺ����{��~ؗ�}M�T�HxvO��]~T4Y���@>"�V�|X�do��T���&�
���Da�a�N�b���hP9GT�qDIO�xcg%�,D���-�_G_n)��S^�㭰�mY��f'������V��ڱZR�ѾM��h�0I�S��,��<:!'�hO�c���`�  #���^:�<���[6MB�:��� b���%��h"�%�%�1(F $37���D���w{'�8t��A3�� �\���R%�#��M�������'�Dq|�*/*�s���A�|z+IA%v�{�h�yY�y�����la̫>t����{�:�YY��N�������l�g�-��OS��ܨ���QzDOù�5�䴈�;P�aڌ�h;�W�+�yԹ�e\�Y,���K8�Ma���z�h���]������47q�������q$`��>-�2������F=�������o��/^r�%a�߁0�]��56*�:�m�;�p[*�m�"m�{����K�?�j���ew�W4�vg�۴%���rr�����$�H�5��	�"�8û��˪d�ò��e����x�@��uD�E�@a����&���B��ɫ5��������a�?�cD��q����CpP�J�rx=ѣd����J��Ù�!���;��v��S6j}J�?�oN)Y�L�eJ�����c:�A仾�5l��*�҆m�f������s�H�D�y�#�t��g),j�:I�z�l&R��$�èc>��1R�M�Ύ��Z���Ϋ�_�#pӥ�(�v-�k4cV��EcE�y�U ����	�Yv���6R����ߍ}S�����
����*�6�N )yV���3g�"O������b�]u��H�<�2�-f�����,B5���a��{������wA�F�w{��!PWE�D����(V��\lV��
M��2�s�8}\ԉl'��
��2w��Z�{�Z�t0WW��"k�4�9��� k�L��`�F�˨!�
#�i����.4�m�]v�u��N�����W^�2;���zM�Cs��n�s�C���A�tn������u�����+�჌�PC�{:!��&�Q{.�Q��{�,�K2��/tN�����1�����%go�$�P(<\��*�Ӕ��v[E���g_����(��_j�Zڼ�y&�g.�~��I�Kv��M��;��c%��-U�Hz�/���?��W$P�/�: ��\l�y��6�E0��:����ۢ�lY���]R1�?$���b����0桂t��,��3����)�J����Oq��t��N�`RA<��������T�7����f�T���� ���`��J��_��)��A ����V@"|���u4'�2�e~�?B�W���d���׫��!ϛ%��U��*B���l�m�/%���r��ݲ�<è����ۘ<.�Q�E���qs@�u�k�C
�)�a�n���A����!'V�eRz'dҗ��Y��(�N�.8tƆ�{�HK|�sRbޢ�P��d��_O�p�CCI��TL?��z��oy���f��uʍǖ�Ƚ���S�B�X��8Z�_�3R	�.#8c��&�4���钝-�R�n"�P���OGb����Y�=�zC#�����V�h��4��b��+/J��=@�'��w���UMX����^���' �����Ϻ���?@��L�؄��r�� �����:ԟ�Ų߶�q�Y��@�m���an|�6�<��>VKP2`�d���B"(����i���*} �*Zkxn�a�ډZ�������E�`��Uy����w^��?.Ԍ�WP7rJ)1�/�&�.��0hR#-��E���g~ZƔ��nh��L],�f����	�Hŷ��R��y :�p���b=���Bp��)��S9Γ#qK�Ԅ�EP�&�q�`�M�s�qx�'f�Tt�����M��[����9�k���Q_���!���/�`3/Z�ż����>H��K��Q1}5;������|E�2�S9,- S��2�L+:�=��ZL�귚\F��cU<�uE2�D^A9b)C�qUx���O{O�mU����@4|��Ҩ͟��Y�%��[#ЗRT����7�	"�%oGh?¢{��FE3�#4���8ͨ�Ń��qZ>sj�(�X8��qlJ��΋�]�=��E�?����d�
U���6��b�R�Nꀾ�l{�Z洲�����w�	��)��0e[�"��?��I �l|�1'��{wI���<u�'�!��5ֈ�f��N0#���2'0c��:ʚ�����8bz&��/<���@��)G�;��Qcr���&�2�i�a�e�Ts�@|?��aq��oB�\Y���x����ى��&(���{�˒e�\���� ��ǦF��iyg�=�s�&�&��1�Ꝩ�\�9����FV�I��%��i��p���E��:c�S�;����Ѯ�\�����j�gM��vV�jM>qO��!Pt�'�ց�X��`�aˤ|�P�́�a�����{5��|E���FO��]������u�,�D�o3��j�D�����h8S���XgT��1�V���ASP�ɬ+/~������Tv`�6��]� ge�X �Y�I$g�M�vO�
y�U2K�( ��]��aau;�S�`���	�p��}V6�����\��_hYyB.����P�7�獅J�{��N���lE*���4�Vt�w8�;���5:4��D��Qzu����@���
k ���'�/�Q`Z��Z{DQ"�1��G
Ο�P�h�eK~U������!mOἁ�W���	kj���!���{C�NE�*'�� ��P��<qYߖ.��*e��`��Ot������ߣ�>�2�$A|�����o�CF��ܒ>�!� �w/,�?�#�=�L�S��O�o[�S*�id�3pה�hTy�_ �%ւJL͕N
��c��G�SW	o�(��TҒ#�Zm0�F� �~��Z~���:�
ho���M_�I_�
,�qBN�s4�O,�%�U�yd�����D{�&��cФ��Gp~�XZ7K�ߋz4���2��|�<�In�%�#�XZ���{r���x||ib� K=���l8��ںx:�%�$t
+"��5:ܐ٪j��"�#6�P���8-�	r����g�~>�iG�A'��]�nվ��Z��1�v��"'S��s�5/���r+�v;8��ݟ<j�.:���U88=D���DL.�tDs�^޹0΀�`�),��<��g���Q�& �`[�Q:�1'���[7)���bpIL��y��5��3x1���N��H7�Z�,(O��>��$�bM�o�s@hJ*��^�U��of_q�%`Ԋ'���&��Y ]Kei_f�����P*cS&Y��uf�w�N6��H�;�	�����f,��t��.�q,[;\Ɵ	N�+Se�2Y��^gz��c�
EMc�
�}�����T���C
\lJ���� j�}�or}�2�>@�۪��;����Z�����%���~�#W#���çr����V2{��-!�,�"f�*�ê�<P�E�5Y������9�r \h�+$6�j��Qz��]��t/�|��b-��w��n'��m���o��L�O��"���<?XZ;W��/��"����(��K���C����V
�HmO�t���644-�3��_9���#��{������`v�"�l��;}��Rř���7���R`zlH%{Y��%o�;��������.�$=�w)�;c��@� nZ�8q��㧫��!DɂZ��ιyڟ�.0��j<�š��q�P��+z�+������1G�d��0�|�^��dN��!�M�c�� ۬���TL��^��BC2�����|_���padܾ=bv���7����t�'UǇ*�G�#)��JL4oƊ�~�K���)d��b��E��w�?}��L"����:]��;�H՞����uh%��w~��58�⚨M���R���*��C�Ѥ�;%_�^���Į�3E�U��$&���j�W�֊X�J�0���z4�OǙ�CK�$J]�i��G�ݪZ=#�-*�U[�-��s�"�@7���V��"��H[�_Içou��hhJ/8�bâf���D�w�5��)�9�J����4>L�z^g�M�Kp�����ٟ<������~���̊�zb�p/`ήm�q�ݜ������Do&�{�a&*cgzQ�e6n�M,?�Į�����E���=���'2| �}8�趐"�+�(��8�p�U4����(iMl�gz{.�RN�`���G����L鱷7ec�����)�k�9�cOYV=I	)Z������p��X���FZ�0F�W��F<�����E���7˗���I�$)������P����(�wL>v����GS���!x�K1��ܠ��P��E6��%�m�>Ϛ�[�^pL����A��r��7�,#���m����^nGbʈ'��r���G�zx�]}B画�ѿ�d"=�G����\h{�z#���k#�"i(�F��wx�<6�|����DE���>[8�.�an�GP�Ԁ�`�5G'�a���dTW2�îC&	�=dQ�k8�Sniq,<{��H�b�����!��i���k-�9�
]�7�ϿQ�� Ezg���7�ݸCD����>X��A���S����(W~��
ʕ�䓼�~-�̱\��N8Cpw?��ժ�\7���-b��)����_�d���f�;�`�r9H�_ž���<�9t�ЌC7���F�X�W�����'�Ȝ����o��۷@sex���@=>Et륾�'�[p��pI�?���0�
ߨ/*�ۧ��N.�X����Tѯ��/��i��:���S� [I;�G� D�AP}1���L�9'-,���\c�ZSO�eA��Uz�m���<�l���~��J��[��+�����xg#���V�7��T�D<(`���J�9-�c[G*�:���2�l��D��~G�SG4>	��:c�J�If,�@-��kuE��a��1� �y���Q�@��+R�X�{����]�����{���Ġ�9B�T;�+�.���Mu.�,OU�?y��AԽ
��>X�!(ׁ$K��G�����>�j;�h]��^J�߆��)s��{,/L�Q��9I��k�\y{�� �˯i�1��ԩ}�FI�
���Yl��$�+:�Ķ��O�8 t��G5|��~�,�'yp���?��γh�v�!���l�j���Y�wt�ا��yB���rWX��.�,��}� 0j<�Ѣ+�7R=t7�4�;�F 8�Zz57l���[fzE^ڧ"��V[�^��m���$`6�QS�W�j�)�'NLT<���� -�q���Az�bn. � KE�����}�k��?�̣V+�M�;�<��Y�.SG&o�l���៛`?�F*K������h5�G\�s��o��0x�0��y�"���R*Q�*Ъy�?.����94�tPD�􄉸�z�V�k�[W�����1�o���� L�aںI|:�o5�b�b+_-�5L��hY���IN�d����L�L9�s���h�0I�%z����(�����vҧc��{�ק���r�2}GZ�Ap 7U_��!�bN]�pL���@A&�;���Cw���wˆ���|~%(�3�
��kV�ｺ����@����##^��}u�QQsN?�<�e�){?�>h���7�k	�������Q2����Ө6W�@9
��Q-�;J��vy傜K��Fw��B��g�V���i�}�g{z�<*�[��4Y�S��%��E�x�� ����}���4!H��Ԛ/�)6#���4�4���!:���焕���Df��� �`��/ ���5C��)T< ���m�H�v:�'�x�WL૫�B�Xy�S��Ud���Te9wmN&���w��I����8Е;Wv6�o�N� !�V���Pp���t蜏���|ww���
{C�)-W�-Zկe�}x�Q�gk�L[��a��{�2�9 �B�bH�&@/�1�����:[�.�~�%W�&�E&OY�le�<Ƅ0U�KU��ʁ4�?��@����'D�b�!� εҥ"�d��c�.�G\=u�5�B�J���&90��q��M�*b�WEli	[���"����'�8�� A�������r.�@X��>����y���5��{���4�G�n&	��>�3�=}@a��D"=���;�p�v:�qK_(][�W?��I\!dh^��I�)hƽ�B�+��`�.� �}�{U�W6�l�K	��
rNG�ӡ����rd�P55῭�v&�[LR-�!��=���|ն�~��Ȱbθ�#@bS�4,�C{D�l�Om�u�s&��t�؝����v��b\��0�R���"r����J��l�Q�f��\��f��j�5�3���t^��P��*7��9ٰ�����Z�<��]R�,�ʄ�A�����/Y�q��#O�H���9ح�:�rc�m����*�%b�|XU�P5���[!(�?b��Ż�ؗմ�i���v|&�@FI��rN#�#�^�un"j�p@nL靯�F�a#��&˗���Gi`)�?��S-e�?o4�rt���?{S"�ȯ0�x �9k�|S)[u���+8�G����=��}eQ��/���A��P����������m^��S�^g���
����u�gau'ǣA~q��c|��&�K���T��|�:�_j��b��\gԔ��mX��
�
M^?Sy�\K�vb������d��?��*JҴ#=���#����O��/@%�16�G�u	d�Vԝ���=�"Ƙ[3�X����M<��������c�x���U"�:�c���vZ3Q�p��Ţ�ca\�����r�v�����??�_��L���'e�Ɯ]��X��y�p�Q��>Vl����}��|	�^��������,N%&��B#�5yRj���ۿe-���^�� ���o�vg_0��`yp�(K��ʹ�.E��.�N�������
����u��e�h����@1��.�7-�{���'��3���@��<\4'-�P6>�1���|d�r/�F��Q�N�𓷐k���T��q0Xh}S4d�ɱq��NU&���jOsԽa &��;��y��f5��[�4W���!���Y,	�_ ��(������+���q�DZ
�Kڃ�>���Au�#k\m܂��sG5[��i�NG��b�;��/�@#�d{h
�ld�(������C6���!��O\U�EH���ҍh�.�7S��1rfC�Zj�K������G^�$r;f����]J�2��Un$B�>�_��$Q<���]���ܸ����.��u�G��}��o�MW]l��Wj�n�d�7
K`XO�<���>�f;�����|�k�k3l�T�!�a�!����C�aI�pe'�i�`�T���D�x������Dj]\
p�,������*��H�y �B�^�����Sc���ɩ�u�8���
�Iz�+�a�)e����@�D�G^���k�5�,��9�bR�[���M�)�jk��h��:��=I��� �?�
1�������f"��n���nM�h3�t��9U��J����o��,{ݐ�o��6�0���$_nd�WG�tc�)t*�Z-,s�;KԻAG\���!��#j_z޳�g�6c��<����.p:�}�l �/:�k@��++	��0��� �J� _7Ã�f��^�� �)�Y[<�,��!?�	�쭉�e���/x��[VJn�����R���(����&���p�O^�!��j���Vie7�M�D!j0j���<ũ� 
��B���g'�����=�_p���,��7j�O�yb�)}�������z8N=�̡vQW�Q(�C�M����u2�)��wɻ��EV��g�yd��jY%u𽃫'�T�ˁ�;Vea��拲�?5V���
�G�8 .���Ѵ�?���`-�������]^nVm�֭�� Nu���S h����Պ��K���vz�"7��T��~��u�䰂G�Z��,a?}�L�Q ҹ�=�ۤ�����ih٘������@ �kdݟ�C�G��W��C��A�c$���6�t}�E��+MR%�.K,���j,�D������N�Rh��M^|++����Hma�XpAtQy/�1��H�H"�%�N��E��g�e���\] �f򡵌u��}�	%]��a8��M�����C���Щޮ3�v��K������/�+�v�|hL(��&�K�IN�d�D��ܹ<\MB���Y���Oq�'�*���N�_3L �ۦN�,dEhus�n7��������()��?��� ���D�P�i![�e����Ԯ5����	��I��\����y���!E��nxd �
ѓZB���|�<�'��ƨq���4����O��96t���8TG,�aU�Y8�Od�y��������~NB�b�tkl��HHab�q��X�֯�1^�|*�j-�G[����QTM���-�T+�=L�H@~r��k��W|���(.����8����P�J���͈0kH!�[0�Y�����S���y�4ЫF��Ui�iP�	JR�.����]Q�G�$�7�����>�r�X��XC-xe-���~|.��.�V��&\�{�6��c��4V�	�Х̭S�x����`�J��I����b1!Z{��q���v�2 "�z���U��G��ð�hMJ�z�r�{6-��uMTB���0��H������Y@��*�8����&�1���W�uy�\�,��y�/�����3��+$1�X�o��G���^#',g�o�Eg��Pz�����V�`��iF��R��{��Z ��}jݮ�7�6:#��Lx�h0�G@���F��{�s�!`�e/z��V���~6�F`ӻe��-��(�]Q�U�<���K�)��Y`�rE��\�'j�d<R^���tkLz��@\Zw�}�n?v�T��9;(�w]���c��?��OP�y��%�_Y�<�����S�A�4V�b���h�Ϋ%ΎmE[�p-��C�kb�l�Vֆ��kN�fx���&g���2��g(�Z�PmUg����x=�s� N.��!�]��R�wQ�Z�>��2K�"2}���i�wc��@�e7N�YSZwܣ[B�p$Iծ�� 0��Q8��D�3^����k�����`ӥ��t	�(�*������1+���;&ҩ��@S��
WCװ��^}Y��ܺ 9k���Z΅��R�/Ej��ꖌmP�o��� ��¨uJu���[kE�Yճ��8p��7qac�i�'��wK|Nf��0�?yWnm='�FA��?眲�Gx�'�[nM.t���eZ�K�8�@�h����O��Sζ�E�8E���54��%���`0J�
��뢋��� vdgQ0��+�d�:Gmո�V��@(8�v��al�>	?&"�I�I?�O�apnԜ���χ1`P��郎M����Ds���{C��ێ�O(���՛�N�3�������C�m�����jfN�~_Ky�<ǘw���ٱ}.+��N����xI<�hF��XU�> �H�25� ?���U�>T��X�#w=��|O�F워��G�����FxB���Q�#e�� *�+�0P("Z�ǆ�V8�[5֤&+4ͭK�K�����O��x��6�	#�P�ȁfP��`�ݠ�D:����,^���ĎW� �	�.BN����j}����T�@�^��@P�*X��&	v^X�t���_�5������(%)�S��.%#�C|�z����KpF3�\扪�:���Oc1dd�FlM�	�7�t$mz�r�	w��͗FA��3���NDN�"��g��zм�oI�k�����D.�Ǵ����|�j����=h��y5�9l�gV��h|�c+�b�~'�5������"G�J�s���N]�3-����@��<�`'"���(�bzQ�{e��ك{텵v��x�u�N6>�"���#�̘a�����~���G�k�t�GU����yV�پw�ct[&�A��gK�K`�xF�2@��7O�0�d���V�W���\��@�'!�2 Z r�����;�).l������%�h0,�5W#�A �c���rf���!���5��&F+2����S� #�`Ox�ݒՒB�.����ꉘ����=��

ú��"\ێ��wǹ�m��֟x��\ /��-m�F68(X��F~ԑG��~����~4�P+��>��ՙ(xY���<���_X7�3�%s�:h6? �~��; �Z�o�"�����Z��F�EY74��s-��$vEpҩ�:��G�z]�,\!��7m�|g��ZG������x�b�Oĸ_����A�Mg^�鋮�OFz�H��Q��`��u�g)/��;���uoZ�q��u@2?B��~��O���v�g͊GP�1�;Z:�l��Ė��<^A���!��砻,�1�^��!��~�#M7P�Y�-mQt�B�G�3�n�ƾj|�e2���B�{$���/p��Sg��)�|v��p]���|��Ʌ�M	�'*=�c���������
���z-���ʍ0FS���3�F`���Ȣ����d^��/�ԟ�����<�����6��[�T4˼�cT�s/ DK�d��Q�%�lOf�0��R��턯�񲔴���<�G�+}��;�<��8go�<S���)�-����=�|����2.�R��ú�0�����ծ
W�0S���g@��^6�1&�&,�Ls'2����N#>$���F	���=���]`##��my�$N��S�<s�O衸�X m��\���˞�4�C	�k���슄:�ԕVF<z�����P&,��}dC_�]��&�������$�.x��w��c��
�/����gr��Z3b��u��������z���1�P͵�6����=��ur�̠	��v�^�9�"
b�F*9�C��X���
Rh�s���k>&��X+eS�`"��/u7ikN�T�^^�?�b��$m��e�L��=��P���s��L���ƿve�'� �2�&� ��J����ƿ| +����Q��f"P�]�S"�6��:E���R)�t];�n�mf��P���HA=lxk�@p5�%��Y�*(���C~���G4:{�e(��^�26T�n�鏏�wҸ�2[���]��H�{����=��G�69�����>%���Ы@'�GL:5���$�͙p�0��+��y��uM��@���1F�/V��B��lkQ.��I�oW���I��x��!J��6�y-66�p�Zˡ��t�>�>P^�C�`��I�Ψk���(c��j���6�é�{��?�Z�%~���tѷĬ@�c�Q���C���N*�~3�F���!����G��}����f��n�~4A�,*)�5�.ۣLB������k�zL���+ܚ]���>�#���q9)��U�Q�1�*��ӯ��҄�rm _��Q=��W8�L�M�U-@\�"��2�c��mc��E�[����QI9��_�`2m�����񥇠�1�nU���un���� �疱3��������Z}%�Qa���m���� �]�����a�܉��%�^G��fJ�{V8Yj`�3�=8�ݸV����8�����d�U��
����@��R�{t����D��ܕ?��|"�8�i�Q� ���C���{|���[gI���|��-���Kۡ[�Ǯ�}�!���1���{�轎��aGW������W�k���2߰��dע}0[��_&�h,QH���5�.���i!�e�֫y��*'��Μ�^��]�L�[��YZ��С_n7do����?�3�ڹ���Z�����X�3�ǘ�:X�~�=��L"�Vx2�/h�\z��{��#���V3�ɗŞ� [2u��̡fj�j��zXd��}�,�Ԋ1�<S1ϼ��������<�0a-҂��a�v�\D��Q!��e2y!J �9;��	�Ϯ1�ko�A�" �Y�~��d�u8��06��H�m�cI#Ґ�bB������Z��l+u�
`�^����lA_[Q4�C�=���4>[�:��Z.� jV�<�,_��U��w��̉��eLGr���R�?�~��Ǔ�ʸՆ�Kf�,�"��au<\t�U���)��|����a墲c���
����ܩp,�w�6�=�F��D�w[�L
�H4xŸޜ��u�y.��I�T>���]
?�}�@�C��AY� ���v����_��~�}Y�`��틃�iŸ"���G�p���K�:��hh�5�&y@�G��G�"�]A��R��+_V��3e�d��}�'��^��n%��e3�O�ճg�;��U@��*R�sKVD�k�Ά�~X�}<l�������Zs��j�DE�s�g�a'�,q�S���a��8��q��M��<�e�<�X4���ہ��?d�Diq��<��:�-!�LȺ	s]:K���k����F���幯�ܬcQ�
$[޲�&ݯ�¾
�)O�;jZ�i-�_#��� ��%nI�_rs��\px�a�=whɬ�ۑ5��+8)�/�.�$��״l��d�й�N�^�>qAh�oo3T��S�ic���psKi�Ol�Z$�	r�z��~� �J�e���kc�S��},��Z��/p�� �I������PKj�r��u��La�uzI*Ni��{�(7m��76�����ee�� ���>�-u�z3Z���8��Ʃ02WW6`e,TG�q����ɒL` ��M=JB���Y3qV&�rcR˼�ڌ[g�,<�����
<v�ZI�W���O��3W�'"�����Ikx�rF�+m.��{�_@���G���u�6�ܓА\u��A۶4�x�9�Λ̣K�|����+�L��*C<8ao@�#��if�O�JO`}(qZT�7 �DU������%jc���>�Nm�����������Oa�>��CK����E������Z�=M��:ͳ�-X���X`�:���6S)�pL�:�nNYy�Q�i�������~����E�a���5o�X}�~�{@��i(�F98)jJ��T� �:��-��E�z5�WL ��PX4���Ñ�������	�[\�2�����`?*:2C��멻��.�޷,�� ����Zd�ӧ���W��Ml��z��FVg�g5�3
;��%Z]�X��Q�g�:jj�QdE�a��?7C�����<V�x9k��gn>�q�Q��v��DY��u�i�,�5�#�%�8
y�7p1���/}�������/Xr.��B�}�1Ui�#�z$@����~;t#ыR��Fa�;�e(8w�R.�w��~rT���nvؚ`����~��"�(�����ȟA��k�i��J��{���Y񭕲^/�t�K7Q�ț�L�w���z�T�V;�,`�r��C����B���*��h�WU8�'�ӱ����(��?5O_�Hʷ����CP�vo��le�-�P��Di��dc�װg���c��a����oc������h�P����p��F���a�2��(@�i�C�OF�*���^�
���ܓj�%/��b�K����5�b�WM��7�����4�ί]e���hs��K��y�nH�m�]8�aqpزۿ0\�A �)�6VXq����!!.�L�w���H�^�
Ur�z�孫#OC���н��oV��-mI��M�Ol��<���?ƍGX����'Ȼw��Ϯ�T<�q4���z#_
C#��~�,ʻMU[���>LC���԰>��Gg�G���"	e��A�C�z�k`! �~jTlu��$�3��K���z� ���79������8�w}��	�y���U���Z�湨x��|t�v��9d���șaؽ�^N���L���%*�Þ>h,1Z��vİ�j�<�G�Eǥ��9(��>{�KZQ]�C���ع�X�F	9O�<y���Wh�Cd�L���H� �N�D[�3�y(�~��\QM�>'����3>)�i�A�u��Q�=Xv|��|e���O�3� ����q���Sq�С$.���`��t�?Zd��>����!��B/7��@�bN�5�r����x\D�� o1`�3��j���B\�RY�Ű��H�n���o����t�VtBM���Zd�g'�i��u�๰����e�8Nݝx�̠
��d�C��m|�<!��x�fu��tC�4��xc��ΐ����nJӏ�NT�d=i��n�>�.`��L����6N��ȹs�ߝ2uC�#�H�fI��({�`e�7	k��\j��;��z]�y}sLb�9B.8�`_&����!M�[�x��K��G�=;Ӧ!��� �牥w}�l�D7��yCf19�s�9$�s{�s4�Ko��kM�	sr��X���'�_��-cJ���|3i�l�$`%�f3�Db�W(>!l�:�h �Q�❪�ӅmQ�v!�r��=����Ǘ5VT���:%��'��&�Td����LL��;����/�9�[L�;�@���6�,zF۟�=k�����2OR]�q�-<�����!N�7��&���[��OR3>��(��5P���:d�1�;G��ߚ�6d��[ĉ'��^�S{�����J�&�3s�R��1]HG;~7Yx�GH�A�x�g�1TiZ,�;��u<�R>��i��O˗(q�4,Z&�s��I�]'���Zb�#$�5�CDp꼴"�����H��0�>_����2�O�#*�8�)�2`�#A��s,睟Ϊ��_��% U1��SJ��|&������!�cŁ��&���4_�n@�0�!�ZY�}mfP�?�Yc]z�%����4p���"-<�\��r�]�^A��P):��Z��TO. �h`K��� ��d��B 僿�@+0�{[����U�ʶ4����� fy:���c��rX/g�wW��4-�����ZJ�g��3֩_��F�S�l����!=��;� ^��<��u�ƴ����P���C0�hGrU�3مH��JPсCr�.�g�B5�i��E�Jcy�����c9�N^�&��_�����As�����ߥ9#��S�Iտ�ӎ��U������s�O'-U|jl5�h�3�= H@i��m&:$rLH��*��	��v�Iu|�E(v�����u�u6_F�����>�����OH���{�4�rͪ�GH�~�ix�3��g�V t��$�b�j7ʙ!@�Lˡ/�Q�p��/8�w(%�`d����1z^Oi���C�4o0�Q������҆�I�0��1̇�#��{�(�n�V='�D R�o�t�hN��}Dw�;���o��C���i(��n*Sd�����ǯ�-�0�ѽv�`��_ެ���g�:a�0:N�XJ
���[>g��/UI��\ĩ��x�#)��kSd�U{l��QQ����q����UZKZ�����Pk�G`{�$}OxvD:�����V��"+$3�c�'�6h���QJ��T�g�J��Q'����v���"�?nX,łŚ*--M6��x�:���n[�'YG|�R�Q]X��7���\n���T��j'�������m\�\X�	%J�@eeق�o�oWG.���o��e�o�A:5k�I@��ki���|���`�0F,��f��ueP���IJ��g��H�z�.ȼ�7�"̠s[&�FμpG�V�]Rl���	w��)��V���h�֗���{���cƱd�צCbK�z����%�����%8�h1!)Y��
I�2��I�&����8"������Մ��U�r����M%;N������$K	IJ�9��v��3A�q���v����r�'��ӟ���j��Q��4G9�̞�#��JP�����|�5���
"�
�(gi��a�UQG���mI𢌣ۨ��zcO-n��!�N�:|�@tn�.4+@w��r؎���7�r>!%��đ�M^>���o6�ꖚ5q�K�.���B(�)��@ڽ�;{�b�t�g�xR3�0F��ޔE��"�����m,[�;��d����Z�枰.
3Vs)����驂�kܰ��n�*?�k�(��_�*cD�-��2
\�o�C�Z_V#�#7
�E��j5D}#���0����ݘ�D��z�����=�?Z�?�3��˝�F�I����-#�1ūMS�=�X�������s	U2�;��W(ù��03�� k�K�O&Nj�����G�� V�z���y�@�#�)߆�"ۀ�8��D�T�eE�M�]�}��J�_��r9����i��ØxD����b��-�̮�bӚ����on��]3���� �(��2"Wp�L\�ț�kSq.���U��is�p��k6�̽�3(+�����X���"�B��A��]&o2������r��MV�z}�c��砲�.9]o�k���-o�ۯ���?��Q	A��z��
�>i�0�Dऀd��Ƚ&e	�R��B���:><7Ս�����'�h�N[Zk��Wǒ}���V�l���V˄*�$a7J���o(��?5���8��/���/�J�dd�*{ MM����Q�/�a�A!�֣ �I��^>�F��w��W=g8��,�6�py�oV@O-#�~GE���2{Q8�Y=��;��C�W!�C��gvЎiPa��LSƤ��z�ʯ)���6����qk��Ig���k"�"9��`�q$Qܳ-8vī�^�w*���B���.v_^�j <_F����n�j�2zX0��{������*+�/�h��J�`������1�\K���W:o2$I5�&T*(V��V�7k\4:b��[�(�bg�'�������LX�c���me)"�ş3�����;P�M�oЉb |���	A�/0@�Զ�K�)ۣl��-�S����7��+�Ɲ��&cDi����;/%ƞ@L��N?.�._莘�fo���ݕv 5Y8�ԫ�L���򼷫K1"����M�,H��"��d��Y�S1L$s~Z��$�[w�z����Bn���W):*i9$�>[�6ᙃ��B^wL�Ⲡ��%�;# �~s�����T�ZL���lWL�^�K��kq*Kg��,�{v������VbT�\;�a�Şpu	��鱬��Td���@N*���`�y
D+�H%�$�Q.y��uUwh��O�����x�lZ������9X�ߎ��f#2@V�u�Ѻ�x�0�Zo�o�̓ɛ�5��*S�|��\z��̎W���k�_j�^�H���߽�;R�� RK�y��o�>��[`�	3�C(W�]��,vi���g�#W$����W�E� ��R����ꑨר�)L�l<�1���k��v�| [� �k*Ev���:�ŗ�t�Q�!\�z��� B��e�UT��C�#���afG��.ՍHX���
�g|�^E�n���N��;���ߛK�J��Aw��[QHhؔ�	�U��/�>�R%E;��8��-�jU�����[�ѣ�ӿ�&�W������K�8���XPbS���bZ�T}�a,���ゝ�SC�,i�5���*ƪ���c:����"�&���P9 l���n�!Tɳ`r.M�&�f�׫gӘyi1���lP�����SM�x�H�/0�9�"ݲl]���c셀��N�xM��~�V$ua�_]��e�\p*���%e��Żf\���Zk���� 2>��.j���𕡑/Q��l�0���A9Ɍ�|k�Jw����zv��5��fgP��8�#�B:��!HX��\Ӟ
 �I�a�/�GC�w�������D�G��V��e�Z}���w�c�~�1o�C&n������Ȕ>@^U�8@��92Z�C�D��	�rX�E	4���i�yg��t�=&��%�ܛ�p�]��j$�c>֪��pO�/2GR	���[�_ҋ>���$�̶���2���@;1�(I�?���"�e����T�_��b��W��zB�C�R�I�te3L#��`�$麷~Z�Sv0�3lX�02ܫ,��XJ9�F��V��E)����-F�9�c���=5��,ɬ���Zh�`�X�Sw9��t1|�8'�'YR�o�?�T���Z�U�~+PRښ��B��8"X��s��m�1?v �=��;)��l_Н�!�	��2C�m���z�CFv�I=>� �+8��c�P����������
��?��%���
[��=���5y�����(�f&f�CP���w*�P ��;���H��|��rc���N�������@���xqir"�i�����
�u]&O4��[�>���sܙ�O磧q9����Yc�@�7�tw�l"b
��:$�k�3��}�o�HVL��,E���?�`�G����L�?zh2<�Fؘ�m�����қᦼ�v@,d���RfO�.��/w�K�����^���j1��Fx�{���.���	f��F�%�0N�	���j�ኒ$�  )�b�R�N�oX)�T�2����]XX�Bg��e׸Ǔ�q�v�+UJ�9c����M]��^�dˉ�d�a�~��zƅ��>�[@@S+�Vq�I����㻓��#��e��7�����^T��''L��#�%�ز8���g��bWn $�Z3)�h�v�PV|M���!L��2���VD����Jh����>TGZ�X�xo�C{�X>�R��-���;�������&�Ou�[�'J�Ю���l�(����F�����"PG�7l�^ ɛ�8��\+高� �~$� �����t���� ȃx�q�f1���8�"lm4��P��TϴIѲ�KW�U�z֡�[�!��9��f�8ɒ�TY�gr����4�Uaq��$&o�����Bu��B�xW���K��[��P[�`�
��6[����Y��B��(�������8���2M�5����I��f�&���<�)&Ύxu2P.A�Ugk��[����Q���h������4ԝ�)l��A�8Um"
o�����20�욧�a3 V捣�C�AA1�2��W����b|����uvU�yt-;c�Û���-ڒ-�C�ۣ��Sr�b�#+�e54 	@'9�fX��G�$���7���G.�1�4��~\����l&����lfv]����-�{�=�9��-.|�z�|�;�͓�>�6S��#�����]0%Ȏ�S�K���OG�^��1����ju�����D3J��8v�V��3��۽l��ȍb1������:S�Emy�y�39�U�_ԋ�N����|�j�=����Fp�tي|AE�n�I%��[)��WY�i���u!�,�����`��6��Ii%���Q�v��I�{�+B��: (�l si�I�MT�C����kY/̚��TC��cK�4�:#����_ȩ�'�<�4�t����%���W?��K���+W3��q9}��F���o%U�lē��X��Qi3�} � /
f��-��V�
�v�<� <�Me�!�NJeG���7��/�ת?&��q�ݨ��P��� ������]*���s�9�{�W�$5FK�ow�̌����j��g�9��W�u�2@b�6�Z����ި�cG��^�.���4���M]H-I���^��{�ݦ*K/VP��~u`�=`��=�zDR.�����6�+	�rz�� �o�t� ��;#�#�y�J��k�!�Hl�y%�C��ڑ��ӓ�ޥn�~M{Bf�ώ[FΎ�j�*C�@�G�_�a�J*���E��M|���y50����l%�������͙}�e*C��c�[�W�� ����;0�R�8����%��� NJ�\kS`�C�L:Θl�����A�^iq�mv��k�;��Sܣ�=v񁓆�[���j���,�����긽L3%� ��k�+��[]6��j�b�#ǻ����npNB;ȶ�~��X$W�#�ψٚ������>x
V2��l3��6R_��
��U���b��z���,��s���oH����O��m��
C�����Y*�Ez����|�F�.�M)0�[�+�-�`����䛌
�7��,CSf�DU�5$C�ߖ�;���A�A&�*<��/;9]�ʌ�fld<
`����5yl?��G),�!QZ=�)򑬴Ō����dXt��og�&Ǳ�P.U�%Gk��m;���gA�B$@k9�^��������S�6���Wi�WN��9
���M���h����g�Mt��-�3�Vh:�q��a�v9�H���S�τ�0~\���ןN����[��|��������R�����Ad�,�W:�n��>�TT<Ү�dpC���C1�^{����c�')$���E6�|��s|� ��0��4��c]����Hu��?�u�=��kE��y�d*l�f:�P����b�>�8��;�S�lO�-h].yvC@tx���2�}N��2M�����@eHD�����W�/s���BnIq����?_n%�����r0�����%�z�Y&~��5\�|�����{�@�ٕ�j�����K�iG@�}��.q��Z��VV"�b-Ό+���Jb��P��Rr��ʖ�E^�X�זW�����ݥ
_���o�0�f<�k��*�������0S:PO Kx��WMzNҗX�lR���m���]젓>��,�T�Q+�Ma�%B����N�z�����v#�&,�6����q��(.اm�+�qF��/�fk�;t! ���B �����R	E�>�hk���-�l�������C�����!��L����!ћ0��q/'��(�J�&I^h���V���Pn�">��z�Y>���yɫ�Smт*�+O�B�@���ՠ���{��%u9E�=+�-���R.6>ZU�Y�K+��w�pč��[��N�/#o��h��l��$�;NQ��R���Q��{���;�{�~��͢�@�TQK\�!�fjȣ1�w[�q��ceα���%0/L���{H��� �o���Q�M҉{�ǒc��~���G�z'5tATb
����Fց�?�S�#�j�sn_�{��\��]�Xй��(�(챷��Yo[;� �֟ǂ��й�E���#B�U/�=7����l:�L�[^��\B/:.�&�|m<�8�e 2#�_+C�!^���n���O�hc���>�&0��͕��T��z���5f��-���s�1��yH�B������R�+�^4#cV;��8f�8���k�)��l|����;��۫zf3�2s|wU��/c�����B֧hIx��K'����\�0w08.�f?��lHP��5��1���M(�n(Dr�jO�-1v��1^J��<@X���F3,1R����˩"�Y/�k�2����;�1A}����� �^������IU���L2vȒP�2�C�#j��aA����%/eo79c?��u
�i���ÌDs�5*ƸbR�_۷Gϕ~�F�\��ݶL�e�eD-k>���AoɦT�fX�������q����d�I�l���yIk,X6�^w��۩/�8�s����ٽ��H�~o���1�-J�������1O��D8i ���&/s�F{Q�7#���I�Y�	D�4E9CPj�ֱؠ������/�N�!�}�JH٤rk���������_w�/����Yb���鵡����e,���DO;��n��2詀Ck�Ojx�Qw�6O�5�?6���"�U:}n��Aᚵ�R�gEg-�r�.|���zNq�&���ta���9[D'c���L����ڕN[�����ҺB��Լv`媒�x��O�8��KJW��%]F��bZ�� Ⅱ�����
��v���A�_)W^�����]؎�Y(O��zg3��(��c���/V�tn����{ݱ����J]#�%^�t���u�ULv	�c���i_�I3L��>�E��#*�<mj�P��hY(?��p!��yt�N��w[��疟+%6��ʴ�:���9�
�֠#� (�U���2�ӕ��ܓU�����W�$���[�d��AΌǹ�m�:���0Ld�)qX30揽I�[}�kN��5�v8�S�3�H�Ї_�Q�g���ب2���2�`hspbW'��eF�R��ʲUq��!���/�)��ᠾ����c��͊���[�a%�'�����Pj��C�1 � �a�n	`���҂e����<�FJ����q�Tn��sE��͏,��p9T��,H�坏��/�=f��Hu���Z�����a�~��Dq:�K�d�!h߲F��҆uO�Η�j��B��N3����S�1�^���8�v� P��R�IQAT��I��z�7z���nKۯ��"�("�9�@�iF�<�^�UyΆR/@���T��݁g�?��LGi���!�g�!�K,�usCO�u8;��X؜��.-mI��}���=�	���ZA���q�ÌAN�:9�V���~�E�@.�p�n\C���ۦ'�RR��D|M,�C�1G�0z1� ZF�C�23N?��|��w9�����9
��uY�)&O��!``�s�����}k*	�hc�:d�	�m[�$� )OT��7/+r�iw3�dd��߄���.X
RX؆ڈ�<���K�7�F{�X~;.|��J��5Z��*�?�7	�YX�.�@CS(h��M���-�{��B�h�0h�0���-n��k.&̤��jLf��K��~=;L��Q�ݒ�0���YvB@�L�}�H�1�w��3J���,"dן�:���g���;Y�c̲���ޱ����Aj"�8c��k����">�cj@��9�܎��2Y�,��։�!>Ɵ#b`�\��1ܒL��G����������;�H!��ޑ2]?��b5��}�z_f�Ȉ聈�Rofwt��8��8
¥h����''�r����X23����|����ji�����������.c�W���E7��"WTp�����u]�&"/K[5P�p��"6a}7������dDg���=�j��M2oĿ��r <�d�kR`5VIDu�ӈ��T7�P>���'�~p���i�RPr|��y���"y��:;Ò8LpEL�S�?�37�������\<o�Ct�!{%n?JS�*��P�xp��3 3>2�v�O��
�Zg?r#����T���<&�� �+�&�.{ ��G��/m�Y 3�-$���Eǆ=��g��OaK�E�QdR�Ϋ�q�}�c9<h��Jz_T��]'Ľ!f[IݤH����>��5���2FLO2�mzt@���vF�ԛ����@+�VB��!1��=*�����1�+��t� BWۦ�@���vaϮ�X��"H ?+�>s�J{y���\�p�Ƒ���ƍ�չ�;@Yċ1C�Vq�G�lu&�� �� zT�av����:3�W�:���c)c97����x ôz�{��B��g�r#zm���{�q��e|]���8��v|t-�E¤�Y�/�0- d�6`93r`Gi�\:��>�0��3�\W�4�S�3*l%,&����ıU���WS� �mP��ŇZ���o�@���"�V�ŖTI�ݫ1���#�hu��(ԧ��g*�,�<��l�m�bF��n
�`��\(k�1�^?��+qzYs� ��7_�a��"�T9��D$�A	I�&_�w�|M��p;Z�M����Y�Ff��{J���_t�GѢ|��(��NA&� 6}�7v��lD;�ό��ׇ���20R3�h��dmP�jMvH��I��20������i��h~HB������Z��CC;��'���]����+gGV��ږ:E�L�B-� t�`H:�u�%��ta)�N�H�Sb�Ӱ�%y��2N�F�O)M��\�mfb�</�K5]��E��άW����/q-������?ķN�;0bsQ���瞰<�}��;�"mT� �8��./�2�ʲ��v��o��߆Љu�HVA.���Rv�'Qf6��ݾ��u�^e�o
��'e������>��̮�+�p��Bd�c��\fZ�qI.�a��|�o�<�@ܫ���Gߩ�!��B�IE<�s����'���9o�DTBun�1����&�GЀ}4*D��h�ȇ��e��jr�f���.��J>z��M]�	��Y�!���ڷ(�A��5�۴P?C�W�����?b����0(��`V#������q��Lr
dX��H�O�d������M'�B�A��`�������D�Ð�9��ׁ���PF�]`�V�?���K�l�޷>���N���m��I��t�aY�g����R�@c��b�{��[�1m(�0�-b\i�s�� ��T��o�ɦ��[86P4(��e��`���DV�n�!w\yR�nv��p/�~� ��Wuz��/-_��\=qm��U�bK���fV��7�ra��+vR/@1_aS���ㄮSgw�B��hxV°.�W�^�0k��J���3|Du��H�n���N�a�<h-�ө��ŦM]�W�ܴ������g���aj� V;�ܮ�Tl�8� K�v���oD���J'�@�2�h#k�D^�@���{�^����)�ux����כ�SRY�O�;�2j$�.��[h'�ԝ=��/�����B6O���v=x}�]����IИ��n����m���u��וT�zu�m��(�@e0�����9�P۴��UZIWѮ�#=0[��h�o�K��NF�.[%�K�5�D�U)�A'�G�zO �9G�f��n��A�p�7�,=&���%��>��L�n��8�v0�`PG��/�P�����\WX�0T �m��T(�'G�%D�cr���?hx�j� �:���z�b��Wȗ��jaR�^�9��=��|S�ײܙ 9���*�j�a�?���`g4���1�	����U�#�� ����5��y/6������p���i��>{˭�}VL���z�Ł*@�}@3;�7���kˤ4���fx%�;0HAw�J+Dh�V��ڕ8��7��# 3LM\��c�%�{�����D�5/�zz3�D���t�?,�I���=xE!����v�:[�9F$��,Ԋ��>�ߣ�y5z�=�̖�˱#8�'B�s^�"��{:s	�r�a8�vŀ����������
V�;�S�V���L`��N�)�D�c����c}Ó���/����������1c�DCli���Ty��}}~�U'႕y���� ��TP���^sJ��x��K���Pp��n�~��+n��(��gL�k�c�4���ܯ�� 	�B���d�,Y��]f�K鳄k��q��{{�e�v�>��G��A�=	w��="�D�7���%��?�E_�=c�GHţӓꉮ�\!��7�����S�l{����V�lI��B!�}?<q"'?h�����i+@>�5�J
g5�3TV���?aBNɰ��V�3v�Ϧ�ίy�G�;�l�x�e���Ł9#�a� ]8$��}�2l4R�S��n��ّ��p=L�%�b&���g7p�I(���\�o������.�~� x͐?�S�ò�T��Ъ��I�K�O3�?��*��h����F�@dH_��W}c�6�)� �x��M�+�/Ӗ^S�XF�Z6�-�-�
+��5
�	���;����X����lf������.�d���<4h8yZ`��ފZǪ�]�M�ϹO3�y���t��M�.��G͊�,}9��yo[�^���(`7�*"3���MZ�s���>�4�8��\���)��qڨQL�bJ�h����ϵ�9=�3 ���B��]����D���*�Ɛ0�Ȫ��b�Oʿ�T�� +�F�U�)��2�l�?�z0�?
�z	D�[�>�"��xx�����*�ܕ�
�e���Q��h���+e�*�2}�9�竏Fqw|�@�Q�a*S�w ��E����k�Qe	�`p�ؾ:!�{�l��^N��W�^�~��S*��{�h�?h�Հ��/�f�gAX)$#����C��z���[mW$��D��	���L\�b��,[���y�ye�Ĩ��7�֡ASN��4������U�v��P���t�s:�l����62g�h?�!�� iNɡQE�$q�[��܁�}�:���\kǳRbM��H,+�,T��	�������k�(��a$��5�����Ʒ����%}ѥsH��m���/u`�xQ[�_��?�]/_6�#pz����5��*WXv6D,��ai���2�3խU��g	Y�E�夐U���br�
�n}jѧ���z6�kǴ���q�����Pu��)d�&�T�Mɖ ����\�g��G����&Ѐ�+�m�����������HG}D&�U�E0 4$j������q�ڥ���,��R��8��#`C2�����	Fg�I���/��� ����5�`�e���E��E����2+l��ًS����;�`
��ԑm9�cP?������٬8��ϳK�44l�����3�e�zYK�Ќ�f�����yY4�@Y�	�+P�;����޸�=��g�(��m����������/�L�L��_��>N����AJ!ܪ��ܑ{ɥ2hFn|�&'36�_ �������W%���0�a��|�*�v�3�$��)<�-�S�.C�X7�A?�B�^�8��}]7�!�f�n|��Qb�[9烝�����?M��{�ݝ�c�E�_������L��b(x�ΩQ�im4GV�I����9J�ꇉ�'�q��1�JT�VQJ�s�c�X}�TK/�H�-��2�'�g�g���N9��t�;Sf�A��v���N]3s�6F@�B���r�ߦ>ηݲ8��a��`����"8�ܨwC���2�Ay:X�rw!�����I�d`��`J.���$�~��!�2�f��?oڃ��PϹ��x��,����Ӈ�����7�J�U�>���X�)ä]��%p��=}�7~��.b��@?oٝ+���,���K���]��u�������¢Lp�ǃ-�X�`"�
�rې�_7�/����[��uz�3Kt+?^Mw�š�?������j$@�����ZFsA��Jv�	mf>�B5�y��-� s�}�3I|?V|�R�_=v^�U�HI�}��d�uc-C�!�����z�F���X�dh��c�ay�!$�bk��pKyf4�H��S,�I�iռ_i�����Uk���A�lp�'�fKy���
�	�y$�3�4ɬs���w͍RX��I�K"�Qs�{�zao��fUr�2�ű �KyR�V����R�CT�2Ci��sf�&Bj�H����X�_��b礼��h��48�&+`����w���g1|��*E�7�<kZ=�V��I,�ؖw!f���2OC��i������°��&���a�(K�/ Aո1*Xɧ~����T������l�c�h4�#�'�e���IS�0FH��I2�u�$B�/CXf�X�Ҥ<��5�Z*\��_q��my�Mv2e��;N�j�W;�� cl�k�9��'�����2_�U�'q���4V���{)䂴������Ɠ���_�I7�
�M�x����ZD;��bPq6_�?�.1�Ic���X����Vb���Jr��(��;&�Sb��h�V�CD��]96(���'���^�w��:�)�l�*�c+��w��4r��sK��+g�,�
;?��]`Y�Z��NV�7y�A�L�*D��@`��Q�򋳈��ؽ��_�?h�c�9�:)��w�1sg�����4��F2f!��f2j��PS��w| Q
�3���=	�A^�6 ���0|�&��&Z��ΠPM#�L�&ۥK�T�X��vބ�1KMD����3o��@�6�)L�k���%��ʼ�=���L�,3�����4m�W�C�Ë�����jJ��֪�P��π�nfi������K��:��,a��-|��|�*�3(3����v�E�2�0�1$׆�A��J�4*-᧕�0Y�pЦFI���~��CS�4+��	 �A�y�*�� nⱓ��-oy⮬]�a�!�;�7�X�I��9�:�R��݋���Q���2�W0������;.��a��'86a�o�]L����,�p��1L/O��H�bvt٫���l+�%���(��@2�z��rdλ��!����h�%�7VKT�⦧�D{��}q�G3�} �����aŖ�I�_T��)���@7'�?sp����}f��c��PvN$�LE,�������s�uRvD�`^n�}����s*G��72�f����.�0���ˆ���:�0��Ŏ֗n+��{D�z6�\ϺէcS2�S�b���C,U���dQk�`R�*�AX���h���_��C7����M����#�5��hf �IB�G��Lj+8�N&��ͼ�)P���2Β��J�cJ��Ie�o��5�i�w&3��q�&君�?��VU	Q�DZ#�g��v<����4�Ͼ�lF�����y�\}C�2}��C��\7�JU���E���j>�U��Y��(����zྎ�R�c(�3ol�p����!�xĄ��N���Ya5�u��dx��	���r���;Pz�D��в�+��E���$�I�[��W���`�H0����2X+l�$�����SQ�d6�9@����͂>�w�z����N'z�4����de�w���ϼt($KW�x*���l"?n�3�����!o��(�[Ἅ!F��B�}�h-C�Z͑�����( �ٽޘ2�s���%�b#���%b��f
�A��IG�dMZG@n1{ -���6y��%�'��X9"3Q�q�8�_�cK4>�K(��O����;������J��x&������bQ��>��?����S�$J��O����H鴜�z�P���SB��x��U�b#�f)� X�,�bYe6ݳ��	��ud���N=5A�0��l���6�Ѝ,�+����.G�&:Җ���\�W�5k�3�v����$_�S��^���\i�>i���jH� �l+O|]�hɆ�S��b0@�Tu���GR�5���ӧ�0�i��bS�^�u����-L�Z�ÐH.5�}��I3�T�"��Hh��gG��DwB�xS,S������~۬LP�oh�,凌__�FL�r�4����Ϻ�f��=^�eUB~�Avz��c5��p���/��fN������Ȅy�=�L�ʬp��Q6��o�g��X����Z��%(~$/'�(�D��S�1N�X�wb�$���hz��)�iq#X��c�[��	��5YU�*�@B�C���e0��E�#�-!���`,�d�����r������F�}�ɝQU�y
'�	?��|���'�ﺚ�u03�#9q��#j7[�۳ƣR�X�.vU����j3��r�c'���%�{��k﹞[}��!D�S�[1j%���E'�K<~B�m�yV#�P��?�Ni����[� �kE�
	�!խv�冓�?���SА��%�½��;$L�d�+�P�!^*C��⭸��-3�$�z$}Zͫ�<����ѱ?��Y�ׁc.���a�)�4�����v�C�ÂS[$�rRێ��S�!,1fn�CC�c��7]O���]-s�-H���(5mz��2�ev��3#j'�C�T����o��^�Pz@�gF?!�v��E�� �&ڼ��.�\��@�t�`���{�i�;�M���B(�6��to������\��g�
�SU����(=�`�E��l@C�z_��S.3�㕻�ڪ�@���ڪ�y��!�H��-�u���M�e�G6��i�⋪��d�!<��}dg���va�սY�i�V<m��,9j�W���3���/�w�D�*�ȈW����*b���p�GU)	/J=�`�yD�끾d�R�r{Q��ޥ����T�W�0H��w*����=*�Xj�P:A8���U�?_���;��s�:�4KR�JV6�����$J�w����5�G<�h���Z��W]
��]>th.Ϩ?[��[8��g.�UDj	_�*��7�����S�vhȺ���V�mI�O}9H`xP�x +�-��������09e��ϲ�	�����8ŋ.e��r�HT$
�Q�*طW ���{�&�^� r�gV����7�2�8E�:�1l�%_SU�#��]V�>��¼G��96'��"����chw3.:T��!@���zX��b��[���`���U)�b���;��3I	�[܃��lH��D�Bw�"��@v����f����b���"�-�bw�xy���{#69���f�/)0m�f˞Dk}��=͝�/�ZKB���H(5)v*��<���_���(F�3�����〞�1\\	qH����|�,�^4�1��G�	��|�j	n���1�<��H8>83��ϫ/a�z_�v�;�+���d�{�as�j������	��L-��1X�w~JϨ:YӚZ���WYXt�<D.t[�h�� :����DZF>q͇�����n�D�43���j���7�g�I
TB��-�_�L�- U v��g�Mv�
(e	��;bPI9�����<
�J_��ٟ�*��-�qӍ��=�ڠ3_Cd6��e��i���\��a�A7����q������yۢ�;�i�Nc�^����>�9B�0y�RQ"?��=�@K%܋b�R����n#~�@kӂ��v���l��\��kīCF�o��L�^��9)���c=�#�&� �fu��p�+�>H����6F�EÚ�\v;�W�5�㲏��D0����kb=�d��&1R�֎���X�\-��"�G�}�2wv�Q9U]X��/*�D��[�J��e�ް&�����':�_�_D�oHD���
�(Xǲ]�u��0\�J�s��2*�4I��r���"V�BX�7;�a9gLQ����A�z�+�Y bn�{=;����$�S ������B�'vQ2��ؙܽ!=V�Jl#�s���b�.N��ʝR�K��`9K&��7�l��xs�[p�h�fVwN���	�^�)�j��]��P{�$��گ5�i��&'�*��58Lv��
�w��bQ����nʲb/;ۆ��e�t����T���2��*Z@�oM7u����=@�&����X�ꙋ1�:��V�<60��>��yWUx5��� K�qϱ��u$z�\b9V�7����,�6�#FQ�;��^��d�M`��/a�UO��������RA�� ����Igh��G��Gg�F�G)���<�	)�3��������Y`<#	�� &>:@��U���ođ�O�{ɦ,��3 �ъ-���83>���q�+ �ބR��[e�x4��i�͢�p#��V-AzK�!����c�c��T�;��lk�D���>�9b�=$�|���X�2�S�TC�h�lsʟf�x��p������7ol]�PԾ7f�"�ע��F���X�w;��ʹ�bB-�Hg�-����+|�&!�9�# ����p���<l�&���Q�H(�H��qՙ0s�o	�"%���p���P�<� P�-�'߹��d�@{���rB���|mFp�����4d��K�����u>�I��;Z�$��$W�����é-c��)���YRC.�;}L�;��S����>:v��Q�3{':9p��k�.��Ҧ��c�q����6j]����}SC>o:���[�j�aj�Y�8��mtٱ<9u��ϏY���n����� �~������J��6v6ԁ��Vb�<�M�$��E�^�يj<:Ð��6 ��&ZO��2;��R�yb�/喐[2�Q ޯ�{���c�ozD��ǥ��չ{r4VO���ħ���y���$���Jk���.n�&OG�A�4����4�2�sP܈ٮ���tB�F�jƴ�?-O�
 �{Ws��P�P���-�
H��о�
�v�[gY��[�R�%2�q���k��I#
�,�5!�!d݆,�7�U�kDB����L���5\(�Z	~zM�`3Far�C�4c^!8��܉�5����[�/%*�v���6�y-t�YӶD����a�R�BG<|	ϩ�W?�a�{���g�����Kr%�Mu0C�*�ytP9����9좔�K��Ddc�7c@6�rɖ��#�K���m����/b�Fb���wuZ&i+��oob��C��s�_�i�2�cȯ�i����0�E�`:u��ȿP�%Q0E�І"y+1Wr/�*)B�8��n�9�h����$���,�d�O5�4�
��y��#O�3��Xs٧P�"�� �x�d��n�}�9�0�eK����K����BB�B�����ב4�S?��	��!"�dn��3cc�(J
3�Q8h�pjL��ڸ �D5�1��#�,���-��&���:O��R����R@���D�������8�q�	}Ӱ�	�C��	>#a �]J|a_���@\��G����V�1����Viޑ�Su��z�a�"��� �,�r6#���(m��^.�!�*�)���s�FU�� Yz��ԉ�Y1o՚xb���E^2�U E��Љ&�R~���欤�rV��O������l�Z��̺�ǼL��NG��Iϛ4g^��cYe'�ǰ��7XcL0:��6��}�j��pxm��h�5-���^!c�i���f�LZ�P+Fe�+!n�@�Q�b�xV!��4)�$4/z�mܑ�{��񜅾��<M�?.�/�Wupv��G��ц���f���O�v^ �J;�ِ�EY�
,��	�2{-~�9��=�2��	�x?��>���s+i�Y���21�io�#�AWC�:��+k��i�i��Ԯ�9��f��^^���6��5.d�������N&��C�,���g�iMva�2ؙ|�,u�R�6{��ӑ<AC�n�=aL�eD�eUP�����()N��kR��P]U���x1�=��^璤�3̇R���R�.�<8%g���o�5X(+��({��N���QC�P��\' �d~�s�����x��h���@wlKG�TK��U��D����db��j�L`����b�u�a�V�.�D�65�=x�VeBWЋ;n����vuU^6z׺m�C��	$N����+C�A��ҫ��\6*�OR�4��Q��.�����"�ߪYx]�!ٱ��%����c̀2\�l�^eO`���1"pM�������?��oډ����)ۜVZ`� y�L`B��_7n����N�ӿS��iT������s5��˲$���P*l)uy4� ��d8���D���ĥ����&�<�R���{�ٰ�gPt���{�DY�߹�: ��~��y�����攋���O,&��jYI(�t�������Â�����VYz����-L��.��#<��N㔻"^�����ݍ�{6!���aI�^���m��f�*O#�i��׸W�9�<N�ө>8r5Gڇ�hҐ�5��?��,�ylτ%NSL�4�U�g��"���nl��
 ��JS�%	�k����n�;��5��e�λ#�w`���~������#�J���}J�<�v����o06��[�����1Y�ʹ�S7;��O���2ۀ�!���r�a�h���i��C���sW<��+��5��n�;-j��
�4]A���;n�0N )����5W�-M�aS��I�����!��%m�[�I*�6}b2�V'��I�}��ԑ�_�x;N�D&M��`�zhu6҆�M�٨d��	�<S�ڎKi>"�e[ֽ/�����ߪ@;��F�6b9Z�S�ǡ����cA�����5J6�f����L�W1 &C!��[�7�Wi1%�k�҆�F a�Ik��f�n�U9d���No.��lE���43���ż��,�$�
1T�.Y�-O��>�ZR�@ *��`3;���A"Ԝ�΄AL���i55�e/9A'y2!EsbN-^���!�_ƨ����+�"��=�9����!�c�͕��Q���(n~�����W$w�C�.6o�������C�;ǔ��Q���T{�����wg��u8ɎAw��F}8.	7��0���V�UM���3�?B$fL^>�{a�� ��� [vFˡ�D�l|#3R?�V`9���!,i������gκ�~V�y�����fYy����Ș�`��]��PL#m�}a�d�Zl���K�a"6z�6�_jrd!��T%ZFm|n/��M�D�!Cl*8�
|-�E�!�wvaE�9�.:�Ɲ.w�n��9���Z�ص�9���B����Y�SQ֬V��m�<D���%/������VW��{Oo>R0Е�|%99��ҝ$���$�$x�r��t�b��w���x�Qݿfj{�~�� |�Y��.��A�o"PeQ�����������	�"�s+��m�َ�򩩆dOFo&#mP^�[ي̺�!������*B��7W�`i#\
8�+����hd���/�n�m��!��S ��zo�'/I��5x���ˏ�#�K��'$�+�w=GgN�,n����o��m�+������i�L	���P@4��F��9�\�gj�qT�C=�&����_d`B�� >Ǎ�㋱&�u�HŮDs2��8��(Σ�KS��<}n�SU���9Ƃ!S%��f� F_��OY!����t�E��G���ۍ��~sy��)/�{������*r��&��'�� �a��܆d�򜼳m^��W(��=��Q���i}� e��Vz�3�DJ���Fj��z$q�b`���fL��u�Cx�Ƈ���E����(-�BE�*
:e�����?M��,�J�AM_�F�%(�gf~ˌX@k��&����즀���t�ZB�ɀ8u�H���r���9n�3?6r6XTQa�h��de�[h/oڨC���w@���ɯ�!|�ȸ��ݚBLM�A�����}@��ՒAM�4���*_�WS����}o@ڥcv�H:t'�n1&EE�z����о�ǳ�SB�G���uggp2W`-��j��L�wЗx7�����)�%��d��HSZ�3鼤���S���&~�Y���PS4Ji�"bk���hԦ���O@����\:��A�v�-��HM�a�ʔXi����χH�%=�T��S���#�Tݔp��0RD�`��3�5[#w�C��jI]o�2K��'���G ���CMī��)��SBnǈ��)`�wl��S ;��h�Cș1�,��
Y�v,��0*Ҳ/��;	��T`�!�����^���A<�&���-�`�1�>��9�h���+P�Tb��i����������$��{��`2�l�Î(�.���/���(�k��I��J���-��� D��YHfV����Z�aW���B��J�ע1��K~|�Q�3'�����3�Z����u�4g	�'���a3XhH��ev�Iu�4jIAᦤ|"f�G�M��
��I���T>��e5j6�0�\T��Z9�� së)��8���T�Z�� �趚�_<�c�q�-���"�ЙY�����r-m	pÐ�nQ�1��s��/�O�,}U ��rb��.#�jd�dRA�}N�#�aE�^��/���� �+����)Ӏ
w}��{�\���n��߃�{%qė�\q��q0t@5ͣ���UI��9�3Y vn4�w���ޘ9t_l�2D����Ye~�R�ue��T��f�gtz�����v2��d�5��F;��T:\-PXP��9K�MB��}BQM��<;��a����~���zȔ��Th��B�Fzx.��~~v�>p��Xq̉�^I�v�t+@ ��Q���R�OY�k�u�2y�_�q��v�2������:�x%]�$��U��m"H2�l����6����Wh|M�*pRx�2�F�V�v�ɻAns��0ty��4_�V�J����s�����%���N���덐K����Dbä�GZ��U�4N$���,�^��J��.�����_��v��RW5��|4]Yt�f�6ܚ���ɐ��/��o Q[�����������i�A0]��Gr#.���
�㢘�)��e��fk��~���J����|��e��S!9�?�#�\�y�AO4�n��<���<۠�0���p[9w���x_�]T�r�V���&�c��`6��Z%���K�yѕ�����D�m}J�U��(5 �|���[��g��^#���%��r_�|_Y(!���9{����U�H��a�zN &���D�h*���m������'C�FӘ�����#0����~��Be��E]��y�v��7~��T��	�0M��0��퉱+eT7�uq�x�NJ�9�0d��I&�%{?2�<�t|�4��@<C�.D�� �v���*Z�����ͳE���<,	�P�gֻ�^=���Q[0�*PA1ct7m-�Y� �(,�t>]�D�	;|2�����@��(����a�}���.E�)�/9�����x5zӬ��<u4�˧]KsF1c��"�;��E��쪇D[�y�r�O�|���8J/��\*>���%v�E�;$?A@D:}�j�������a�}:�a�GMNIVT�4r�	����3�}�U,���Ћ��7����%��s�9H�� �sj�\B��v�K�,K$	����FЭ�7p���mB�}�iC�4L��p��:vL�ڻ�q����rS1竈�M�*�0�IVq����q�7�Cu)c����v��o��S�H��E'X&��yO������k*�yM������QG��_��R�kE����rM�g����(�l�q��]p�'IPO��������Q&���dW��B<0�x��'$Ш�?b�)�0��OV!hxdoO����x�HI{"
�h�UR��$>��A��>ϙ�Aq��=�_�9cL��g�u���{��kA��|�|��
�-�h1{���.c�1�G�.L���AnB�XR97o,ƇA��W2��ߵ�cA���[Jw3�W��b�F���9O���l�؊�O�J��=�>u�������:6�HR[l�/H� %�X�X��X6�Ž.�1�&�2��9�BH@���h����,�<�)���|�(�q�m#aW�L���Y�WȋƉ�b9�hNU|��_�4�c=��p��oy������	g��ˆ[Q�tW��j�NY���k����?�q��[|E� ܼ3"X��	�|3=�ܱ$IV��3�B�b��{nr�	D��;������ �W [K:�&;�dR���qB �hz����z*�+�C-����b���=	���v�n�P��z�w=�u%��8�PDSd�^�0<������VRHZ8\C1�M����4�E�(d͞Z�^�*Wb���|�#��=b4]��3j���i�o�'��CM�]:�%�Rp��۳#�ݦgZ�`�a�X��ܜ\t��:k~�5��sr��\�f��ށ�W t��Y�^����5"���7�Q�F�tDB�Sq��'�<j=�:�����1�ϼ�]��z!�0ri�D����uL2s@� vbG�RqY����Mbѧ`���L���|�����A*���:��	�?s�-~�"m�M���ɜ%�/�����HZ�#U�β����与A_r)}/`�������R�Q�h���m�`�1�ڻ�2�9K��j�/�����1�w	BX�|W2��P�������+��к�N��xq����$��P�_Ň4�R�)���v��~Q���WdɃP��߁F��5NVZ�#��1�d2X��#c�c��=������o�9+����pA�t��kD�:�-�7����v��Z���8]0���=��BYڢ(y���`���I:��&�t�`T���\.�����X}�8
n����\��ֺb��p>��h��*�q�4��1���2:�C���Z�>��`4ܩ��닟t�ғ1xg\���"�v�5�!OC�a��Ec��sQ��������^�����.OŐ_s�U�(-���L&94ƈ�W}��oUj��Ge������w�5��l�e�w�GgE��3d������d�U��Z����Ƅk�O�g7�B���.���M����bݡ�_�!����9�����D̰k���fDˈok�/���v�dp- 䍷3������zZO\;L�ω� K�ڦ@{��]#C����n�\���	����
9���}�Ѧ����@�ͼ���r�=����Ymn�So��)e��,��8�3d��|����a⎃��@��0���{gP��C,�1	}�U�
�L��V�� ���ψ3�,���0�/L�Yf�)n�� �\Zf?ƨm��W�Qw�r��<��/A�MN�R&`Ԋ���%>��cU�/y��.��FI�i��	-d'�&�tf���k�z^�B ��KC��Y��{-�ظ�s��?�T	���N���n�E�ךX���^ɉ'�i���L����֡U��2ܲ��:}<��ف���{�P��]�I�sk�B�n[�D�
�ʂ��Υ���>�1H���3�,e��Y\��K
>B��cUA��Bj�x����;Q-���M،N؇�����c�ߝV�6[\���-�v�C���>����d�5�����R���*D�ߍ��k�� �= S�o�X��k'�|drnnB��@�����]���j_&x���C�d]��\��BAӗ� &Y�N-���0b���&����5s��g7�uhh���S!��$��A_��*�?�����s�t���a"{�Y�=�5�Y1(����j���!��un'�Z
-�^��ݷ�;�;��]��^8�b��#8yK��V��g�TҼ���G���W;����N�F�E�$2��`K{e�,#���H>+�r�����`��ƫ!\����5���������/nIOe�=B�Z28<��i������Z�c�,���7?�Q~{OJ��c��o:��% H�[�#2�ӿ�۳��3*����Љ�D��~'��6�DE�\P?uu�#ORE�O�n�A&���m�,S��%����p��`#6�h���vxęT�Gq}PmL+�@m���O@��#8��x_E�����0"���0���	:�UÕ��S���Q
f���י|���n�G�Gr�B�%�T�16�@q����wZd�k��l"r4�|-=�th&bl�n����������̼��c��"�5�������C�ɦ��$c���H���bl�G��ϳo%1�)%�.�ûd7����wn'��'�z6���_��%�k��WSdݴ���8|���������=��,���S�ӕ#��a�_(M�/�k�$H�Kb&��UI�\ԁ�� %�e�h��6&ٲ�]yF�W��3#����ku�
��\ٙ�"�ͭE�#��\ݜ�cϨH7$3�k	��j�;�U&�
� L�+���3h���}�%���s
qXhoW���}��G+;{e��j8����� J/YF�V��/4��F�<��X"n,ä�R4�?Y�j���	��i^c��-�0X�'�R���'�%�1����y9��^��|�� ���T���۾������Ǳ��݅�k���	����k$���$��4	ޔ�k5y�;?F�{�**B��\�0>)�d��g����\�� =`��/%���b]�9<%@H�mf�\�G:��5��Ǖ���|Nӣ��"!��I��v�w�a�.!�΂�B���D�Mj��<�8�.ue1�G��IY�y��p�(%��h�k��� S�!��v����g�E��K�H�j�u�b��8���t�Ņ[����|g� ��s����a��&T�a�����,a��NY�y>���~:��N���C����[��^K�]x,�M]	�l[����Ƃ���O� �*�f)^o��}R�{4�$����\Q�w��إc�!�6b�E�W�d�-H���}e�����<�e+� ��Sw�{i��<��]IJO��\ ���A��m4밊�n#��֕l�z��{��z���z� �����/��"FD_�Ǣ5Ŝ���J�K�ENA�?Yt�;\�o6(�'F�,��o�bm�"��I���9,z-���+����u�����]jn�u�4г�:L�0O����|�����荷�fn�c8A|���J�@v&�}��s8�/;���P%B��m�MD2�4�F]�/=!�����ëq�e���Ek�K$�9�' q��}N��(!�$�������)��s��t���ON�{D��5,�\ZRpU���T��UlSy�qu�E�'.�	� ��y�H�#8('5��ɁĠ�\s��-�Z����ޘ{�YPyu�>�	���{:�Y[�^�]�|��<֭� ������J�b3W���X�q���'���f_U�a�1�#᝴�	�����,�Bv�z��ZԲ6�9P��l�.�2U�H�l�R�٥���˯��ޤ��!���/ZJ���ϺX�c���Yz�~��+e}���p)FԄ/�jf(�^�c֜��.YoK�� �@��?�����7��J���"Ĳ������(�_���U��*�;�Ie�ծ�����T�c��=?r4�����_y��*<�����kA64�=I�ƵJ�+�&D�H����K�lWRj�z��x��5Mߔ6�щ���Iui�p�ou@ϝ�ls���3#t����o��\�*iQ�_F'%�	+.[E����B�"�	�!>���	�K}H�֦�rV[�Z�8}y��??c3��|�q��S�`S�E�{&�?���AI����Ƽ=S�
NG!Fs�<��(�y��t;2̔�ۖ��x��!X��V2%�]i��)�ÃT�����l�j����\'}��tW�#F�p*��-y���6IxwbR��lq?�$�BD��0X�o7�YW��r�GWX�5����s`��K�`͏��bsr��S<(7�7F��=�-��5h .�8��[�.>$}?��c�U���ѓ�p`L��9ƪ�ǃ��iup���m�i�
'M�L*u�o!mC��I!U�Z
��Z������V���ؑ��[��q[2�]�y�m���ӂ`E������e�1��	�~X]�,�uO��b�6-n�T�(���RN�+�[�C��Tg��@@��GI(��)��-<ge�Y����=ϝe��@�<O��V�	G�O�<A�\hB1��_�	9�HG����&����	�H?�+�	ƺ-�'�[?�6[ʸ��kQ��:�H���d�@V��B�@sH����fY��E�F�%����� k��A��)_RG^"�'R��mP�T�܅�����ꄢ��u�L�F�g�,�L6���^8p+O�(@m��/����a��&D����"��\鉀|��0��毝V'�J�*"G�2�p�zb��C��}���fC�LeCDg)�K<��Y���2iJ������]��*J�C,5/�8���B�|����k�2�R��;�X���ُd�m�õ�l7��d�O���B!�6�&�n���E!>o`T�IL\�l#g��5����&��Y��=\pE�����lF�ǥ��7��!>пZ$k=	T�k�F�,0��}TX:"��b��q̎�EM�0�V��%��S�gUΐ�_l� �d��Z H+j���=�M���G��B�&���)ys�T�g&�%�J�E��<-:E�Z�1, �ҧ�� 	1@7��L�f+`
��ks�������%,^�_	�Z����������\t^�~�R=�H.��Ⱥ��P�[�"#����f��$Wl
�y������ ؍�0���}�^ʏС/���?�괾-��h��6{'�޼a�U�]����3�5���$_U�����E3*I�:�k3�un;Ŗd��U%�����{o��A��ϵ�}LƊNţW��^���������uY��#|̼>A�(Pp���T�V�{�_oq�G������S�S��Y���`�a|iu�?K:s%С 1�rB�-�Հ��<P��*��@	��Kc�"��B�ZB�nh*��Q`�|RސZ#>�!�Ef�j�l����������͘#ʮ�z�'��j��]~��ϓ����"�R=��`�V��̠|Y�oyZk�^�$-�q�X�.~�/Ư҃u�,<D�JO�W-���J�Xi+ <t���\^"��~}3]��)��r�xs{tZ�P}��Ѣ���������hs;G:1�g�;�n�.>2�9Pĉ�fԗp�'-�C�M"��뚌��*@&|c�#�>fFt-��{Kyj}t[I�����N�u��>:%+�����z��ժ���Uǁj.���.$��D
�P��j������K�x��8f��&W����E�,cm6�Q`��]����1x�$��؁M��SG&�?�c��'�}� L�O]p����,�/E[���p�M΄&[Q3/��uӊl��
Zz^%��4����O.���*�8��nm9;��8ַ{S���6;�c�c��R��V�S��K�	��*��Zksɨ>@�����]��S��"<UVv S�����%��`X�t�-�\R��j���`��72����������UQ?ED$�`[k�W�nk�y�H�3d
X��u(xY�N:�X��7-��x���#�TJ�I�6�zE�E�3O�?�c/�Ua��k�������\�C�h���¬V�?�0X����cc6���0��ݕ���\CKwT�q]@�/ń���~�=�/ �
�	H�Ǵwu(.d��N�ۗ��:����d&��),�!|�FE6�[NRR��I�h4�M�F���Fk�� xE�Rh�B��࿒]!�
s�.��x�Q�����J<�s�2J#BA������v�f���V�er`��=p2���	��|�Y(N��8ʑjN��1qu�X�a��v��V�BF+wC�4��0��&��Ak�^���8��_��9�p\��� f����^�����8)ۅ�c���ܬ����U������yۣ���~����o��"�OG����x3A�����V~-m%x6�G���-�}*�M�#�M�$ɰ�A�V��m��T��9<B���@�ݮ��ǐ�,�Qsr;A�ڱ��SQ�_K~�K�*7����������X������)Yh�@A!w�H r�@e�������B'�}�L�:�Y��t���M��J޵i\;5t�4�$
���s�>d�� �M�JĭF�
m��櫳Y�		��F���m�J
Jm����E^�_z�ą���5/�U7�ޚ҆�k�d��Sj+>����8(qt��ݚ��k;n�F�|�6�4�rn |����G�1����#��Q�z��FԾ�t<aC샾�֫���R\��2߀!�`_�W��G�>��^�zp��c��d�Ū��gN�~��v��8�F����f���W"�U��k-ߙ2���iJH�0Լ��J{��?L�vM�����ϳ��/�s͹��A����c'�)��	Q�%��$��*\��A�EئA��(�%���s�o[��;�\�Y�rɑW�i�?�)��yE�D��wkF]��5�3�	���	�l��$}^t�C��*��wM���j�����w�z��F��}�S��]�CS�k�}<Ƭ=�<)��~�ΰ��U�j�]�*���g�k�L��el��<9f)����%qȖ���Tq�Cq��vXaH����C�a2��"��r�p�#Ӄ�Զ�&S�h�z���-�d+Į,
��w�{�\�QH��Kj�ҘƥY)��S�;��U<�[u��E��я
 #F��x��[���ZmZ��r��&_�G�����U�S� �ٍ���@D�J(ɢh3��ְ��uO�m�.Я�z� �:u�6�hXu�{Rx"��e�)�3Ζ�7��صA���2�5�A��6�NP��jvb\e�y*#B��W9��@8�`��,�>�m�𥂺[��=�vjY~_
�{�P��}�Q�$ ަ��&�ޔєM���O�쯝�v(#�����*V)�F�
>��F;S�I䙌��:�#��]������d'8���A?�)����E��c˝ܠ�~2iцֶ�BP��E1�<�ƚ��w��U{j d�|w���������?N_b�N��+���k��ػw���U_&���[7M��O����}� <V��^̎���c*�(�V[T�=�����g�4"� +����P|��JͳZa�4���t�Sp���ċhw��I�m
 ����-��YZ��գ��7�}��Sx���|_���([�XsDj��ޝv��t��`�<x�1�#�ӹAG.f� c�|^�!��T���2V:)S|';rۢ��5η��2<[I<2�3����-&:�q,�z�� H�A���._����=�������J����b!���~�ؾx�hZb���AV�	M�]eɲx�(���ڱ�c�f�������Yw���:���|��c��"��Se�H�9�Oξ�pgu�t���z�D:�86���L�>
�0:<3�"ɞ����qO�B��A�0<��gP�Pv����n[�%'��������7*��R�%���1�ax���e�ľ8<e��n�5�t�Z����^N`�5[o��E$O�Gv��.ڀ~�Ŝev����jE�=`w:�Т|c�o�'jֻ󽋳u�?D��`�m�� X�ț%툣��)�i��� ���嫩,�#����ܻ)\�������Ϳ��|E[��4��0Q�_=���@�	-�,��hz[�W7|kO����=.Ӷ�go���x-��8� �U�6��c��޷�;��v�����+��c�aVE^֖����cA�o�,��/1�$����L.��V���5��ٳ�i��-�U|CLpN��	=���Flϋ�G���қGDbAVB*1��n� �ã��a�u�!9ǜ�z�Zm5A�5 �	lE 2���*g?	��m'����F$u?�����b�q-��y$r�J)/UKjݛ气�·��Z(�IC���W�Mĥ-�l!Jiۅ��8$��\����e1��3��_��~�p�}7��a�|��K�j����s��s$�%wt�r�!b5�f�?�!�!�^���E����إ�/K�,�B�.�6��T�Xu.
�er�H��@�^Y�"���d�RR�ڃ 4��[��<���7�|��Ǜ���,���Y�&3���,yw��/n4�X`K�~���,��̿���- k�g�������K0G^���_�^ù�|�D����=�*�$v��q����6\���?.����)<�5:&�$��o��t3���)76,E�t$I[&�M&�5�3��r �;_�[�pąPF�)s�,�T�`]hA�l����2�H�F����uQwn��;¥˪-���i�9�4ح9��{Bb��'H�3}5}��.d�����m������z#��<��d�A�G��ݡ;5�)�&ePt�F��(����̭�����͉U��@SNQ������i)#� ��J/~����H�+ ��v3��#���b��\^�h��z�//8�;���l��%�(Q�>R2\�x�@���7D.11~�;� g��o�f��-���l&2!����섥�Y'O5�`]s�}�6����cw�q�:���w1Fd��d`�=9ǧ�0 Ay��F��������-;�DA3�����E��"Χ{-C5+�e���ŀ���b��߭ː�i8�?9�2��y��m�zc�p<����/�h�
�qr�P?vQC�u�^���� ��`�F��cf�p8
 YӃ�z�Ǡ��xv4 �F�,��$wC/૲j��	�\>��3~R
!��wu{<�K$El��>	k��s���*�u=h�j�l�mBBU-?��G "��F�c�O�������[�Q7b��F��k_�a"������_��YYݻpN�^���T��'��N���?$K��3:k�=�q�\$&X��9�Ð�B��(��(�%I�.���'�0��OPbÈm� ��;%]�:���Ŕf�7b�:.�u΂���N�����f͖��I�:h�1Hk7����7ƭ��~�%+\�C,v��Ħ�*����h��vؐm��Z���Oj�z/~^6��+����P�Q�����c�E�wvN�
�<d�$�	1D텉�rÌ����^~�.�4Q(����K�y���LUn�0^"�Z�Õ�����H�p)�C�j�b�#�`��O\��]�y�fO�e�M�2^����Ĕ��հ<2��[չ������8�X����UBzZ�k��f�&XF�Aأ��S[/�u��@�n�x����btu�#EOk����DKK��3���_{\���TmU;,@�Mh�]��`bN�����ȱ@f�H���J���1CW�຿جvg�CЅ%��h�}��5Sҭ ��͠_�^��r���?�%d5K�������b�T��=J�7�F�����XkZ��깨�������0
�p���U�A���L�ga��|�]}���Ρ�����Y�LVH��d����2MJ!�v2P.`�>��0��q��j����H���z���l�$��?}�:LfUI���l�?� <s?��l��'�?.Ϸ@��R�q��+�hC��a�c
h�қBQ��gX�����!X��*��̖�y���i\Z
����{Z%���g-?�dj<of��^00m{��ֿt�h��}$�*����pMa�)V)m����S��+�]T�oG��(~ms|�����0J6��"�/.C�����|���.�VnUqΦ�_�4�!��<�¬Д%*�T�ZS���:��i	n`k�q-H1h��n+J�7�*�>%U�R�SN�@l�ڞJ�y�Ո����SY�荛�����
2�x���4�!C�	��*T�2�9z�S�z�F��u��CO�,��z�F�O;΂"�D��X�~$�_9ܙ���#�'eZ�p�ϨP��~�k.��"�|�I����i�Є�n�!B��앨�P�^o��"=��!F8����Y���-�Q� ���#�{Q��i��}*X�m�3���l��;���E�ۢ�]3֭����:�'��	��¼����=�9��kr�9�	<���C�Sn~��sl���l@m�~_�n�~�����.?݂�����_(�ЇUt�e���8�B�8u8����X����2��ˋ�*��0���vٿi�� %�n�:�O?r�i�Ϳ>�N�u��R�9�!���P�'�-X��	�˗*Ͳl�t�l��HP�ZĄ��z�z-���Rޗ����b2)�f%bY+U�[71��yĊb-b�9z-�8�+O�X�9�Z����Ã��
��P6���O"ЕV*1�wZ�[�2���>�)uA��_'K�dkYX����4,".su�xV�[�2<�4Ӊ���z���H�魼�AK1g�,����t�K ��E]���)�����e��[���!��,�vΟP���)�-rl5����}&�Jv��Z�dW�����ݱ�{��j�
�[ �����饟 3��f��f�b*�N�u�{�]UE�?]�oS��(���\��H�K�҆�Fq�D|��xٶ����~�u��=dVh�J�7f.z$j�}��br�`��SW{��ٳů���^�3S��\�8X1"Y��'��K
�H�����p�gSr;�|I��E-�pRQ�y#�b3�)����]��vd��u�Ei�OA�����f9OX�D��L:u�v��ȳ�p�S�]� T����Nrb�DE�,��i�Y����Y�_����4��8NϥŻ\nx��>�+�����<4�%�K�"�k�4��K�l[.dC@T$�0��ȫ��߉?el~���2��Ō�O��*
LA��^LI�:�X�	���9��E�h��At�q�K� φ�X3�o�.��ul��Y���ɴ�T�ٚ-�P&��0���=��40���г�J�$���Y�>�$-*��!��^`G�OC����;G��`+Zbs��#{��%��a�n:�v�:�٪TQe�/��/���ya�-b����@˴ �Q@`c����ߨDY�oZ���SUm���;Ցɿ��t�e)mm~W�A���Ƿ4y!������F ��9-�m&��1��SۊBm�0*lN^p���\7i�>҅{8���8�"����$7M���apX�C[������\�J�L��I��IfH��U��d��މ��Ip���s���x���A��%��M�gK�	ܗ9'�fy��=�F_�J0u��;"-�o7�_����g��%����,o�b4ZʴM�h�����@�`h|@��؅��ۂ��Ҡ�\*c�b$+<����������4LȪU�'�X�����K��YVPY��+Y�9��'J��)�7Is=�Df2u60� *���v ���RS�'TH�瀽Z3ޕט���_�5�7�p�5ZR��&���E&�8��/9�MDɄ���L���^5��Ω��1�#K�0�>� V�,�z�T���{��(�ϝ} �]�������K2��Y�c͹ T;���Щ].�y�1�`P������|b��y|��5�0��!�m�W9�?���|��e�鎏R<R{mUs��:?Me���}�nc�jh���*~�*�����&�#	La�޴�u�Ή�?��A��@E/����(��6ŉ��,TT��6�X��	B��U5���rdi��k�Tt�u�RY�u��_�6�I�\��
�:�m38Gs��J)ăN�27��Ԅ�}su�j����1E�nT�d+�mq�Q�ǿ~���{Y~�2�z�v�d-@ς�L�2ɒ@�'�kΝ��s+��p�Ų�V��ˇ)�u��?��)ʴ9����40�㜨�����Rs��{:#J4���w���?���~d_��M��GgH��H��"����|����2��fA�S��=��rmd���^�,��aU�.6��<��3l���r��}�C��[^����EPa�2�k�7�� ��@RKj��}��0g0i���Y���VͶ��E��������E�_�gѪ��s�}F�~$���vJ���Ԥ��f�q�scAF2���n`UW��a�iՆ���b��JjJ�����j[r��/&��c���`�?$uSiU	Qj��ͅ�[�rc��S�.��;z��#z�LÐǿ���d% ��G4�[7�4ZIįD2:L��l���7��
��Tмp7� 'z���c|�W�g��9-���#�'�t+J3$���zQ���pX���"��8_n��\�զ���l�T�H�_�H�q��yd��r�D� D\��\�@�kn9����,�1�*�Yn��U�,<!���Q�Vf�ߗ+���D�k�i.�� �0I��s� ,B\ǔlz������z��CW3�6[ ��x�ؔ���f4��v��߆4��j^�iKo#lv��+�,9�,\W��^(���r_#�nUd�d���#� P9k�9�~�:p�7�����;������V���~cI��},��zMc�3z��ۉ4�/���J�oC����o�XidGd`�G�[i׬1�π<��n���L���L���.[hv}����_���t�o�X�e��.w��d�m�m�;(j�Z���_����m z\>_X����@#���]be�1�p�B|�.�3�x'���>]PE���o	娫�v��U>\б�c[7G?ZɈ�;LJ�4�k�}6jCR�jj��3U�����1��-?�A�s����\�}�r���A�5�����7�ƾ'��<�0�m�N-k ��?�u���.
�}ڕ���UA�B�V1n�3����ǔ>��s��� K����,R��s� ��@� ���Z
2:8�5��/��>*�����Y�w�$R$�7�l�ؠg����4�Z�Eqʘ�I�Q���WH�;�m!U}A|M�t6����nt鲽�����F	�5�|G��Wa%:�����g��;f�Y3^���<��-��`Δ#�9��%��n.�+KF4&���E�*�7Jgu���
Y�)(nB-���ms�O0�#������E1Y^2�R�s���q_�|�X�!�<t�[*���ѥ��=�_����R3y�g�܎ʠ��B�LN �X���ՌfL�xao��?�_��{�s� 
��)5�R����&r��*p{��I&_i%����f��=Tx��R�����Q��K:�Ǘc!�܆������IU��?֒�g&�����~d6C�;����b*��6t�*z�u���U�7�)��=�^�;��ar�ߜ/�契�[J��L�ލq���f��O��on�@�MF�ؕ��;�v휬H ��L��=ȱ\
T��c�}���5���0J������Lk��Ѹ#k��t���H�)�41O�'��4�n[�d}`��%�Դ!Վ΍�}M6�����Wk(_Cgԍm8�u���~q� ��E'���w��"s���ܳZ����d���`[���6-8���Q7 �3���X�N���'A�F�3ˎf��	�.���Zy����'�CA���[:�ä����`�����4��bjAH�xx����Y0�.⇡��N�w��ȺRz�3댵�m��o�H+CmK�7Q���ґW#ʐ/:?7��%� ��?���~�7��?�et8'���*��"a*��I�޶��sM6@��w���|!Cn���9N#��5�T[�/%!Ky-+�Cym���2�m�ʖ>�*
���I���R?k�=��`=��ܿ�������1�t�DZ��CG
%�3ÉsJ-@�n��~�}�xR��8�|�:�������`z_��WhS�|�oG��K�2��P�/���N��f{"9�����q��\�I��+A9���f%x�/�h���M��N�.^0^�&�')1�)�;CksBk����\�Uo鹉M�ςie�/�˫��/
�/��Ꮻ�'���m��<���>�:U�U?V��SB�'LD��)���R����6�7<F��(v�*;� �K�)%��͑Ti �^�l�e�%ޖm3�g�e���@v��2p��*}T��0O:��<��!K!��<��+<�*Lb��֨=_16�ć(h��{6����k�"�e���+|.	�u�
�}ȭ~������Ib~ ��qfVk��ǟ]B�,��kV)8j�lznn*K�4U�
�l�_�9�f��#=QB$�_'�]�,�E�d��`@���#�;؇>�R����Rj��x2�EMI8���s:��*��ܗ��F��A�`��7p����T���
�����0�c��S
Sc�l]m.�.�^��������	������L>�[�in'����y���Q�D3����(됑<af?�0����V��y`Q�b� �L�n[�W��e���|*��7�S,0q��C�A�0�w	|�(���ͬM��Q����9O-/&<�˗��GD�n�w�Ѧ��;���krvy�$/8�B�����+�j�JV��ZC����ř���	���OUtk��П�Ւ&)�m�@� [�YƎf���=s��P���iţm��Okf����R�Mv�8����9���],��]�Q�O�?�,|�udk�±��=��د�T������?C+ɬj�q�ͩE�����Cr 9*�B�K~�G�<�8J��Z�I�T}ߢ�"�����*=́6!"j�B/��=�z�>jo��_Q(;*��NE�Plp�#�Bg�p.��i�t��-�YP�ء�>���~���!�ؕ-A����z��4n�KBhE�Th������Tݚoj��s�&{�/Duz0���~��K��#[���g��#�&wvY��d�%) �i	
�њ���kʗ�M*`7��@#�Ι7M ����Ơ�ɉ��V�������@�I|^��M<>.�U�!�Ph�9�,9�@���jդQS(l�g?�l�^��g�Lz>�'��gk�C���N��g'�u��
c��>�M��]�{�6�;���E�L}1I,�X�C3t�I܏}&+��,�u.(�$���ԋ*Bѻg�_n���3�u�{Xc���'��X���|�=�0�� �RA�zGx�����+}"�<�5.)��*i�㍼��?�m�E�v�$��I-����e�Kfa��a��8t40pi;MS%-�s˴	}oUʊF�QD{�tDu�1F��o:�#qH�	��O�:h�a�W�v�R5T�ݯ��\}$|qҢqX���~)� �eDU��\)z��Q�:���9�%���*5c��o2=g4����
wǄ���j�A�|�U8�m��ݜ�B�|�Yӑ�X~g�U�1����<7Wj��YFjf�/�����'z���CXΎP�n$sO�U���X(�7�f��չa��a�K��,nb�����:`���m��Î��ٲ�^�i�͚AP�NFY�Y"qK�iC*��N6&�f���O�Z�0~���%�%���^���#�lna�x#L~�����@IA\$�(�����Y�^<�7���5[�?�{1�R3(Hώ�̃��K����y�sܤu5�����+��0�Ph��/���s����:�I0�����$C���[g
���E��˞�/2;����&������|t�������f.u	5�t��b��c�@}���AVF�lQ�bܢt�1�\#*#����E�D��H3��e�B���@��@�&4�Sӵ�N�o|"\JV�k�5+���_D�4��ț�ce��� �%RO@�I�!�xtZ*�6�7f��h��u�enQ�	Y��k��ЭX�{�����4�f��՝��2�� _Ths�{:��&�P�̼����T��^a*T�jt܎ ȯ����l��Ҍ�ÀkZ��Cmt ��/0��l�W�]�����P�0��lR�Jǰ�V�ǫ�w�e߶�j���q)l�fZ%0W{���I�}\�I\ϊ	������K�6��g��0'���5�e�߽�:�2}�V�>�����mr�֘%޸��q���u��۳K��57��4��I�Рi�@#�pI���<by���ҿ�󗨤neJ���e�i�q:�Q����G R�<S�h��R5��i�#���"�ϑ�E���7:D
�MY.Vc����S`���]��w�vH>�C?��Ử�yY�X�� �Nt�����3�k�Վ7`��'��P��)	�W���/?�3]0G<�,q2�,â���-]x�� G!>�����O
:��.�����g���RF"���7�<.y�BpF�h�+��n�ئD��DxO�>�΁�:�$��O2N(F
�6F�ڀC.s:�(0f�1��F%���BV�m$H��cƤ�B�6V?T�������\F��դ{0�����'7��6��zZ���N$s�|t����W9L��4/y����pq<];����V�E�׻x&/��K��w�>����)^����M$��`v�:'�f7�
�H�\��[�����|���,ļ(�S���enj��A�I�w�F�+M��ޑZz�E#��O�lٜfVi5: 
T/��M-����i�}�X��P}^���5�[���,�0��k��G�D�W��h����9��۞�{��aUT��K�6�O�I��h��Vo�P`�꫞8UK64���;E�\-2�=����-�W4�3舦����u=��������3��<�|��}������K�a.�\�/h(�-�����a@�A�ި���RͰс3Ȱe*�L=tб�E���z�����ק��x��̘��U(p�iۚ)�}P��o�+ULK�9���DtӦ����I�ʟ֪a��c S�P޻��ĩ�&-�����<c���0$6?q���!"�t�goM��}����:�X�$��?�
A&'�N�`�;e~��R�^`N��˥���o�Djhm.��i��]�uz>�)"/.H��$��wta|�L���)-Rlj��� �%:�Q=~j�0�^K߂J:�!J3�7.HyD#�%u5/I��a�����c%)>�g������	4Du���(8za��LjA?E�`E��(�r�Aa��O�>��{¥R�����Vo4����9Wy�d@w#�S�A��W�\�4T$�HG�R�u�e�N58:ˮ�:*0�j�r�}�Yt����k�{�q��r PР�<�򬴓��̵��Ǘm_^�'p?�̞�tn1=���p���+����
g�I�D�f�[B�4�8:9�9��\��fv�]�9Py�%�5v����觞�x��b�-�sa�$&��q��P�^f*)*�;��_��3꫸�?Л����}��.>�-I��\�y�4�����S�� X5g�]�n9��z�����x�������o�᎕�}d���\�G��s�b�M�u����%Ǆp�]�2W�%�#�=�Ǵ�g��j���܋��Y�iй��/'4A,��7Z�>��l
/��0ӆ��UIϑ�`0�l���vG���V"��� R}z��kV����)G�G �����[�d/�1�O	�dXE.�)�6Dat���_�ى��:���ξ�y�K����U�݅�ćc���]�9��-�L��@#�n�+�GJ�XH�	��������>�F��<g�%\�����m��������g�vI(}E[Ɣpn{$eq�	&iQ����u+��x��g�"�����-�ΖYUIwľ�v��s&����@6h��1�Q��k�>-�AS�y�i*�H+�����_��Q�-)��+�,x��;���|�O�植�qhkgås��C�c�-+Zx��/�ӫ�e��O���$!�)0P%`����9�\�~f!�N���vA�b���!ʜ�Ϣ�Ч��Po �/��٤w��/I��������"d.M�:��隣(�����NI��Gn)�A�WE.\����G* ��V螳�Pv+��{	YuI���R��.(l_j�>2x��%H;)H
��5�R�7-����rs�XR�n��t�����ll��������s��-�8�M��V�3�a��m[�#��z��K�X�s��Ev�ۃZh��tW��f����fe�do$ݠ�}ڪ�ZG
���N�bи��7�Y��ISo�6�u^\�0�R|p҈gk��E�x�2��~x���$B˵�8/�p�?�v*�~�~Ta4
x�[/�s��Iw�����x�A�O��|Xx����4�;�!��<��N�(�\��z��LMwt�\�;�T򪟙�$~�홹t�`�|>����(�� ���A͔_W��$u�D!�w*8R?I@�T�ކ
�e�v9)�ܷ�vWA�_�,~R��L��>v*����M\��!1����C-ԺZ��9����1\i�X�m��Tkh��1�?$�i���3d��A�=�O�9�}�NH��q��I��pF���6�����qq}M���'x*�#L�'�C�&[x_�O�$ҕʨa�x�튻��Il�	������
��i�s?��4{�O��hϴ���pb�4�oȿq�c�'��9H��M(dJ��u�[[��9��#�f��Ǽ����q�1�VO:Ce�l��[IS2��H�5�
w�>�h��ӛrpx�I���Qn�5[���~. ղ,�\���{�dcI��[�-�G)��}ᶻ�g{i͚���'�mE�	�$3�����b�Zhx����B}]��*^|��.�g6��F��od��)�d-����8�9�go�� ƪ	Z�Nhɇ2d�k�.�V���3s��x�x���ƲL��7���U�
x��WT�h"��v�\����jz*��BHjՃۮ����.oqEs$Q��b�>�V%��"J��n���~�F�W�=u��9(2��1>d��|�R#Aup��D�N(��WW�<��)�G#�3}�?��y|xRㅊ�܅p"E?N�x�������	���]Op�T��~��l��+9iw��OY]q�1:�C,M�����0ު�ī�t��v��V>6����Q4C"����yHd4�O�&�m�nb6��!�]Y��������uq��:�%M��e��!惘z3l�غ�|rpn�٣��M�����?�e��%�uY��r)m,�YJ�M�X��Og�5��:���?�㐧�㑧2�`��/
��L�yYJ+<���&��B��+uQ6�P�n�`K�(bOuؙ�FN3E����?��`�.݋ }:��fs}}~
�����fJ{�m�](�mi� �ei?�+��1�O���u�{2�T���җ�ɯd�=��GF���/��R@t�Hg����N`b׍Q���X�7]�Cn��S4��
zXd>��PY�ua,:WmZ6���˿;|x]�4�bz7`b�r%ӡJ��\\��(<�>�OT�ߊg9�Ӣ ]��C��	���跬�>��:Oc�]��3����&�kZ� �]�KE],��pA�+��[���EF&��߃���,]!�.oMҡ��r e�FF�'Z���
�շ�f���܉#9���E$VsL��[0��.<�B/�
!����d�φ	hFG�ߠ�M]�z���mU|V�X\���~K[�F�-�����'[+l���mu+����r��0PZB!���4�z����?�$m����@�8e�@�L#c�3����R����]4�"P��{���mH>����>kW#�ܪ�y��2ry�-:Ü�[�ڽ����P��3r�<Y�cmMz����&J�����-��z~�C��3�����ܬ
�iY��p��ょ���߀Ϝ�u��.7�t���hO�,ʘ�g�)u���<�=���O��h��:S?,�*i�ե���a����~����s�2m���x���#��D;g͛xrz����]8��<z%?#c���"��/Mju�"2��널���S٩���5k�*��a_8m�F!9z�3���C��q"b�����g�5���r�v��,T�����^h�2�:�X̥!��A��;o�R /J�e�{ү1;*D�_�ÕK�NP70�ٝ�c�i���p ������	��-u�����2PT�X�bkg����,z�⁉�2�E��Hs���Ĉp��D�� '�%��_�0̠��5'й�:��H\�V�����qh�P��T�rE,j�_sP0�n���!�B���޴!����eG+r�8&\��Z&U{�� �.9;V��N/���nY�;�j	���L�\Fq������W�������#��i��:u���#D��:TH�sO��N�Ҫ�ޟ���O��4�sP����A0�tuY.˖���n�w8F����_�kc�+9q����њ�j��:d0S����;��M�eE�����]�g^g{͇Ŗ�WW0���\���.KE�[���?�{0b$n�j��2k[�I�A'�Z��%-��(�.Y�A��*�RU��[��{6¦L1"��Ln�0r ���h|��AxuH%��?*��ބŸ6	�k��� 6��x�W�a��B�K���,�����]���=�[��6�!rT���kh�
�f\�Ϩ����k�bZF���������Sx�^�6c�;�i �2�oa����9�#�B0��?t��~̢4����ݙ~��7y�Ny*���
���q��f�˞�#�nY��Y��׌s������ӊ��rm"`P|�8K����8F��{��z1�Ւ�\�RSJÑ@'�ca�6�_j��k�:Ew��;�藛�#ٖ>�s��[���%}>Q�,�ā6fn����dk>�3��bD�z4�,|/0F<��ʹ�w ��7�}v��K�Erݜ1Ū!LZN�+��[�2����p�" b��,�A*�j��� Fo�������5�jE�-�#$��u�f�g|Z�u$�:ݵ��>�ҍ��$,r���kR�3�՛�2oqY�#��9*s;��xv���3S8��GB����q�!�z;�$"�f`��mE��G>���S��
)����Bq3�I����~v��@Bׁ������.���p�����0rwf.��qܼ4�D�����EX�ɸ�PG��ٿ,���,Xx��˚�Ff�*����o�
&q���\�n}:K]<(5Z�6$8�b�h�*��-
�(�� �ͦ���-$h~���m����gw����b����DZ��\0a�8�3J%D�_�����TuΖ^����1ج�m��P��~��Д«����ڇ��m,m8<��GudM����:�c����J�>���ҁ)�N���&��J���
���� �U��wcuԮטw�6�w��.|����q��r�{w�i1�����:���w��9#�#�;9��62��H�!���3ǰ��xs�t����r�#{�\��E��H^��|r��4u�=���̗��h����G���2
�����@��ڡ����t"w֜��â�o���C�Ól*P�ޡ9�"P+{�:&Q#�I�4:OGU�bmd]�GH+�8��3�;��R��#�O���������F}�����������U���G���E�3��<���Uer�HSN"�@���D�X�����H�l�ꒄL�컌�ȏ�*����=][d�@�~&���o{��|�Y�}is�<ø�6L�M���V���	�g���i9Q��b	s���A./PB�������0����� �Xn�%_���G�J:X�t�"rz��p-3�aK�����E3M��?tR���zE�	w�ּ��5�+EEnqS�T}�<�=��͡� ��/��>�U�1/���>H�JW8����Ҁj�7_��O,^���Ǳb�W=��-��!�{���:5b��
�s��3/� ��YGc�p�Q|?؄��JбØ��m�����J�����Y�c��-�_d�'�z�k�ׂjo��`�7���+�����D� �Q���7x��Ft��*����?�g4~�/~j&�K/���,(���Z�'�yTtV�Hȯe��]�?�f��$���]jj��3IL_0ᑔ�l�y�E�����4����dވh�'$�o~w���������E'�E����;��ұ����J�j��,P�����o���;�����|���,[��T�:��)9Q�9�icY>v�Y�R)i3��>��m?��*rp`��g�����ZoSN���XJ�Y�+R��Ke��|�2D5 �7�����IOr�ٵ��N��N��V}�s�q�87�˵M!�XKЎ��+j�*Tɏ�x�03<���H:J5��,<�6���i6`�k�^���.��F1K���/]��lgߒa�"G@S�s�[j��Ae��N�Y��&c������#��&%/�\�yy�Ǒ��v��ҫ:�0�8�pNd�j�됖j���J%�-9p�Ȥ�*C^C�G�.)!�΋×L�4�ո=2 f#�d�|��H,_��aiQ�FY���A�+�C{ٞ�k<Gj��� ����M��ۻ��M��.�yO�����F���&�318t��CZ�%~���]$��`�D5�����G�r�珫��-�P0(���!�bZ�EoU�Uj�Z`Q��JpݠV��H���24��/C�6�'�(>�쨀n��3Cl���m�p
۽��K�X�v�tp�n:=`�tO)����[.%�ͺ0�f�3 
M��}�s
,�&���n�N0�>([����,k���5��?�U'3wT��É[���H|7ǯ�4�S�>��-��SpMxAX��z��/&��v��~ְq�|tI�?|8U��,��=ŝ����1�\
XK<L�L�A�%�:_ ���ca�'"!G`zܥm������?���J-�Rɸ���b��U~?�,�}c�Ʉ�ݖ[�#�s����l���NN�ң��y U��%7��b$��>"�w��^_y�.Db)e;���[�2�x;rX\2\���/5�C�=�H6�sl |d��>y���K�������,T. ���'�(����E{���4m�F�s��5�N��a�&v�d}ef9��,��]�@E9�ɲG1S�;��LD[	�D2�Y���z����L0�t��-6�𝨀�=��*�#�I��aj�w%��`��h�^�|�	�=a���9���g}���t[������"�l��U7����j���jB�áRz��� QFىYw�FN�/U��w���Yy������3@�O*�lT���>'�u�hGظ̕��yo�R/D�QQcDĖS>:��a�#T�YW�F��7gP㋙��4���U��R�Sv�W���~��?YqPd���$�cB��p��-s��KK��;��$5!g�J��pb�.��wE��T�A�|���y�0�O��*;ez�+���m�Uo@%0��sXݺ�S�ex:Q�R�A���6�|ͽ�&�U��T�'��W)4%�$L�O-��_���\i5x��� 2�8��ID�����QB�o�;1�K?�YZȑ�T��;��sU��8�{��s��.�Μ�l��q3�o<�Y-?�	Jb:I���{�(YXgK�2�;cG��U�� �G/��L�I�W�J��2���]�_���,�r2�RA��JA�i%a���X�Z��z��4������V���1`N_^�*��T�j��C��{U��~��.e�8��̸�r��H.�B{_��މ�B��c���+������wv�Ꮹ����%M��w:�&۾���|&�e�i����Ƅ����,]�Du7/{�� ����Cv7_{be��]�r�#�x���4�6*KR�DU�l$��27�3�O&��Ϊ�92���9k=�6�A>1�֓�рk��[��� �v*��V��C�����s���ҭ�d�A�8?�a���O����{eN�|SS�7n�{7����x��1=�,�k���JN�T!.*��F�*6^2J�^�[��;�����a���	J�u��%v5�h)����W� 5�s�mP�Z���.2�P-
OM�3mk�'pCQU���_�<H(�y�8�J�O{ǐ�q7�D�V��o;�Ov�d�;o��<9���Q"#u)<u�b��KjԗМ;ƽ�;x�aA��`�EK�ʶ&�wWVl�*�W4g��de,��)?^=�H��N�"�M;p ��d
)��?�� :e���fx��h������=G�Ֆ϶?og@O��ns��	��tj�܉T��r��g*�_��ʯز����<n�'tv}�w��N,����&`Ǩ���Rl눀鞧���h�|&C�d}�����3�2��3�9��W��&z��u(L���=_e�<&���WdB�K?�9
z�	3inAa6�|�C"�*^����S�$]J�g��e����n2�ʣ��R
��x�Z�e��$���"���ר�#��٦)�F����h�o���0�:;�{`o~u�T@u}��>�*��r`%mG�u�zq� �}'�k{��C�2�y(�])����B*[(�̽�� �˺Bǩ����	���)(�4�����@c���j�]�T>�6W���1�X���H�_�PK�Xa��;P$�9T�Z�]{9�T�Y�9���
z�DUC�*��}�w\���a��b��z4^�z��zI�w���3+ �	�{4�䛼,�X��IfD x��8T;Te-�Nd�=<5���1���	3�++�k�]D<��^m��jv�s.׳���ި�WD���f��/UWTd�n�C�M��r.�2>{2����հ�&�+�^:LJ��ȣ�dY�Э�cNr�wY��C>L�8Q�H�R�P��TJ`���d&d4(3��í�U{��(�)�*�Yo����>����54����3��l�6c�,�Ś("]���	I��Et����g�s[īl�uɢ���o\��嗲.ff���c����Z|�.J��}4��gO(�o30w�1,�������͕�-7|ăDn�s"XaǰP(�� ��x~`��x��7�5�[hؾ�°DA���D��0�s?�gC�Xއ�D�dZ��4�9Ίk�&i|��a�,$�<�� P8�¾S��`iT��T��Kş԰ر<����&��/�ĚI�VG��o}X�{4]W����r..�p�^wg��d��H~PYw�Nc:��)��e��wd�D|�D.��#�3�o�ts�6Zsَzo��b#�{V{!U�(w�^NU}hm[(Ⱥ%1��W����%dХ7!�]il��" �zآ��C���8�u���J˞�n�6�ҷe�:�-L�,�Wkr'h��]���T[4kւ
��)���kiI�S��P�����i��c�t�X�дA�u�v�>��?��Ӿ�׷����ҾEE_�yY�.��#�x@Hw�Zk�c����O؛Q$�������R�m�CS����HR|��%�|$<�H��E�9F�/��[�m��g�壢�Oյ�lV���գt��S� �G�wb�-�@Kf�-�k�:�S�@Dju"����|t�<�@Y�l�qX8tns몜}��O�j��'(�"���r�N(�]�WV\��� &�ץ(�^M\�3���n+!tK���E3��8~y��Z�v�q���������3K�p$��2�����A�R��� Мcbk�8�i�8��uz��_���(��|�����TJ��Jt/��)��T*��6�������U��U���@�
��mrK�I�$��y1��i&MR�.��g����~@��T�:D�r��V�F�
iL��|Yz6�,#�o�^��&�nC���D�e�B�=~5/ƭ 6�$jwxW������ O�ڳ���rС�-@��}�^����}�+�Bk�6�tی���U�&`��O��FQ����f����M��t5�KA;	[Z��y-����0�Z6Ҕ��p5��mEp��O�$���,>�yt�1]S���W��U��gKG:5mqɦ�{h+�vo_�2��|���O��e���>,�v�T��"=yz�A+9_K�+'0ȴJ$s��\a�E�<��.��,ä�Z.������*,�e���U��A��G���OJ�lQB�����M�q�8����l<���;�������y�R�l,n��o��j��5��G g	W�"�7(>�M�!��y2�L��Q�n�p1`�btShI�!Y]5�>F�
����'km�UG�׈<V�̜f�]>�b>���xG"*�XpЃ3�,�u�Rޠ�s�� ��5~K��"s�_�B&�XL��f�9���>�Vĩ/H�M	e�m.�ʧ��^J��fp��"h#��#M7��NH�ߪ��!Xh;n_I��X?Z����RD���B�42P&7S�/�j��5�T&�����RI��d��:�E��V#��dþ����Da�Y��A�0��_��4:��h�Ŀ���q�X7Ms^����=hm���3(�n��'G����l<&�zF�R��vuز�P���3��'��?Z�5� ���A�s
�;�9�uY��9�_��M��y� ��<�S��sOw���Ռ� �"��Z)F�Z?:��c��2�m�[��VA��"��Y2R{W�~{~�>k��>i�qg�i�V���}=�����2E�����o���crdc,����L��h%\H���m�2'Q��yE"U�����
���E��� ߗ
'C�2ޟ��gQ�O/6��q�aytR�I��i�Єe���:m��L��������卒�I���R��L8>O~���jӷ���)����*�<,�5�բg��vo���fs��L������As�2�C��\�}�s��:6m�/V�q�;©��O����E!��k�����=����1��C�����wX9�W�X[�*����ݔԼ<����i� ���7r'�<m��L��	�c+��##-��%���M�J� �ʇ���,GV�?/(�X<��d�@����5��h"����46��5_��?s$��֩X"�:�y�0�Lytֽ�	�k�F|��%�����~�R��av�ir�j�E���0���YB9)x�ǣf D��<���G��/Ԁ^͍M����2�9��~����&��6���5�Y�!!��΢C{��K�sO���O-�:����c�*��aM��p'�|���3T.�����F�pRū�4C3o�G�ĭ���ۭ��M!�V��1՚40�W�*�|+��A���a|CuSO9��"M07FC�0�t�(Hr�Ni�"h�2rҌ��`�p��pm���'���El����P���%�'5�'Өq�g�`6��S�^/Vjnzs�*H��	�q �O�v���ڑMn�gR���!LX�,�?�]N�[���
R�%��D������A�d���:h/�Wv,ɲf#.��˭gh�GfK�fh�;��� ���u��	����[�~�0G������0�\p�b������|�	((���=&�>����G��i#%/����p���WW!�
�{�Ïa*f:Rbqq��ͽ�Vγmc��L�k���^��u-��l"�����{h�����x؟���\�BK�8���@�a^T�b%e���ٹ�֨;��3����q\PJ�ܱ��\'�c�=�@���W�'���ϰ��%B�r�~��"����r��^w��i�;��ٮ�&�D!��J{�ˍ�1}���q�xt�GdE��c�G4Q~H���~\(Q�S��4�x�ekrB�O��+�3r;^�T�6_��#��ko�z�K���3alϠ �Fl�*}W�C���M�nO�Hi�7�%�<���T��3��s0��'$���b��B��Y\��4��/�y�T�R�W!Dy�X��g�rq�Ai��'�-�����[��vf��@��S��ls��M�͵3�#*}+��'���ި��ƭ�	4L�q��D�j0ذ���b�"���a��Q-WG�^J�Ͳ�ř�B�b\Ug(��fEhh�m�Y��&,��\�$0�t/�L�Xu�5��9�>= r��ٺ�<ag�b^�W˿<��r%�K�]���&�z����!:V24E��O�[*��~�cw5�>u'����N��v+�Ew��Ċ�Y�y"r֩��M����
��ܯs?�e%�: ˂�����G'�"�9ɳ� �Q��K�?]��D Bx ��C�ڗB��T������Wv9��ѓx��'F���K���Ԋ�Fb��>����RL1��꣦���-˱J1h��m
J(��(h���%�j�/n65ǡTG"�Z[fQLw�QF�Bd�@>��?(�D͉)��"� n�D/
ܭp��;x��D���Rt�(������H���G�3q(��)|����%Am���\���q�aH+a�����-�?�L�lޡmyZ��"�%!2\V�ҘZ�>��x�#<go��d^��S�ݔ��T�08����fƘ@s+�k�3I��D8�U�O��G����t8�0�o�J��[��3�<fղ�?���B��M��E���?}��q�p��;�9D�8��Z�ް$U��7��0<�94��X/����g�7Q�(K�&ރ�)6�V��1��8����$6Ǝ���Yz߮Uz��0���܄�e�h��DjŲ�0�n?�Pd�w9�8�g���)��N�K<��������Nm��(`���C�G�]H���}U/��%�4O��g�>���#a`A��'4�!�4D4L��}i�DX����5�Fe�5��N�q�jm
$Z���ޜ�U��"M?�%W��[���a����qS�w&c��楸�\+G.V����OpW��8Sl��9���A#�z��M}N�⮈�khz�U}�$����`;��%y�Tzq���������b�Wy
����<\�{,�í����{V��$���U8�tk �hR�h��^�fU">ܣ�[#'��i4]����}z�;�'r��]�qWQ��2x��9o��B���`wu�#��`��`��RN�G2�£"�z���Ch��J\��g���Zrk��co*�CQG�{�5��9���N5G�N�ܒc�"�y�ɳ&�iYnY�[���f����R�x�)T̋i���JIʊ�5�M�Ip�oo�p�P�R�~I�&�]� 7�h�X�:��-H-�h� ����=�3�T�-UJ�C핱�㺋[���<���MpidSY��=��c7�f�5ѱ��i+�69�Kŧ
��ovߍ�+E�r�2I��4�'��ٶeT��|>��6�o<̌q��� ��s�!��K��߂�z"E�)�[IF�+a��q���7t���P" s����x��+�Z���c.k�����y���6�u7JF�ٿ�@Y��c�}�!':7�l�3Wc���lhZ�K�6\�uc��v\�M��`���Z�*#�NYo��V��E�JN���Q�����֕}�C������]�3>�&z���$��/1~M�� ���Y��� �)����&��
(�
�������������Ŀ: P��ʃH�G<��9�y�S����1^�$5?����t�w��1"OPL^�!*r����t�~��b�4���e�w8_^��d4�]C��Y��E
0x8�Lz�����8or���%GǇ��<��J�.��Aal>yz��T��&Y� U�:B%[i����}����4;M���@����]��v���;W��<�f�?ru��rJ���6q!ѝ`�����
xR�
0qP|���W�ʽq�+�Ө�&F�rE�5	���i��g�&�a�VF�T��	�.�n�������X��Nn�%���Lxf�$���~/pMEE��OVk�\΅"����i].�:��p}�g�Y�Ojc�lh�@� �E���4�|��UyU�1>?�@�?\��3���A<B1j�F�ڙ��g��Aj��H�9z���+zeul���Nb�>Xx��= 8*�\k�F��1F���	�Q�dH�:�$�ϱjo��U״�cu&"��m��HI���w����B��;�4:�|�*@�T[�D���԰\�{yJ|C��VG���sxX���\�#�r�B�IQ�V!z��@H��Q�Fqf��n��1,4����=�)�PMЅ�H�pd��V��n%�>��"��y���t��W���R�E(�Ò�@.m/��QT�sFs7X1�S哖�����(��a�+\�+��G��%��:f����Y��C�	گ���V��d�u~���%�N��c/���r_^��?jX���#�w�R�];��R��_�:`��,��Ϯ��,Uo-���̪�e�ߋ]�5C��,�����<a�B5��2�r�������]�Bz�S�F�����9��䚭�ScH����o��:`B>�����ߠ�O"�K�+}g��t.��:+%�,]�|1Vm4��|����������*���i�6�皢���T��WQm��(K�ٵ�k����2�·���������b��TK�����z's�T�|#*|i��ӤG{���LD�^N;��*�2���⸾�$
ל��47C�{�?��?�����[�0}YĘ���=��)г�HܮW��}Ug���V\����T������K��I�)� ����p!�W���W�5�L�Hj�K�4䆆�8FqG�
yfpK�6-n�f{�;�Y{�62~�&_!L+���l"�����h�}��P�l_2=��v�bC����AFliWJ-��I �ԞC��mmm�� �Jzϩ��:�њ�,n�kQ�3Y��?wɆ�	�0��W�b�%Zu����5���]�o�e�A��Y���b>X߆�v��u|([~���8�M�Bq�-�T��9B>K��	wr�<�n�%��I�E��GY�⬔�+@��kF��<���dq���+
�0�pO�#�S�]�9.�#w(�U���/{yG�k������q$`��,o�V-\��>$,c��h��2�F��)epd#��.�������s��*�]5?�<�$)-���ʳE۹p�L~4 �GdG��w�1��,�yG�N�糡B���������������0�{*��yL
}�M�ֱ����o���U`�ݫM�;���LVD6i��K���=���b�I�wudLiM�����3y�x��TF���Q��3��"A�mG3�l��k�F�R(F���B�=��� ���o����!�9��sc�6zP� ���H9r/�1jb��l�9�o?��pfL?_��̢�ݤ��L�#�)�Z�ث
���	M����t0��+8��h���Y��'n@��)���sbv���ФWa�*o�F�Q���f�8)��6��*!��Sp꣢!�e�އ�?��V-�@l�6�f#g(/?��j<	uu &E���eV���MZ�,�R���J2�u���r����!��r��D�p��K,�a>�~��C<S��'tM��9�~��d�n-%���.!�mzu��P��M�5WJ��7��ڗG~7�+7s��@������^?�`^UE����	��s���G�{�VK7�sF�%ozf9؏��ϧ��x
���_z<�m�8���3��9H����i��=��֡  ��ڀu��Hq0���YH;Gy�� �l"��a
���$3]fV��j��B�2g:0XW��p�F���zHP�v�6��G�u���OI�G����&�?@�0�<;�Lq$0�I�o:\J���fe���JP�wn_I��t�Mc�T)ެ^�s�+T����]�
yeD���{���i�?�ο�Lc�6����޺E���P�P �'��~�5�Uܬ����ht}l��RC���*&îr�����[q� �k�V�	�Q� j��ԑ�D���+�%&�� F��yJUX�-��
�]���/�V��
�\ �E�L�	��1�SfI:Ai;�kOc�V���O�!�q�`ٽ۠�L
�o�EQs�ur��G�t�y��z��-s4�dmX&��Ay8'�4؉��@иr��П!Rf�{>`?�a-�oD�~�E�/��T�`�2gX��d8A2&i�����G�Lے�Ы�Y/�WǴ�yn���!P/.�A"E*�9�v�g�q���x�U�*>.�V�5���M[0 ��AP�ԀVE�љ��z��+����/�G����x�Z�F��~[Z�����QR*�s���xjډ���J�~P��s
�sR'��'8��|�]%*��R���B3�gĤ�/�dw/WS�J��:+�<9 �U �D��$QܱjD��W��H��hs��p�΃�\��v���q� ��y�<�("�.	0��LEj�ZZ�ۻahp �0 m����``�	������v�~xL �dAw�=�Qo�t;L�aR����W(�ēh#ȷ���<g�K�!�ڛn�\q��#v�����kw��R��&�g�E���,��Cv&�G��Zo>@��i����ni��ׂʵ��Ԉ�7z4�Q0�_��9翽��'�����߳r�*/穜|r�
�NN�vKQ� �:���F�S:x�3�T��~ˤ�	��y�9�$y�%*;p�c��;�DV�%����G��W�s� ��~f���BU�	 ���U1kb��.���/����3ְ*�M||��F����[��.@��˧��黱�s���'zWґ���S;�8��3_���/1vkK�1N`E&�6��[:�,B��*��+d�s���W�X�e�IQ52~�[u�d�*�ɞ�4���!͕��)ڼ�Jnv-��iR_3��O��jW���$�\�wΛ���V�ж?���6����)�	��	Xe__����X��|0��Ē�������6g%}���$��������>���A��IJ�2SE%�w]X����[V�˓��-�|��Oh����nR �G�|�LH��-ߨ�܄y􀑆X@#Dx��0L�@o!��$�fTB+�����Rl��j�*2S�<(�$����߆m�ߺ
�����(���uՏ2�p`�yc���p�_�e   cJ�G[�)�mq��N����t[���3؝���(���[jc�E��j^϶���{�be�Y�}�f�n�%��ɲ}(#���#�fv��^B[8�3Z�����ϝ���/dK�c���ON�Y���yJbQ���X����JaȒY�ln*�k_'������)<�V��9ɂ�$�o��|�5�ا�.�_�o�mĖ&J����s2#
C���������V@Qu�$� ,���O�&��p����-�jխ����e&&*�ƙ\��lG�3�x���A��"�u�?��k�%_%�@Sds����e����=ʋ�?<�H�0�C(�J+���#�(�	�Q�I�U�V슩MІ1�%у
�Y���V�$YL>��0E���Uj��cșp¼���.{���V+F�Q"��kʻ�A�$*��JH���+�Uk����hZ�~��è��L�-�d�B"�����@�������fڲNd�p��0:a>�.�o>��ρR��hF+�/�U���GI2��+��x,�����+��.�įZ��,�3���T���KK@9j|�}�%c��&�9���������1�R���,�T]���XFF�5E�YA^R.}�����J�ĩ,����ɓb�V�p*y�����+V�A|��1fdr��wY,�ě"W�h,��b<�Yu���72�^�z?k���[��7�V�0)|������7ʦ��z@1�Nr/.�����E�cJ"};w�O�8�3�������[�,p��}���J�)���AD<�5i�����~��gUt�F�����c�M�QH��2�ˢ��1�B�T���?�~W@�]qz�ʺ3�ѕnPr��HS��C�	��R}m�)ۄ��u�Љц��B�IeHc}��ݰˇ�#�7V)ÜVPB[�(�G��(6�A/�V��X���o���3���zmg�D
%�4Lv�=�دċք����bH`�%MXM��D�;=��gy.�JUA:�gW��g-㱙�ZE8}�������##[��^��[FI0�V�:�Am8�H8���)��_G����hf]K�jl�<���&Ez�x*�-��y���</
�O�ah.9m.��o���L�^�z�!��T�j���9�r�E-ϻ��?�B9��DQ�+H��( �����D�;�S�>�TG<84g"�˦�q]�k�~���S(j��0�L��4�]��͖mw���RT��̻&al=t�>Pya�y�g9��@��z<\���G�/��0�L�Yb�:���_��1T�����y�6v��yY
}p�R��cZ�yoqc��t$��3���S����4JQ�Tf�m��jdW!�@��_`�$�#�Dx�ӥR�p�eb��:���Z�Ӛ�~���h��́x�J���,�eY��{'���*�}�='�LˀY�wSy���¼�JV�wT2�Co��R�����Sg����H��y�\��U[����~�˫���3ar��g)��ML��d����Q]���I4i����$�k�%f��-��G�vx�@V����]����'7#^���|I�q��ql�;���q#��i��������	\�&�B�M�C!}�T$����'ՈoUU��=����2��C�R� ՇJ(�O��hG����$�.�!b�!P��|t�}$Y�pXBe�|���y�%�2�û�U���6S���exر��Ô\�>X�᠝ۘ����~�z>��~��
���)iz�U��Y���D���%#�ߟQC�NNq�;/WB�{��#:LZ����;�1w�ɆS�ܺF���[����[�Xc�Rx�_n��|��Z�/d�Od,�X�ˮ��[̮��E�}g��;������0���Q{�<�-�6�|\�T2�yt�}�?&��d�{*��{�nn�f�/l�+�(R���RM���}���.���Y���z�\T�xfId%�6�-;�M��S������I�&�R۝�BY�u��)��r6n�Y���ɐ�!l3�b,�c�F7
�g���0*�g|@W~�!���|�G#��}I��{�Ã��C�t�6	������;|�s�N�|� ��<� ��T����q��{�M
�]N&<j2���?u�`H���y�}Ӌ�l�w|�����v���ߚ��46�:rTi��\Ҟ&�X��Z�gټB^4��R��Cy��k|��W��ΩA�d�A}3,���o��	&����,g�Ӓ�[�fm�>4�b�vi�%Y�0�p�!�� zj�>/��-�`��n����n��%�X��Z����Fb~Ӳ+����~H"lDSp��f��XS��������A��ll�I�iq��@!��qt[����(S&���8�6����l�������a6;A��Oc���f̮�j��;i�����2���/$����8�o�~��a��nʸ �O��� MfP%�L�4���{\W� rG6h�)�!&p������K��~LO
�
1���[�~�l����'����V!S��&DrN#�)mU��9�t��6�bE����iZ�����}�@x<} ٳe�h�ݰ�5�b�<����rDX7}�:eWJ����יo��2,������ ��� �Ѝp'g�?G\a�q�uj �N�����ic�3�����.�Vj
�"�� �w7cn�`>�����#�k]�p1�~a���l>���9�x��\�(�T��Q��(�Ĩ��n,ka���L�590�	���WXE�{�l\{z���4��ii�i�����Ԉ��hPd���,����9h�]��-|���z��8�����	�J|�� FiY��v��~�q�� \�-�)����X��x~b9�/�I)�3�}��F���t�ePQiD��LU�BD(\���V�RIje��j̰I>�)�A7|��.��,�/~�\0}1�m�D��>�ӝ�`]�ऌk&�TJz�B}4��JR�2�a���Y��2����0����������d�~`�2׎��^�N��K�����rH�L":�
7��'�����J�	D��*m{�oA������	���x�bS��c�D����T�&.	]s�8ρ$�ľ?�BL��ɳ%��|�@��mJ��; m:�+��)
�?n|���C��-�O֡���KQ������<wO}��䘇ո��1����n'�:��-��N����5.f�y�
�J�}��x�,��,�o����~�y�ae!��u�Tpm1��Z*����j�v�������o���H��N���G��숉���/���mW\�ɚ�a���q0�X�+Rʡ�D��l�;��g�:��5���eG�"|_S��na��*7�E��:�Hwa-��S=N�FF�������W�5Z�D��w��ZG,ך��L)o٪��W���~�ꨌ:	�H����w�M�E�q�dW�Q�2�X�������#Su�̅��@F�-���M��ɨ*������jJ̞�`�6紭� ��sޟ.~��d��0��/�)�	2����Ήٸ�G<С���lw�]�6���U���S͜�G�'���c��+xV�}D�($�mX(k�~��]A�����rK�H�����G��ꎎ�	�J�L@���fBB��A���� �����W�Qe�:�}5(���퍪����?�[������ʀR�aI���w��5Y�8͵�B���>D�10d��-�ݸ/�xA�q_���n�Ȱ���D7��W�Zî�y�#�]Bp�t���� ��{TVgt��u��dZ�D��0�qG�	��]����wυ���Yc=�W.̂���h��NtX����0(�ɪi�Z~OLtn���<FR��P���mv�H�)bZm]���k)�R�
�A�<���'.�����N^��A(�����P֐���v�)~'��>�c��'?SdW�N���r�׶���vp���C9�aJ<�����Ի�a�홗�Ye'g>�^Ԥ�� 'E��6�/� �����f���!>�k.:J8>���m���G=����ʨd�چ���R����mC%OeK*�6`V&n.sѝ��Ay�͵CY�I������P_��
MS�5	LQ��˟�z:ٺs'k+�+1q�l�P��KPj�������_�� 8�^˗��r)�e� h�Ue4�{�]AK3؃� S��~wW����t̘�YA"V`^��'��t��@�MJ.�".@���"8^���~#�6�_`���sk��D@[�Y��������t����\�g�U�Y�l7Fښˑ�ɨ�U�/�?n��"�Z6�+4 9!�|!x����w��~�csc�#f�D������xck�I��x�.8;�3�2���jA�c#�B��+"���ޖ�Z�L��:`�<Ү&��[�2����b<�T1�V��QS'�kMǍ6�_�Ub��oOK���?�����V�;��R�a�-�y�1�~�)�$�F5~3�ĭ�qqF
�\疧|ѐlO�o��@��U����X��Q���D8��(�M�P>1/H�^d�w&^�W��8��U�&�����EC`Xf��\O-��M-�C�ڝ	��ǡM����k;��"���ƻq���c�	��u�$.���9@	qP�(T��[��Y ���
t�|����_�=>.� ^^ҲszY@��xM[}+���>,P<V���v�UU(Wb��z�Iw�6"��X�_�.���G�e��rk]HX|1�����)q�z�O�G���>"&%���
P6���/?�p*ǕS�@�,�=�#�I�8r�5vp9J�L�\����fA��kȞ&=;�`�A����
G5␚Px�#��.^蕶\��bگMƃ7����3����<���a��IPݐWON\�Xp"7#ੲ� �������n+�{&��aR�B]�.��v�5c�#B��d���UiE���e0f�;5��ښ�/7V��dO��eR�_��{�'�����֑��%+��)�'�1�u>G)���4=K�y3Zg��?�a(�Ͻ�D�n�yhY��}$xls�:����~!ұ*�R5��p��g&L�b�e�1^|
'��d���P� ��~I5�Ca@M5�+|Z�P�\���
 �b�6����W$�4�RI�=����2cֈ7�f˱/.c�A�E��c�_b�jq5��;0%q�%�&��Q��|�v�x�Q܃����iPkpC����H�u�\(�����'�A��"��PS��tT.��c�|�E���X(P-;y�on0���P�!OP�*��W?��D�Q��_F�� hm=6�]�Hb�L���`��%�Z%���s)�{J������p�]��=���E )�y�9ǚ5��K�X�d��XH��5Ȃ�]4��%YU���|JYk>�Q�����0RܲT�շ<,�5:��-�9�E^.�S���s�r,�&��v(�_��ն��c�D��a�����
r�q;�Se��&}ۀ4�4+�q���Q��%�����P+a�t�c[����<�з6��Q�מs��|�kY�ç��'���׶��,��Յ�Ƚ!�6�Z`�z��J�����&�%f���Eɮ��P�É�Vhb�T�Px�*ɴ�Y��>�k���= ��?��_���Jǐ�+���CZ�
���ۻ��v��se�"�]�~��c�ԧ�g��W{�y]q�g�����(�k�ol��g��̀}T���(`��5�=N�$��g�����};���Ѝ3_#���/6R��98qw������Sh,�Ԟ�*���
�Tp{K���R�)��%,8d
�px�"q�- �7U���D+[��vF��tN��;Z�*WA�q���'|����j�V_D�;)ӛV�b4��C���5��|x	����R�|/�'�.���N���Er�\���IHi�u�eq�cUD;�5<>���(���zh��O��He=�T����ҵ�7�����b�BϪ��k��� 3��c����xo6���_A����	;�Փ�h�B6��w�*Ha�����P����n7������2y y�Ç���;�n�R]���t�x����;�ǔ��(|�H������[����4c=�3ǥ��f��i��4�h4��*�6Qt�JY�����sw*��~&�ڲD�mn�Ǧu:b�P5D\!/���%����������3��n��w5���j{���j!=Zp:����(LV�
$i)-��}�3kX�Ϥ㩆�8n���4:QG�[���}�H�G��*Xk=���R3��1�
g���Q������䣂QG� ����O��mO��~�v&��Yqzy�B1����i����=�ɑZ�\��b���ӎ���}7A�z'J��"�cw�6�;�-C.��0�Ҽㄭl�'KtXe)�<.Y\_����Q��콏�S�6������0�"nߘr�YHg��R���u*��;���A�o���7;X'��G�R�: ٱ�j	�>iiZ'}��D�� ��<�id���Q�]z��D�� e���bCs#������%�|\B`@���Tq�����5��L�D�BR��ö�.�^s���jk�P�^����t�ϔ�|YS��]��S�|��ڞ��*'6���9x�Vͷb8؂�b�P���f��~3��h���M
q`�YW44�,Cq$´Q�h�B�yY^!{���^�2����J�Ss�ڹ0��ɁE��+Ijl��+����}|�d�C��v�����~��M7.2��������n�6 eu}��|g$���{���@��o�Bmq�l}�m� r8��:�W������^��2�(l����R��:V��J�G+aU&����<�]Y��3���FbdLwT{�"Z�[ ��sV��B��G-���;P�./�%�����@���)�[�+R��(|����3ذ�ISa���E��.�c��F�v���vw�\�f=���-��~b��#Y��ے�.����W�����i$�}���KЈ/M)I��Mֱ7�<�	<�A��}��3_Τ�^t�</k�]r#iKs�Τ+��9ٮ@��>�vg���l`k\c�D���ˍ�?�z/�Ax[����I��j/�R���
9Xl��� ��]�g̕�@���Tv�p�۔HU��R��uJ�U�����i�D�3�!���KS$ؕ~E)?l	׽�?�Q@�YY~�=���6Т�;ق��FdA�y���H.��4��w��W�7�s�'�Дw�}��؆��+7�q��h�^���+Ȯ<�|�����ۭ��{~V���5n��	�Ly��Y��]e�_&�X��S-k�\�U������~�5Ӗ�	���k.6x��Ư"��r���O|_���V
�j26'�!ZGo!BOr�3e�!��U{kc��@��V��!Kk���]'/R1S���B��z��2����5k��v�$c��(�!��VM��*���hU����v��t��uY%p�w}�7��>{+�T�GD�_9Y���9��֐d)qG{�]�}�-0�RActi�Q�5�� #�,?F��HO���6�me���Olξ�fcZ:�k�Ku+8��5EG8L?�������'�:n�Y5ص��K�!��
%�*M��_��N(��*��ǐx��M�~QڕO$�P�dfVmb;.kX�Ig^���3���MTiώY�=�%a���r�kO�K퇊m�]
<w ?Kv~4�rAen�c+��h<�rL�ߙ8��x���Ò�GQl�nop��>Z/��K�qM��W��n��2O.:9t�.Z�
6���2k�c9u������ެ0I&kߑ貮]t���v�vg���H9�����Jz�!u�|<iyzN��C���*�����"�K�����v�,�Y�\;'�?�R�����{k,���B¼�b�ҙ��v�مm�|I�l�|���5)�l��P���*�M��]�%�&�O��yͤ:hJ��ٝ�71QEG=q��E�n~�z����dc��嵺�{�G�n���rg��@p�2F��@�^ٚ�XlSRe�ǨW��@�OA�9ם������B����}8�q+�> ,a�gi�������m�e�1Un�K�3~��:Z`!u��koP�(L�J�y��s�bNN��l�P�\`#�ڱ��	���&���	�?�d8��:d��}v�?��y!t�`�[�����-#Gje�5��P0�7�._���r�����_J�{�(n�l��ڝ�*#��H\�9k�_�Y��j���|��
����*�Jgd���CB;�G�A���A��
}R��ƾg*�d�دG���oQ�)g6�4�n�b��۠��<��_��(���"���i�%��V4x�5܊�&�'x�]'×C;\\��r�S+8c��O�}��� ����Ma�����.�ɩ:�XW9!7i ����/0d=ʔ�I�f��X�Xۇ���Nǫx]�6	��\��x�D]�aE޹_�W�TWX�6�f�C/ͰL�J@'���=r�����s�}q�5��6�d�۾���T�[���vS>~ck��G�8�����x85}�<*���Q�k[� �OI�Р���N���-�[
���@�,N/@GAO !��S��C���*�L���{W��,� �I�e/w�%b�k�S�9_"��6�����������4K��Zw �w�����%A���m��#��T~�Z0^�"��J<�H �� ~bg}�ӯ_�����3K��2�/b6���d)&��J�(/�}�'�����:�dN�\�W�̘�ѯAnH�r]i
��r��K��ٝj�	���2q��]]����bR�z�ޗ�C n�����:�Q��.�Yh����`^��v
��Jf�\ř��G���3S!�G��j��_v��ُ_�%�'�V i�;HR����Ł�J7����.,{F
�T�$P�. w�2[�KE:\�a�^Ld�D?Y@@pz.;��sYt)z����@��R�ʽrI!Y	`�G[;|sX�yUS���N)UJ�r�dZ�NGCA�d�u��!S~�7.~��i�<�ᅙf�����<��ׯ���T�d��bT�{M�6�(~��W��W����g/3�fA���;�y_p��U�7F2���b�:�J�����:P�}1�Wʤd����Xi'%i"�OW���oi�d~�aO`��~�<b?0ʄ�\��a<{L}�_zgR�ډpl����*HX*��������fDMz:��d���ԋZ+wƾW ��V��bc�嬕h6��&�U/�0�_����6��M�H�\��%�[�F�j��*9Xa�xU�Ҩru�fM���@X0a93^*Z$�!	P�7x ����8�F�5:0G�wъ�������_�|���I�ˬ�v�}xP� |8A��k(�,���*��t�U@��WH��ʯ��2@V��,��g�d���VR�t��_��3��ǻ$�TɎ�� �rٿ����,�����)#�"� L�j�������+/�]9�L�9�V��MyOΕ�\���I[���*�Ӡ�C˅uHt#�T�H�C�e&����:�}��v��i�CES9�-��0��R���T���Qi�*� 2�\��'����([O�y����6s� �v��e�@"c4�.-ĳ璽kt���S428\Y��]:�c�yl�X�'�X��2�Z=~�G�[��T?N�5���)6�ٝ���P��P�|t��k�-^�� �&����RO� �h�1��%���MY 31�gs��W������Cy�p��]��m0�I��sK���j[�I���fП �'5��i��X��� -]!d}OS�M����E TV��$��(��d��ѐ����~�ȏJ�LҜ]�F�8�ï^�(,����`�<tc���'oTw|R5n���ӛ_3D-�+�ɥ����Ɠ�>ֵi8���T^]�����G�';���!�#X!�3I�wW6�8Ȳ�w���ن)]��a�ڰ��דHph�nD�P�� �6��e�V��G-Du��^����@�B��%3ȠX�	���2 ��s�]_��:ru7�3��;[�`\F�.D&���Ўݕ�qyH����l�%]��@�'��I�����Y����#_�AX!��G rz��ᷗ���8c�!ln}`5\�vS���>G�~�z�U7nD����u���0�o�X2���m����:�X�y����=���mЂHT����@��.�[�����s�K"`��$քp�ڥ��J�3��ݎ�45�4(|�2?z C3r�z��>��Z�QŬ��(�l���4l���۱�}+P	p� �G�zѨ�*����l%�ʳ�r����{���w����z�}�>/-�[����)sJ�vbvΈ����D��Au����eN��GO�������c��}�a���]�Ie���u{��?0-�dx �fj���g�����k�P7|���Q��}#]���4����-u�c�:������us�����T����l�:-�^���3u=+ѤI%�?Q��C�6z����rK/A2N�lBnA-1�Τ֐�H��Ż��>��y�"���%|̈H 㨡��V!�[�� 
?x:��&6;W��Ia{�68SR��&!1�~�4�?����S�{�n�>�+�&7��L�Zqb�^\&�n�=)�ZN�{���EL�0=�.�����p7}��*�&V�`�L�ׂ_��wiS�s���z�Gt |r�(;���G�������G�b�7s���_q�	�|a:��v�e˦��tĉ82�JW�ٺ�;�U�0ɴ�]e4h����b�+�pGI�#j{3�6��o��z��m���h~Fg�5�IJ��	͘bv|�x`Q!�:��d�D���+��R���O�MDK�=���e^��]����%�m�?�w���?M�Ў���		?�j�x�|�jV΅d�x���X�ߚAD��wHЅ�u���'�
y��,���O�T3��2�~��;���ŸQn�e;���f@�lw|�gDM�a���c�VCш$��s@��S������������'��Vq���ޝ�Zfw���;в��\�>�ކ�7����L5�vm�����a��LH	�6�Q�DL�e�jW��8�))����ϗ�sU�w�;�F�?sJ�C=SB����	/��[���|�XQm K�9
�C �ؚfřNv��ćaB�f�Q ��:HEJ�hb�����E.�s^�iX&&������@�i�*�[�R2$�0��dt����^��YZ��>|������a�h��1z�� �f"�U�"���mB�ͣ0L~x���ùb��5{n["�Z��Ǝ�"8�Fؑ{,�C'����$�;ncL��Y�U����j!Փ�J����l���]C��ͬb���G�& ��e���<\��j|
�I���6:|J��r\�T�y�=�g��3d��b�5!�z;V��yo��̜�;�-��w�k���
�� z��UÂ�<w2r&��K���R�#4��*Aj`'������,�׌�o��A	$�`H�M!	�\Z��Eëj~~�#��^��bP2���k9�>Xy#A�ց|��YA�� i+w���#�-��`���ڹ�fv��v�U��y�����T3�(�#_f�=]?���m�a�Ĕ0�0[2�̆G�Tf�)�i�!�Le��5�w?M;.���pdh�N�K&��"�C��	�����W�+��_wR�L"f��}�W7�2���p�⏑�,����P��p����fe�j6r��x.�6�w�ݖ�L���G�tjn��_\������=�hd�ͳo7�5A�}�� ����»͸h
gI����|N��p���c���h<��@�l���`9�����Ts��� 4�������)��h�D�l0#h(�-4�Ӭۿ�ţ����)?+6��,�n`�&��9O���~�nX֞�G�*���ψ'�4p��0�4�H�!iT����iI��o�?�	'��ރ�(Z�EE��m�����k,
�?t�SG��kC\A7=����J�ܴ�R��S�9��ǹ<�.�?2����Ν�a�'Q�>�S�����N��fl-~A��)�a�rh��D)�w�Ԓ�pU�̟рs�N�|���uw�üP��,4'Ra��E�֥�w3�B�W�y��O���\YY ْ��&��p�?����k�0w0�g5yf�t��2wU�Λc��7>�/t��>o��C���c]R���H���1[mW�]Um+h�!O+��[i�(�6�8��b ^2��0�S���=i�O�u=�4ZƠQ~���c!��p�� �*��{&��#�~�t�^�LC0{.0R��m����������5̛t�g-���ÆVl��u�B�B|,����HckNh��D�9T	 2]�)aQ�N��p�^94�v�Q{�ɽ�^Wv;���c4�=�*B19�Y��-r@�T��[���r�h�:����K�uR@�Q.n�S�+9  ��*��� ��,6��yۜ'����Oy��F[���H75nRd����ȇ�,�
���c���ηuY��H�E�%[&�JTPHn���S��M�u��ه���Ż�<���F4̧-=�:{]��>�J�.BÞ�|ceCU"E�f�η3;�1t��Fd)h��ltn�	�&�(#�Dv@���G�� ދ=2�ST��I�7P$R{��U�.��E�uB�{���7����ݩUf��3}�� ��[��bu�V"��7Oа�)n�e1��
Y�?��i�
;E��@�PE�5��XcX<XNjhU�iJ~�����W6K�>�	`��t��q�bݫX��q�Y�
]͛38^��-k/
q�k�����l)s�i|�w+���'���_e�&���1�_���yF&f�wD߿���5�i�(p�E�O����FFܣ�G%w�S2d%3���B�ƒxdo�Z
�*���hʧ�gV��烷-4)���L~�����]�`�&�����h76tKa��Z$W�O��{��])�?X��g~�р�7;#�N�'��6<vw�I�R��FɅ#�����y
��^P�\m<H�c�>m�p��������Vc���Nb4:�f��J��˯Z���χX���|�{m�����xغ�N���̹R��&����_��1��.@�M�i�	$���P�4F[.��Q$յJ�o	#��mN�XB� I�i��<B^T7̑��6�5"�h��p�6�̮H��48FLЍP�&�M�3s	�?�x��m���ȣrC7��
���6!�?����r��Q_(���K�l��<�Z����r��5X.&����F(�s�O���kL��.����K����u�dR�]�4Z|+YlN��P2~�&��xw�/�w�<*��o�cm��X9C?�l��x�1����'c�) \+���RԮe�U��om��:���~��C���ϊV��/P8(zDG�N�KT�=W��k�%eڕ�M_!��t�ū�IE_>���2�;w*O
l��E���W��f���;��'ay']Ŭ�k)d2���KH���Pj[Y�"'w΄&2�X�<Z�	:���+ޒM0� �M����*��1��E�^x����![�k��k*�2k���v�h5UΙ�F�G���)�iF���$z =;<�H��nn���b<��\hD�)@0�{�Z�0y�jD�Y�w��q���4����
F�7�l��S]�GY�?�"��x�k$�>wS��q�}����ݪ�%��Ў��S@5�8f-]=��
�aAC�ν.�2f�D�eS��me~ώ��D|͎8��r�ʻoc�<�"��N�@�rU�g蔌����^~�Lh��Y�ܓ���XȥoCh�֙�f��Qc��&�`��$-'p���{x&`kkG�1�x�v J�>�R@	w�e��Ykb�ïx�q4)Ob0Q�y@D�twf���Ƅ� ��i|Fv����u(K��Ll3��NM�FA�� S�c�1��v���_�9� Cì���_5L"e�?�x��KJ�A@�������lʖ
��6�,�<�w�z||g�on����@�Q��^9e8δ�1k�w���c�}�V^��I#���摽T;�v3CA �A���(�q�Qh`7}�5��"���
�ˋ�B��Ly���k,Y�*>h~p���V�sE4�%A�Bh�u5�"��4��yRe�a0;�oBR��?~��m����ԛJ����k*g�4�e�z��L6RaOS���oX@�B��[D Cڌw��x1�L#P��qeke���G8l��U�pD�g�]��A"��_��H���A8^�����Ls����G�F+9�=R0+���v���t��L�5���ioB�Oe���HO����΍�Р`�gl�wIgo��^4\�RzWw��hr��{��� ,U5>_ԭ��C�k3��h�� �+�*]z�P�s�yDy�=_5���Q�ˣ?7�M�`a3^&c��]M���qX�&�b�{�RՄ(y����B�&o�}���xR�	�g��2�RQ;牯T���0��\ļ粇��Wl������{>0����	|O��W�']N+

�D���w�����|�$��
����ǀ)d��!�7J
�Ρ��H'�Q����+���Z�o~u�1���H�!פ�Td;JK�B*�Pe]8Z��V(�ǿsZc��A���G&C���8�B=��x�C���B���j_c��֙\�7@��ki��ʷ�2nz�F�R���5�_���%�w��Er[��/� ��aP���0��ׄ��d����ט!��p���Θ�W��}QCկV�]W�e��U��\��X!�A�\�%<�UGCI}���r&*����faq�ud�|ѐ߼��)1�<Oy��q��@�3T����Gw�p�/4d�xuҫ��G�	��V�;���&�o��m��M�������+A��aڱ�)r���d�ዉ����;Qǖ��^{2��c�dZ�+��dk�#m�%�֐��{#׈��Hc�T=��L�=�Q�;�" s����<lD?ƃbx3Զ7���+��s.b�ڃ�oh~u�k)M^W�Yw������u�K&�n�ݣ�&ڬ������mW���d)O�F�����������V<��W�{��8���E�Ve�N�]��i�[��S+�W�u�����Z�hh�LP ����d����Sx�9���'����(}��q,�����R�@���P{�ʞEJ`$��������m�0����Ҹ
=Y��pZ8�*Ц�Z��/�,l-�*Il��#�|HJ]}z��;o���G�5l�bxǍΊZ�Šc��AN�}�C��������S�9��9Q��&iT�~O�ۑn�VZ�Y�Y�Qb;�Vp��췼L_�Ir���GC=�����!��U�+y�KD��:m"����D`+�?bo�;��:����fdTj��mr����P{�HY�|�"��ɩ�P��/B���u�p�=��:�����?:�R6��P4_&��n��X��oɯ[9b�}���1�e�aA9��V/uY@����yNId�%���w�*�
�z�P�#1�V��9�8��+$�__��a�0g�U�>��� 	���4~\���O[Q_��z� �$��r@�5��i���M��+i���z?AAπ�!�~��n��V��Ӻg �^���ׄ&^�j�F%/��g�g�ڷ���`\�EA��N�l	����'7�N��%�L���L�z��4*ύn�{ޑ�cQ��9����F�[H�Vԗ ��A�&��l��r��>9j�%�4[���ޔ�s��mv����i��4�cK�$�?b�K�(6h��1�!��F�.g�B²�N�7�ُ��������Zj�"�W{b>/p��T/a�,���O��]eě��`�N7g�BS�����ֲ�|غK�l�O��}pȎ���q�w|���g"���~H����)�``�d��~2, �h<��f��;\#��f��}��i??b9�7�\��o�w��y�X��_�%����ZY��X��������-Ť���M�l��F���*����J悅6�7�S#�{��%״o2�ML"xF�+���F�p,7�At�^#yie����a�CL@Z��H��?;����R��\�ۻ�p�BC~>�A������~�m�_�C�1�9����3�³����f������� �{�X�� ��{�K`d��C@��2fm���O��΀����v�4�.w
�bbut�tdz�W�i��ЌF8ݣ3d>���4�(��)w)���'�RFb�me�ړ���p��4�������z�����k����7�p���g���&�_S�����s�
�8��O2�0�t�Wj*H��r�xƬ�Nn�Z��ONS�}�34��n�C�CM�S\�S��P�}�R�|����S�D�F޶�z�'�.��t�ɂ�}�Bמ1?`��+E�{��`���T���t�!��j�0�]�_P���]���DE So���c�
�7+�����]H�E�vR���`(��Ϟ}���^�C���ޗ�bo�H=Z�PA�Euđ����!��px��J�(������Oе������z@��U���(�A��W�KLv��0�vҦ����h��j��0O���G�c��e�-H��J�q�����RJ�t-r�a|�^��.Ǭ}�sD[�k�^x.R�
��/�!���ann@�῭ٺ�h	}��j��JF)-ʲ�:��j2��
R����3=:ޟ0�M�[kH�-D���W^���c��c�8:&j��L�b`lڤ����Cɭr���S4�k�� �~��������uvy���-t��u���Xh�ݯ��H� �ۍ���<�j��HQ��;��"�'�-3�82��B͝�f[:�-D������b)"W ��0�jZiZ'i�gcO }/����z�U;���Z<� �ڒ:���������mt"������BD۫��%�1��#E�<!���Q�\�$=�Z( O���K�	���aW�s,�(x2Ƿj��Kk6�����rk�����G�1��vC4T<+�RxO�ބUm�!�S�Lv����l׽s�����w��р��fӃK��i9��΀&��"gZ�I���'O�|���!i��F���|��Oq�$�)�m��F�i�hnVYF6d��^�����]�״$����ؘ~�e�A����F4@"�,���
�Wu�  t��^��8�*�G�Y9v�'1�,N�2���QK�xB
��4͗�;j��R�]�!+��G��#��Mme����e"��I&�Z����Ѐ�BA��R��g�ҬT�kB�w��U73ｮ���X�㵶ld&��ñ� [RX7f���	�?2��8J��p曐�=�q�Ө����½dX��ni#p<=�J����R�(H3GG��]����6>w�zQ��JXO���soƫt�M�SXCh2��?W
M�WV����z�F
c���1�+�:��j[�MCkd7�;Q-x�J�'
�Un��b�H��@N؇���46|D�X�}��MMAĒq�uɮ̱P�J^̚gR!��]!^X;�L��K���~�������$�;�+.C���2��f'D&F��+�c����e�f�K�BP׮W�ߨ9=�m�/�m!�������zZ7Vޯ����_cy0:�P/5ۑ�5t0񝝱*�\��.��
w�@��Fy������b�%-��Bѡ�/�D�$��04�Tִ�֫v�uo�c��R��]�=�v���7�a'g{P�.�������Ԅ�R	mE��Gfwqġ=��.
��P�m�2�C�����¸s�1�TZ�U�����w���K��+|Tه�H�)8�	3? ZG����%��6_��ns��%��~�6�#���鷳H�B��a��E;{ѡ����'N��ݯҎC��Y�4('t4NB�B�2J����N�TQ����DDT^��7����X68wj9�e�C#hQ�<!!sC�%�G��T����/�`����@PV0�������lB!��~�p	CΥ2 32�RK�#½�|nUI�zU7���d�i�N��;�E�NPB�H�;}�P���+�>j�=��+,"�3sO��J�����S��2�q�[D���*[���-O�p���Հ���ͨ��N��G��8s��#�G���2�naB�;����&ig���&"O��L�&�"dvs��CG�O�l��� �;�w^ �Ů(���@9� �)�loǰM&�ɛ���}wE��؝o�RތFd�5t�p���n�_��y���ñ!�`N��Â,v��.Eϩ� �l��:�g�j��mH�3�w�c��N>��5۫)��w�m�B
\g�lힺ�$��q�jo*08��}k��]� $W8h�ٮ(��V������Ĩ�G�+�y-(]����*���6���r�Ac%IU���;p�;�\q��RS�D�������%z_���"�>�/�.8��_�o!����@h����b�GDI�QJ0)��G3�>�Lm�|�
�썤�Ӂ���lxF����I4��@��rk!�/D�}�|�hF�����q���o�,ѻ��+�E�~���,�7�=2Y�������aܺW;ĖLd�?Ҧ�g1�8��EeԘU��J�6��rl˦��5�gJI �r�?>��j]�p@
%��\,��4�� �$�������S��Z��.�~
�yl:��4�y��I臈��C0�:g(�_�b GXHZ���(�bh���#��Ur�⩣\B�/�Me��$8�}�&�A �g���W������X��v�������U+"Nݬ3�_y^��kր����d��y�4O8L���5�Us�J���D������-�~���吣�$�KN��#��x�+�ZT���)�7L�QzjC�D�16�����ͧ�W
8��hi�!Z�Ge�㜊��o?���ƮDR��P�(N"e���88A��j�"���~���F�.fo;� Ҩ��v>e�(��ѵ������.�x��e:�5��U*�I!2nDdwO�P��������&���3�3�"�,�;d2}���y�ߵ<�r��M�Tm�"w�����"=�לn�>��
6s���퀖OA;����y�T�G���f��uL�k?m��[E3cTD�Z�?Ȉ2��������*R&�&�{���_8km1i���N+q%N�+OP�[�^�!�.2��Ǒ�&a����6z�5�g��!��e�)�sW�����N��j���aY�d���#���7������b�w0̏��ڵjp��඲eV9�8�C'W�i�R?��r�ot��_��u�ܻF-���ͶEt_�X(B��T��<f0�@�p��ZP���A��Η1f���G�5�锝��LVΒ�D�Mb��tNb���I��<;�B�-�G�I��){l@@MB��	A1�N ����-�Y~6����7�Mp�&������}��my��x���#���q����zz('V�LQY���Q��B|��ۏ���^�Tv�v�L�b6]n�+H��3���A��[O��C���̭m�����u�%'��:�/�3~S��z%F�C-�T�ʇ"��el[�&�f�J�̢�59��$*��O��gxhE�T��u��n��I�W��;Q���YT�N�������)A����盏�$�^�8�fnz�^px��㓰� �j�1	dB��'�@���jO�{F�	�.��2@q���\Qm�*0�v:u����*O.9H��e���|ix�L��O�ƺ�R����[��H%���6�p�Qmí�(hՌ{�BF��Rx�1o�!{�ӝ���G���B�˗)� HҐ��̅2��F��/��({�fkځޑ ���G�����kl9Aj�,,���n���TJ���I%�I��;�l��H�OЭ���=�k|��a8H���2��+��1��-I�p�[ǋsCSy�0`���'	�=�
�L��G�cr�����՚�h��X�KT�r���x[B$�D�����ј.M̽0��u>�,"w�U@@�J�0P烧�v�Bw��I���b$ϩ)4��ԧ��G�󇁣�lg��#)F�^������]}��C���<!�/҉8k9M�VY!�����:��z�P�}A7ɺ<�ʙ��1��ζIK���SK�}� 1ܡL��d�a�Wu�X�"Ka������k2s�`��&�#71Q�봴�����x:�$퓋�C��Q�\OK��Uz{:$�@�)�5�▬���� ��T�
P�d��@s�9~bo&:hR�%Z��6��2<aT������isw6Mt~��֬+!�u/��^�yR�'~e4�v���Pڷxz�� km�/��ͪ��Zv����:��Չ<d�:�g�j��x�sQ}�������qk��N�
�
T���@�A��4k�,�azf�.��T�oH��n��i����c�pN'hF���q���2E@"�}B����s��V�H��qvQa�$��t��8������ֶ�	y�烎�@���3鷁[���IKiП�����T�ۂ�ܡ�߽����J?�4;��JF]�/@*�I����α&����Jm����i���sI�G����@ް�Iܯ:~=x�55L�_��L`^bw{���l���o�&�}KO4�U��Pj����m���4g~�V)�:�0s���a� 1�<g������]�Jn,��ugI�$�F6EM�K�o_a������_L	�����.�{=�"[��ˬR*5�T@Č��{����G�gA�"�R�r���'�X��g~��z�]U@���f�j��L�у3Wl���U��k<�a�@�� c4:�C��4���t�s�a�����?�d���g@.��"�
���I����h����U��rt=L��z0ϻ�S���#~n�؀`�sq7k!�,�u(�a�7��=�-o���7�{~c9���J�c�.+�D����D��V�}�aj�6��d=y�&-�wc�߄Z�E5��pic��.�^.���[�4�w����;Z��zQ�J���3:��zt��A�~��t���ac9��@����#M��j��w!�줯�d%!��1�<+� �~<)��I�yR���=���~�bs@��g�`[�6,���"��YG�K�-�ԯ���Q�l)C�R���2�~Ū-�{䂎��(ʉ�s_cˤ��?b�QO�a��,�86/3�.�د ��-(�a����ٱ��2U�\n����g!|��2�����c���y>]�1���Ő�\�*B�,�8�w6Ww�nn��1���1���ܨN+⸹����	�웩����gU|�u��Z�1Q�E�¯�ݧ~#ma��X��v8�C\EϏ�B�%�
�xGp��	�%���sZ�L;C+Xⶦ�;���*�Pz���� �w}}������|�C��r��K?g􅄬Bn�z��
:�v���N �����ӵV�Y��ڦG��2.�O�l�-3�m.su]�l����推)�"&��龚�����h�T�gb6O���t`��#1�����6����S4>��8�k�d��|6�G�&�/Tb�jS,~	�]����rE���M���I)4�%G1*�:�����3��,I�6����9Bs����>�%��Q��9T_f�⨅*�UX2��R��ʓs�TDC6����X���^���� |�*����`���hC:$�в��ӂ�{NٺKkyR������zi?�����؜��7qr������.�"��5CL\�K_w�t�}���i��y���������$B�oڣ,��E��L{%;��l%��Qg��R�.~��_�qM�~���Y8{�+��q"K�u)�DBpmY��D.#xƼ��o�����p��.�i�i?h��Nk�.J�mZ��!}��Z��s��,>�GK5�1M�H~._��@#s����B��e7^�[I9f�3ެ&�H��U;K�a�S|MZ�ɓz!Ǥ�P���%Z=1��&� ��"��+��@+J�d_g�8(K�D�)�O�����5� �Iu��'�|H�+��
>��l^
4��Kՙ�f^4˘�h8g-yn�"�z���[�~'������;D۝dj4�ڼɁŪ��j�  �c�N�{��� z p������ںIho��]#gh�
���2Z^�:��B�bms�r�|�n�T�5)YN��B�5[�ZJˎN��������>����bUvRF\���u�:T���ů��X�K2��ĩ�&��-�R�-�r�[ei+uݺy�- �177ʩq�l����yh<,��[�B���9��GHx��-�(�4�7�u���!�YΣ'u��:_ڦs�Z��й�~�@���RҞc�Ϭь�Wp�
�%W���1<�!Bj�il���z�=����N��фs���m,����K�c�@���Y���r,~��:�w ���^��~��"�
��ߧ7��dӶC�L�|���atL ��p�7Lf�������	��D�~k�a������y���s�
�����Һ�BT$���?B����SC��c�_��*�T���HT��������Wfs:�	����KUes���(�t�.��*�XARI�p&qŕ��ٽ��1�(��>��T�S�X[g�Yә"�o��rF}��~�>J���L�ɁG_3ʌ��L�����������m�R��Q��J
���AI)U.,� ֒�3H�73��tomx7x�'4 ��k �1�k��8����7A�J�6 f�����=}�eTn�Ay���S�X]K�69`��7�52����N���_*�w8hW�
� zs*�RT?O1��
m����I]������կ�j6��8����5h6O p(��O����<��m�Lxs�CϠ�%�p��V�_���U�f@������5ከ�6~��'��p���k�|_vڞ�`�b���T-U��YJ�e��4p��� ���-	�6�O�A�˄-|�*$C�d$:�o��y�LMDyHXo�\^�Nu���g}�gP�Lx�JHF'������D~�WF�1��4�4%;� l�K�LE<?�ucx�6P�>]�V��>����]��ʩ�?{3�y���	:��ޣ\�ʟ�ț}tf����pO���@W�a���	$-⠀&�-\�n��40����Li�����Yb4�ɽ��)�N~��.�"R��i�=}󏨙��Y?�9��K��`�x�K\�9���77�D���ʎ4D�/�JGY�u����ш-8��,ߴ*��sK��Ee[�=�i\�ic���U�t���!kb3��)Lף>�H�(�n�m��=���2C$&tB�2��y�O��z�k沮��Ƹ(Ƨ��N�Q-0-3��M�?���t�I�]�M�2g1�pV��IT݁��Q��8��u��ܕŽ)Ҍ _Ǚ��1f���w�5m��#� �zx4��AL������$[0�=�$���osD(C�&@YJ^Īk&H��������0�K��zv�_��X(��^�\k>��/�q�c"����#�
O]� ^q ��rl����M��B�Cﺜ�,�������yvJ�#;8������G5��V� ��s�_��`M��Ś���+�D��>�S��ϗ�@��⤂��}X)�+ �Ȍ3��c�a�
\�n�7���Y�8x�n(�p���J�L2�{�¡��`��㶵��B^"����[2���9��F�Wsy�u��w���W��y̾Nl�^sO��I=|���������O�Ký_.�!���@Ͻ۷{�������]�^�a��ԑ��р��l��MŮ��0��)i�7)���ZW��)5��Iӗ���ٓ-�����\�f��s=
��d���@��/�ɛ惲�Ԍ-�� F�����۠ ���9���M�N�ot�l�!�B���g�����|_%�mȝE��� z }'��.�l��s㯣��O�`Vta�����S~���5^:CSbL惫o�/7W�N�#��֔�\�Ϗ'�� KP9��Yjd�m㑯4]���
��	����Ў�����BÄ�����g�/;^�ucT����,�ɝ�/���ƭ}�oy��6������wE~7a�-lW! ��Hʔ���Ӱ���?JM�3l �
�"��(��J�l�-f�h�����9'۾���	M,0�)����Ռt9Ӟ"7��K(�YUܜ(
coV�F[����1h�2H��}�[���JC ��d�щ���q�[�g������EH���B�J`��m��,��7��w�>o7���M9#N��<����Q  c���`*�;�� �x��]�/؆`i�!a�!3���❋�������SݝX6f9�|_5N�#{�c�?�א��	6�>G&��(Wb��i|=Ⅴ�ҟ �0S$}�V@b��o5<��{H#l�dbu�z !(����-Q��q�(������8�d�"Ja��Br�6Y���)��X�w`�Y��'�#�u6hP�k%w%Y�X��V�(7-&H&an~�EI��)����~v�HZ|����"�������p�G����6V��n�s�C<H~�1�����?��<͘!x ��`���oyj��T`���(�����uM `��	u3H5�~,�	�gO�!<:Ӌ)�0�+�p[h��+n۞��S~y�1�w�A�j�1����c"��0�b�$���o,���J���8�+(ȥ��E�}��3���ڻg�A�榚ʫO`�ܕ[׮����1�?j�+Ԯ�5�|A�
L���l�j$;m��rd���/�	}=�J���[����:*z�)T��K`kx��s��СPx�_�6�����B�dXCΐ��D0!�o�O+��Aܹ��R[��^�JA�9��� d�s��SOI��!4��4ǵ��R U:� ��ΜU[u$���4#�1m8����h�)=ަ"x�_x�l��Ǒ�m�(�o�n�ǉ��1�Т���7<
���N�� 81&l�1���즍�l$QX�*0�k�h~�8R�(�m1��V3���%��TC��o�!�h:����kP�H�js�xxO�<\���/$�4̏f>��ru7S�L��g����-�3V���[���Q꼽��xAUz���i�̧�i]եQ���<XDى�IY^�6�e$j�^�3E<�1y=���n��.�#��X��ږ�}/�%����܀�¶íZ��u��5+�=F�-w���)���{��v>�t������+29v�܎��G��)�(jeZ�ǫ����e�>�}j���즮t�!�
*���k0=�	���T?4���=	�i����E0D���P������T��y_Xq�u^1��rZs;��t�7�^�� ��T?o`�����
q�#75��aαNch�,�r�;�.�hB��-H^�W���ZCct�۽�#��	� �f~j{D}��u%��S�y��������� ^!N�6�OS�FX[����VbMvB-��R^�M��Q�AU�2p�^���]��Ń5�4�F��?6o¤��#]w�f���*0>֦�ʞ:J�^�Ӧs�Vً�Kl���0Gj?iz|��F�D�U"r�D�