��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VYs�<b��3H�&�fE	ͥ+u�tZdx��t���4���2�@n_�'�����>�쫺i��X�������E��Ӄ|;X{���?5�dӔF�:���<���&R희�g�kxbV�B}�㏥f��0�ks����c�;��Lr_��#��c_����G����b<Ô1��@,�b	�����d�C�٭MO���|�Rv�
x��C���p.�x�r>2���t�qcL��bR�8���O��A$�79�5��UL��,D�9�N���#Ӌ5�	9�T]�[&�&[�ˬ�I�S����G���]��*f�ő���l>-$OY����� �ԛ�|���%��h�^�곝{���K�m�a��}
K����QS��S��4����"�]�P���Ah���+�׽g�qs��I��M'j���:
��5�=��ū=Y�6�E��QJ���xO�h�<�~��I�-�t����������&��.,A���b%�O��L�AAi
��V���g>oI*��˳>;�c����3'I�#ʱ8�t.�����J����O����9�H*�6!��,����Ņ~q�U�/��Ϫd83��2`
��-eG6$�$F�bU�r^���|�H|G�%���I���?��yg2˾%
K�˅��~e�Eh�I�4��q8�I����z�������𑪟�o���3U�P�X@�G'�7�J��
���l\�aI4�uտ��b�9rm�[�Y��=a.���:��΍����rÁ����S�G���f�!m<��'��2�(=aH�k���qZȅ~��[�x�+H1�\�1D��4փ��g,�xf0殮���������v��{B�X�jl���_S� �n�D��c*�������{��l;�+Ͼ�0��((F���-�V�ȈOx�;~B<)D+z���������82$&�)�$���Nj��HҧzFt�o�ڝN�)c��h��;���5�q�Bh��:��$����U��=:v�y����"s�n��Ə�O�Z�Vk�q����HA�X��f���+���<�0�	��^���x�<u��q90�*�i�5�P|z"��ʓ�.^��^-��n3�n��6�Mss\�v��\r52_�ё&;Ι��0O��cv�r��^�Z]̽G����|7���X�B��=J��rԟ���Hp�w�g
�5	Hs�au��r0Ɖ�
�q��J�|��6�F�sEr��_qh�R���O���Wn/��?r��J�Xy�L�|7"��E�SR0Ӧ�����z�)���U��Kw���p��k�2nujAG�^��<�[�"#�e,O�q1a}��EK��G¢Ķ��to��b�v]�|�� K�����]�����P��rK&�>	�3]�`U��XV3U�G+��<�C�����|��РE���pdm��<�OA��T��Z�fU�T}��Z=���Q�R����}�E%`N��-" �y3��)��^{�uf�����P,�_��>��g�Mk"���O��e���9K����[��7?@�J[�ܯ�g��_#�, �"���V� 2��jd��]d�wn�^�~�-�s�i�1�u1a[���F�·0]����;,',C}:.J�a�	XL�
3�W�o�Ԍ�<�\��<Lg!�X��U�AF�Z��Tr�0��ֻ��I4�{�¼ɼ�PK}��(O�״�����#pC�>�^���jx
�)1���`�'#(�|-�\C�4Vb� ����k�̉��eF�!_�a`���3����_��u�з�B߃�@ ��Cp�u�.�� 7ԩ��k����3i5x�'[�V�iw����
���<e�漇b�<��	b��-G���6m=�q�52���8�����e'�p{�}���y�㣡U����XY�:"�  ��
'��VAd氕JI�����0�#�]T�#��|ǸԊ�]�ǔ�����ɬև������(�xX�Kg�`���:d��g:feދ&���n��0;�dZ}P��R�e�s����[�'Қ$�3�B�a��G��/����Jݔ�-�X�y�|��t��X�#����El�wu�BTLb���|^:S����*������F{Ď�����~�P�~3o�f<��A�����Kf�G�-�<
����@A�����GkN��6º]`�#Z3�����A��\�>z�U�ֱ��a��[�B�8~L�hp��d�svc\�gg0��˭��H���H��զC)AN���o���c�5|�Hg>���'|j��e���p4<6*�������cp_ʖ����$>��*������k~��� ���4��_�.KC+/i�R�?���נ���g.���\LpZk����~B@)�;1̪jXū��bn�WU��:�l����m�3=��W�N6��2
^�a^��		����9K�F$����U�$���3��`����U�8�%�3y��rhL��j3�A�����݆:6]�g�^88N�u��1c5���E✊��CDs�>G
�1s[�E	��ƒL*��pW�[vQܚ=;ޝ�
!,G�\uV�������Gp[���V��T�Z�i�A.��r#��� a*�ҍ�k��IF~�S@%X�����UԳ�c�a[⩉-Ñ��D���-(�TTtz����̳K�ku&���� sbс�]ض(����*��5Hm[��Tg��S���&]:p��n_$�E�fn�cS�g�Z��	�Jk 
B3ek)ҟ3�OlL��}ɩ�_W�/�g5B���k�F��o���%����v],gNx�T0�:,`�lW"�4�x��#�%x�����R)]�Ijf��Jٵ|B�$t�/HSߜo)#�xo��K�)��k_�n�"�����xޅU��;C�ܾ���q$��"7w&
�a�j�_���=��-#��}8��}���ڻ���O�}z�'��]���V�Si����~\�d6� �vS�x{��%�J2Y�$�݃<���@0,>���5O�a����Y}��_��$��b�L8�踇j�HI�t��=��N;��K��]sU�ԍkrk|��"y�S�-�%y\�-86[z����`^�����u��Nѷ3�2ÉQhn+)�ၮ��%��礂'�F�5E���;����Cj9�