��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ��nͳ�R[�ظ�_����Qq���G�]~��\�^�W.Z��ke��X�?�I\�zA@���Y"���a`MBl��$���X���/~%�cg��OU#,��;o�w�F�~�wy�0�Sa��qC�$�_됲��ݗ� ���D��.����v��C��k���<�$J��3��I
����<[�P�}&ʁ_m3�P{�
A���-X'�H4Eml�}-���i���[�f�c�:p�D���� Oދ�o�HN}-��{�/�v��ٺv4~l�N��J�� ���/8rA@��K.z`{��C3��ϋ�����G�4���²g$t\�ޥ(��L�Wv�9��M�=�����w �i����+{dB�TJΆ��g��L��]똫�}�`mi��̸�1�J����WI2ܾj�n������g�0TO����ƒ�`c���������;��Js�'����������n��r�tj�`@RUF�� ���P��^��
H�����_SW�B�4E1bBuH�������mFh��KcR�z	���U����7`��t3)=)�7�!�MMhs���Zr��G��gX�MTlJ"�c6ڏK&�-�n#����-紿Q��c�M�}�F'e�A�\����3����7�ڝ#���>8���,+܂��a�k��Fݑ����]�Bn""����n��r�[kg+�-F��i�5��b}��4�r��*O�^qc:=D4�b��4���U� W��g�>ɺ%��ݨ߻9n��i�M�M�`��
yoi��4YLp|S��t���nbѫ��	�h
V|r_���z��&Z(�J�X$�y�b��@���˂Źj�Ow�8����O�FOޜY�SZ��)
U�д3
��|�Qt�!��VK/����>	�ЀH�<+��Pv���
����:����q�U���\����� �(hK��@'(�Xeaf���2
��c\X�l���	��1h~�hw�s���O<� V�����e۩X�B�����d!��(��u�-��c�n�~B�Er�����N<'�}e�;�&_;pm/z���C~�s��� �S����ȵ���`�!u���yg�-�gC. �>g�'(�t�����5�#Ҋ��GmyS��]_ %mH���H��\��U=�iĆYX3�C?�d�D1�o��v��M4�#mpsF^N�����q�E��4*�=�D��1tu@�=�r�h���=�4�E��q.�c�Le����CzF��J
v6��Hl�m�x	��i�4R�v�KL��Hn���)��mk�EYY0+mn)���%p"��
ۚEc�Q�9檞�L ���,��v�pz�rXڣz&]M���T4���4ˆS^���e�r �ŤD��.�R#-G>JL�44�"�.>6FVc��c�2�p������0���(P�V��o��B��~��q^�g��f�s�M׹���p?	@�Dz��&���H�/:"M�lI4�g�3�9'��	�r��.��t�n�1U����OҦ�}V��h�5N\���']����������H�}�`J��j�C�߇NW��C|�� 
.�� ��s$U�g��KA{����;S-��/�+E�e	'|�<Y`��ȵ��rկ��ا�Ͼ8&����[�Ԟ�e�-$��zeW7��3ҲN���
q+���SV���yл�kk�ו�I�ad�6�IO�-�)!C�6/s�ؘ��P��zA0x�5��W��%�B�}ty��V��ǭ��Hۡ�J��pЈK��{��[㐭o���*�*ٮi�]�GX���ru'����Wlp�UԞ���T�^X�%Y7����|A����_��(��)
^�,��.%���Rz5jUPY���ٰ���f��A���-*ʯ������L]-]�_0�UH�[B�y1m��:+���}V�
c^��4�Cn�r���Y� �S�>H�E�#"���zM�[m��*�L}}�#�7��H�b#jV��pY>Z��`��C����X�Ţ�D�bvG�������vB�Ʃ�߂�D۹�IA��*�dw��u��a5I�^�ÿӸ�I|���<J^N]`�'��g�L����z\���ګ�O\���2�.��̴��Ûb�N����%���U.�yh��,r]��\@o R�Lm��#�bK�QEz`I�R;8��Cs����e%��M�����IA˜qB��}�e���xZ�T#L��C�����[���r�n��Ҡg���r{�Z�˞8b�E�
@�R���S^�:%[lz�"=Ƃ>��!^�0O�W��k�����P��ޢ��:`e��B�[鍷�'qlgE�<�N��E�G����"E;�æm6�e(]�$8��#Q5�a����!�,��BI6�C`����?l6j��1��N!$.>��3+�Q#>���Q�9yG�+$4�PG�S���"�<o���[kds��ό$c��,�F囋#�)������h!��c-\5���Fn�\�@?ÿ�&|\GP.���[`��JeE��(Ά�w!_����-t(�1���ކ�[���Z�;�EUYC�-@Aųס՗_~����)Xs����R���j����J�)?��_����ľ1c�j�f�A��ƿз�՜1�,�A�vY�����$S�&���8��}	y�fm/�'��ZL�UXW]� �N�[J0׾��������=��G��YS��F�u��ʸc'����c��p�Q�r��^'bUr�xԀ3ë4��&�_jQ�(JR2�.һ����qH����$��3��|�y�Ls�S�{���m�RJ�׺��%�zA��x�oi^ۙjA�d��'���Vf�nfB��R�p���"��`}Ç�.P�K�4~*��W��ߥh��/ſK>f�/$�Qd��L��j�K�Ɋ6ޤ�{�Kv�-SC6Q��ZĬ��?��t��"������N1�������s_� ��}9,�����!��ґ��}�	�W�E�Ǽ�@`_n��jky��w�T�y�b$̈$����Ip��k��nd7W�D8�ڗU�P��b����׾"r��U�#�M�jQ)��O܊�Ժ�z_��l�1����}e-���X�6�z��i��U)�ut��v�c��b5\��b�S�%Ї���W/������15���0t�3�2��2q�r��&�s{J�?��������&q���Љ�X:�-��)�I�(����j{�e�w�ɢ��,
(8�ނ�2j2��3aK5�ӢWZ��j�M�'$T_���)G�`�9tS5�htS�4���1�Lav�-*��tO�L�u�R�8�X)�5�?�0}���2�w����U��>k�Yz��Y���`�n<�D,J�7= QS	O�5F�T�7�D$8���y.�H��]�PX>�ͅ���,����c+ C�r<���z[,��m��Rd��a̽��sE�|J{i��b$%�%D�/cuɄ��7 ���q�j��'�����S>���E�+���+�Z��2*�lqT��؅���Ѻ�����!;Ӊf�5:��^$��5��qK`|'b^Mˁ)/��S�l��4.��� �6��tKe�^�bd�o�ϻ��A!�gp4�`|��c�����Ϝ5��$�ړU!��I�vk��]}����b�>8���D��wRrH:"��[�岩�����@}��D�:�n�G�2AA�����E?2r�G{;9��Ҫ?5Ʀ��ST����L��k��W""9Wz�>�`}*�2P�o�OH����gޙ䍌�m�P�X��X�:9���Vy��8PI�Ҳ�����~h�Q��35��#(����e�!I\L��"�)B���a��'�]W`r�)Wf��5�5h��H�2����p���	�@i�Ӣ���é�kȼ�5�,��p)�b�=��խx�(��`�e�ބ6�,�iE5S��<в/u�I��L�)-�(�+Y��T� _+*�6ۯI�ӰԴ�c_�Bw�z����p��ꏚ�(�ǯ]�G�q��x�W�^D�
w�c��gEf�S��mL�%�2%���}���#���m��];�M�b(�b���n*�u�t�h��%�����f�E���	nN��W����yA,�柇�9�}f+��P��@�cs����^M(����2�e�Z
+�]� m�\A�M5S8$�YUU����Q��JFX��gU�s�����O���y2�߁���8pQ@*5��xm����V�