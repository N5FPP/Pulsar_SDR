��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY�5����4˔��MRyp��^�#S5f{�}�2Rt@%��u�8�3�� ��ߝ��@R~o$�d�~7�
K9�z��J��&b�9�N�ch��Z;\QV�?P2\2�̴���sܫ���zE9f�Cf�
�T�
�h�0��a��{���|o:[��DLC9;]�6��q�?�V�t�_)�[��eM��W�@����@m�������A�A�~ܫ �a	����`V��r�l��@����H�%��3W��P�*ׄB�P��3��>�]aAY�f�������O�SԚ�k�&	*7� V�1{Ck��߶�I�9E_ð���4,�g>\Q��&~�;Z
b����A�A��D�0^
��z[�-T����p���Ƕ�T��|��`��
����}� I^"�{e���in�;�����4�)1��V�mX��o�Ω.I������`��(��ϼSh��!{��٘���cټ�;�ģť"�R�Hlp�Ok0j�m���~�$�K��w���/����B�:n~��fm-��(0ii����86bNm�E��|�\��ĳK���Q#�a � ϐ�y-b[�AZ|(�lF��jU.Љ����$��=Y�nQ��Ѳ?����Ni6�)=�9�p��2��@6�6�9��.�u���W)�;G�Q 3������N�_��֕�
AM��㥳��LOt�����+�y�����k������#^�*�P��f�hH����S�	��e��HRbA�ģ�V��£L����S�)�'~�W�N��[��8��Q���<W�*��6�:�`ZP�s���b��F���\��S�O����Z+J�
l�*Аi�d��W!SL��3�az=�+��r������+m��u����L�?�}�u�7H���5�∣Gi^�f�f�����w�ɩ�%3�e,I�u��*�T+4�X��6&����=�P�ٰ=����v?if�8˅��=N�|���߁KFm�-���I������� :G(oX�z�g��N�-��$�>�" �3��9���$�3c�O����mK����e�K��4�C�7�$�k�խ%vl��X��<x}���.A��;������s�i�be`���N� Oaq�j���}Gq�
����/����"�a�nm��}\*�팙%Dh�V�)�x�M����O:bɄ��e���b�䞨Rí���+��t>�����T�x�o9��Ko�=������H��2j �͹�V ��w_.�T�	���Ζ
���J�A��8��ެz��qU�"��Ҹ����Ƽ�_2�D�t��d�����y������h�� 8.dyn�'�ꎞ|Q�GIP�/��O�(���Xo0��S�c9�u���c(����Qa���YaW;$��o���^1�z�/F�ZK���?#�T��SZ�����ӞCA����.bT�0��EM���^�C�;���r�)��Es�-����d����6U�u/[������J�6[u%#�+ա�Bz㥤�Bk7��^n5r�tx�#�^��?*��9���G`L�g묳Q2Q~n���61�t� ��a]��JE:�n��ǚ�jMBҙ�:\\���$���YFV8�Ȕ����T���w)N��K�����K���hO�n���H�zR}��!�}�}
��7P�;y���ּie�>ݤ�fæщ����69�Q�yWH��G\��o��=��z�\ �K�/ɿ�:pȎ�eK���® $I����Hܢ���߲`�6�']�9$(m�m��;:G���Q0�GE����$O�bjƆ��-ŚFM�v3��2?4Y�Vx!�K�/�%�T���*ϲfj��@/f�6;j����J���'��0G�\i����~��O�������v��-����%N�_�pi#y�@r%V0ϷՉ^ ���f�������]�]lg���>L�-<�o�g5�y�[G
���5�4*�֘A�E�.[�p���1���\�_Н��!�ѤT�����d�k:&�،*͹��U�=��κ��S\�9���M����es�a�����n^}��%�����AvA���ؠi㒭�����ɝns�_��>�˹�82���)Qm��@VG���α�F�qKG�1*e�tq-4ѝ�Q�q�U��8��84��!7cZO���T~1ǫ�T�⾑)"�Я��f�ݏ�̌�uZ�@A�SA�'B]��R�8�������cv��ɕ9�ڐa��I���z���-D����6`A"���z��Η�*>������F)��/W�����CF(�`������6�<?`_�ϞqT����?�N�(����v�T�{~�ګF��{�Ʃz��`��-	G�DD��0��y���TK
J��;��$�F1 ~�g�f?��س�s���i��VP̙��t��W[�[���!ywx��h�n-��H>��U�q;,��ުh�y������l��@(�j�CDp7��K��^ B?bU���/�0�!lY܃�A��}x���t�9�� ���RŭbzF[z~(4q���s��l��B�kY�S�4���1�ct"�D�SFgR�Diw�	G�'p��b�GA�Yw_��E�Z�����R�������?+�D��z�ڌZ!W�c�`$irZ2��ftw���r�l`�9)����Tc��@n�`1����{l��(���׎��f����A��wp��O�g�SgJ���،v򉮡8�Cڕ!�9�7r��%FZ�ry:S��k|�I���3�v.�Y�[��R�J��jB.�����N!��,d���e+ǃd�F�e͡��R���ƍSiu�7�Iha��vܜQ1��0���&ֽ��C ��� /�8CJ;��"#�E�p�s�b[LU&��=ĤkA����@Ogn�n��ags�eM峕�������Rz�C�cK��ͨ��2��E�h�\�d,MBkj?,�ޮ��,�kpu�ـM�!�&;E��v�f1ک�эۂF�+{��yl�^ �W1Z�uK�"�b�cF�ɛ7 "��
�j��2�����2��"9�|���;��� &Uऋ�-$!�,n�����}��}�v�Ţ��U1Z:3Ĩ�����"�`N���=���[|���A!�O֌T׆������p���q�-�ǲ`�p̈u�~P\��Wg{�S�$5��Zjk�t�	ݤ�u�XP�/��kj�k]sf����Ϧ.�O&��]�����5�v[+�s�u~5�l���gB���ɹt�y�!��S?t�m4�u�8��y���3�6U�?+`	`HѢ�	b�&;X�q�m�s2@�����J�C��iVU�c:��
_�����n��O�$�Q�S֥2��(c7��c_\��̆)M�f5c��� �@GlK6Q�V)RG����wjG$ٲ�cq���+�4�t�=�W�2B�H�p��=k�"\�e����m\GM���$��|�j�4tX�7�`fO/���>uoK�m-}�@�m�ZH<�\Ü]�v��u�)�n#Eυf��=�1$���h����a���(҄�ԝ\�X-�-xlS�t�����&���Mt�IX	���⽕U!���Ol\h�*֟o��	ќ�^�l�q3y��)e�V@�ͺ7�d�95$(�2�L{�\�K��Ô_��\�@�d�#�?FV+��bL�{[�A(�E<�o��o��ƃ��C�L	 h�J�6��J���V�}��x7	���cPRQr���?nq���sv1dUڣ�H^�P��|�-��%��|Z�ZJ�t"Ҁ��
\�T>$�����aA�(�=�t��8e���w�#z�� G$�*����\O�or��h��'��־Ƙ��μ~��)jD6��@?(���M�Ix��Q�P#��dv�	ج�Y��� � :�$t�Z��5,g���j]ݺ}{��h@�����>�mh���Z�%f;x�IS�?"3y�B�6�a����Z�d߳�t�R	`�|[��K���r_�&��"�v����a"�N���e<���z����jح���a��$�*��|-v�*!�1�K��_������zF�I�|s
�'�F�L�}<��i�ь+Nef��ތMs�N&w#�0b	v�qҪ+ٷ o���`����'�)��M��[\f��~�s�)����WLR@ʩ�!�ϟ�q�V�vL0���f)m.���C�'����j�tM֢kU&y�@�7�����l�F�'!�U(I�g5N�)X�L��(���Q�!k��@*f�m(�Us������i�-%� ��|�G������q�8mG$�N 0[�s0������Lk4*zN	P����)̙�L#���ĥ�������w��"�I<>��v�|�`�s��埒&#�S� �#��?C̱�u[��7+S���}{�凋��f��H)c#��� DN۔߼�K7ȃ�O�G��[��X2WT�p~����ӹ��.K�5�lZ�!3��̊�%�s�btY�^<R!�<L{��U�i���$�5Ua��C"4���s���6 LN�4�,Q�Z_���Ɩ�w"�<��$���} � =G웁����~�["�y#4	b�W��m�����ޱ���d��f�s�$b�6�U�;h�3zr?~��lvO�B����$Mv]�_.�E�s�TK?�%�m��+�L�Q��Л�j.{c��1|E\��2`u/)�g�p��K)`�Nz�AV �n��톝tM�9�*d>&�o�5�o���a�Vm�2P
��[3�2���k]�'�9�-������O'NW�pIwr��4E��-̩�����,6r{H�)�Jd�����vɛ�8%��8��0̠���$C��N�'7̱1�:_�9�;�g��	�<�6^��C5z)?��}��k���b�����AY_�S�5�O�F?��_��IJ�����	�_��.t$� 5�d����1Ĵ������\?��[f����(XA��		�펨�	����Q1��
PxI�W�%��+���n�p[  ��VĠ�	-��Η����j*�4X�̬Nb�-%r�դr=��v�&��C�o�!��1"_�E�����Q1�48.XTH�/����t��𖲍M�9ul0ۏ�e���~�yҖ�N��æZ��g��BD�h�GPP�I��a ��1�@�ͫm�#�,}6�>����]E^�	d�G"���-���7�	����>��l�[����&�+ʅ�hy���Ɵ�����o�e
�3�ֽ�q@MrW�5��(ɞ��%E.l{d�68��0���F��M��쁆u��E
��a@���QM�1H�Q���X�k @i���H��
N�.)��+F�`ZRp��4E�yUDy�g����/��5u����}�Y$���ϗ����I���wEC�.��-��f;Ri�×]��ũ�Yn��)2����!� %�9ό�Q���
j�7����aԘ�bei�"��Ԗ�d餌��0��q� j7��G�4[W1����-� �e	�+ʯ�_���o%hE��Ъ}}��q8l���!}Dy9�@���U��ry��u�`����@�jq��_��ҩ8���)*M&�׀%���[��Ҏ�M��ҕb��R����b"�b)_r��g�u�u���\<�J���lN��򁒀S�3�����-�Oڀe�g�~dm��_���p��a����oX62���uc��:�7!-QUG��@���DO�a���v���tJB��hj@QW���A7}��uh:�^��K�7,f�Ť��iZ��R{�H$֦��ޟ�#��N�:2[u`P����x��c�Oq�Xڮ�x�";���f
�KqW�)j�d�"[*���@��{MSPܒ�.m�c�?�*MW�S��w�x1����9���Ⱥ �_"������μ5q�����<85�X�k[`7+��l8
��J|s�t]�U->��$P:K�"���4-)pk(�!h�v���a�E��,��l�)�|bR��q��j4�_k��HH��>��2C��fzb��	{��6rZ�z�KOY���Z�.�5J��@�ś�d�|+��P�Ū��?W�`��ː9 ��ض�p��DahX#Ip#�N�cl��05g~�?o�;{��y��5���F&��J3��?(6��$OP���0X�d�@�t�M�}�\ON�;Z����	M��dw���ǘ�i�����
/$��z������b8�O;��ɋ�n�h.`+2	���i���L� ���ޤ3�4{)��v�$��F�;~h�s��uG<�8��8�t#��!m!�8������Wq��⹉I#c�F��Z7�j��:��%�wՁ%�9����Y�pxo!�t�ꬭ��}���Y�@��\�Ղ�7M��x�Z�RO"���j�Ya.�r�t������ԦzL��s)%kǎ�<�76���־d`C�sa� �>�f~��$/{K��sU�~$5�nLu�>�5B�@T	[=zGTQ,���O����~bV���aQ�/���G� ��*����g)"{����W`�F����b�tm���PՆ�B?	������vAGEN��VӦ�P���v��r왡�U��$�cQ��Tm��*��&]vF	�4�_\��/�	E��P�ѵ�6�9��8�%�d2���d����=e-97e&4-�%(��Y����{g�� F�a��0���$��W�Q���"Y$���Bޯ
�鲝�=�&q�-�w���s�߬� ��9������3��S���������@�F/�Bm���oN&�~x�
����b�^E٧d�Yk�S�00o�	\�͹!�j��8�e`;�!�}١3>��>پTQ��2�c'+�� ��\6��P�( R�I��~Rd�]���oo�g�%�f��#Õ9���xE�vS����y^Ӯ)r���鱅���ĭ�|]ʸ�7&���i`��б<�N�?dV���{�.-�Z�GI5!��-{���;4i�o\X����Ja���T)w\�Ղ�M^8��yw!�q��B���3�:�r���ݽ��ݶ�X������,^.`� �I�����+Ɩ
��T/�Z(�0�?(8� $�±A�����^�5-.�����Ȕ���F�=��߯�ồS��L��ȤIDg�u�]$�<�v̢����8QUUĮ�H�(��ݒ4��&lcs3�S�zU�o�8���~^��|�KĶ�ք�����d�x"E,Vk	��l�	���Ъ������h�ͯ9�\��ؙ���6�4��U���{$��_��am��](��<Ʋ��p^~�_-x�)�K�4���ݹ1_�;WjĊrt?Y�p��h�V:d�'1�l���|�O� N5��A�o���ŏ���5�BGbW����w����7N��&Fî�s��e��B#�
����}�Jw��� y:>��n8 '�R�"*�a �M��0W���ŷk��E>0�O��;��,D�)�a! ��Fh)u��B��5�1<M�U�
��l97+�ED!~�e��W3��wД�e�zD�"G叒v��9϶�W��@�з)-�g	K�7~>��*�h8M���'�_��2�e.��6��-��W�J�B��c{��/6�|x0����{��*(|�zf�!I�]�Pd^���I�j*}��_;���-yj�j֧e�A饨tp]�~�<a-��5V�}h����	m����j�b���I��]7&���4r`s�Ю�R����aTW<��q��/
5#�p�<J�F�.M!R�Ѝ�s$������Q����H���'ƪ���#��?ڗZ�h���K���8V+y������w�<s��w��!L~#_��l��ޔ����1v�L,�v��:<N��D�ـI_�-������?~�a�*�ug6��O���90��r����d$���W�ov�$-t�v�1��P@\9���R��x��`����=������\���,6>w�aڧoВ����7����S~��(�dS_`��쏛p)��)7(�(�e���F�%@�ȶ���X^4��}[	|��R�-]��Vc�7�H��vX�}�EO�Щ�L����7�גPa%������)�-�]�W�YԴ����5�9��^Gnx�K��M~���^QA���b4&��I Ab����mc�3T�e�&Ħ�e@
��t�U��x���0q&@g5�ri�/\��٨C)��