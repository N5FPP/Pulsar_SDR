��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY������@S��#cb*��=��B���b�
ŬtHWT0A@H���.�v�q���h?��ʜsv 0���?�aFo�}Ra+b'���`������yš	�s9kw�>��N$�����Na9��N�h�K���s���H�}5G�+&g���^H$����q������K�ȩw2t�K���9Ε�κ��UE���(@F���R���Q+P6(.����3�U�vi�"��Tp�F������NoDB �9��f�@P9���C�no<�Սd��F����pc�Ɓ��N\���}�q�s@L��O��}����X���=P<�K��9�+6zK�w~�.�?+�F;J�
���s)��qg}�	��Ȇ��?m�ںqö�5����m��f��
�g$7N�q��������-�7�,�]:%�:�/����D�:2zΐe��M�FX��篔�۹bt��E,�>C�|��8�{7�t���B��1ҵ]��E��I���ȑ��T���p�H��u'(���Wl�{�j�\�L��%������·�;cK�7��V'-�D}���|�6��t!�s*����p�IW��A�|�����=U���V��p����r�"�n�c��]!��I_;�(��/i��ģ%اh�
w8nڭ(w4�h�M&4�Ya��}2N�@��6�t�?�b�"�_������Zv�5�I�s	�Қ«E)xN�|*�$>Fi�L��)\;]�(J�H� �Q Hj��s�,��}�@0�%d
Qi���>�B;��� ����3w�A�*�Y��3�[^���4Y1�{[��(�8#�)i�n;�"l&5��ZrX�L@P��S ��5�%6%��S��#��0���	�^�����t�O���ʨ:ǎ|jy�^rX�pG�����M��!�NY�y$]G�L^�F�j�N�ݢ\<��4"�бï���<��J,ۧe��.�Ax/q��O���F�d܃㡩W�:z��Q̡�ݥS��d��*���D��	����k���������_���2(�����凝߶��J� �IPe^�{`'2����F�(m;��(�waL���I�$;��+&���{�>����O�����`����b�zR|���X����1\��}��70iF^����M�"�}y��K\SFw W�����u�)=4E��⫉��'mN�Ϸ���P#��Tӻ�5rf�,+�#��@��P��N_+{_��A��֨�j�a�/��]6�ܤ��Ѐ�RHRY;(1�˗� �??Lwvd�ve1��eu��2���%�Y�R@��^/��[��,��;A��=Q�[��k�O�H�<��|�vg�ZtB��iҕ�HLt�������w�Il�0��7�L��j�&f^�����Ll,X-�R�.��wO��6���{��k� 4�mz׸�J-�זA��L�X�Y`��(�)/�C;��&�R��U����h��U���f�T=�p�ղ�m�/�: ���9F����3kR�[ڀQg���1u~��c�Ҏ��Zaf��'㕸o���{jqG"�^e8�C_���P����:²�&8C���������vy^B���(�_�N��m��;�{��2�B�4��V�ۇ����VD��j���`�G�q���{7WX��X�ȩ�.�f֋ԣ���i�X�i��,��$�h��j��f�Z�xk�S���h!,O� ���Ԫq��E��E_���w4�j������\&��O,��\����6�	R�f���u���`�g[[AV�c�
�>�M�	�ĕ�L铲v$��f��dq������y��MR�๣�mW'���F���{hht��8Y����w��&N��J0��4y'8��0�_����6w�������X�Li��:u�3Q#lK�l�;' ���Z��mO9:5p�6�
��ih_�ٙ~A���'����~8={!���X6�$r.a�ɘN��EU���p
�G���Ϗ�P��)��7�z��o[���Հ�2��tI-�kh�[뉲7(��߲��1P�߿/�s1>�<��n��/���>���)��x{ƍ�>Yhj�Pe]�;����Mq�ϧ�KA����*����:	�}�{��n��'*�sY��U��oW��=ݗI�(.�H;�S��Y��'j��)a��~�퀥2a[�Hg§�̂��F�[p�����!��Pt�
&.D;�lM׏�/P}�$�i��gZ2���$!�)����mOq�8�@i��P���}�����\�0���E�4�?��-�:��M�Eꖛ�gV�9]�±�O�j�#3q�8os�v��y� N�kp@ e�_Pg�Y�ڳ/]��n���~���.��)�0KF0���7gk�/��\����$�����Z.��(a��P��{�)Щ�l�lMIc���J�4�I^�}B�T�=0� �T��Mnݶ�8���W�h���[m���ys̄/��~Ċ�����)k-Xw����n��'�8g�	���]�&'c�V~[��ٶt^�;D9�\��X��넨V�^P/+�큕j�A���P�شu�Y|��A�����QVm�S�(Y}�>T�����.*�34�M�f�=ƞ���'�Ǩ_y3�t�<�d�;U���[.��~�����'��fc�bk��=��S
+e	.}�qF�^�'�y nX��N8յhI͊W4��Eu�*GA4�`_"��fZ��k��[�A���h��Y��|�ʜ�Q��Ո�J9+I��E�s�#�M-�a|�f�]��wj���%Y�	\�PHѵ�?�k'}W���.�l��ྂ�U��.	�P$'�K�TI�4j^�Y.�o�h���~ 2z�`�<9Wϼ�<
p7��,=jAW�z���jZ��z�W]��_p�����5�$����L]n��+� �(0����C��^:�VK���q[{�0ʺ�b�a����gS��)�[ڗ*z�F���~��V�WgYw���M�z����zx2��Ă/�`JYB�*n6�.���a�
����b�ߘj=�����O�'�vjx�S�� �&�{Fq�|3�K侾f*���!�<���_b��m�_d��=YQ�Q6�s�pj��@-�m&�yvH��K�ra9Zu�E����A���|��"t���]֨�d��]�2��%���I5��}V���7q�zy���f \	���Ƚ0���-�Y�HP)8���R��K3P�j]���
��$��oL�s��X��|1)mM��'�`�I/K]��l���>�
�E33\d�����,�Ks!+֠y.��Y}����++�m~
\7�R��{��Ȍ�rg�L����h�+��IŢ.e�j+��w�T�-&$y���d�L�4+��i�ݭذ�~����J�_�;[Z-�%y=��e()�$R��H�9[�e �?%u��V�FS2ߕ�BA9x�2|���GX|H2���^O��"�K�+�4b�/��(�Պ�=E�+}��t��d��Κ�`��H� '�T�s��^�5l(�:Q�T`L��$�c�D�?�T��ye]�V�m.�<�( l��А֖��+�0��<� �^j�w�[���BQ�x�)��ig�Ko�A�V���E/�{'�ي�����*�TUl)�ج��1�����g�
�j�h�=�s���ҟ�bܥA0K���z��(��(����^�mP1u��-Z�l����5G+�:���6��0��jdf��"5��>�^���=���6�)̷=tW�LTq"�pLo
���in�\B�cM������ǿ�Ј�G�2-���]���<�>���[�*~Q�����r]�Tm� ��ǜ �s��{Fl�Gy�1�%߄���}�>��]��a)\�:�������T�̪�%�#�5z�Cs���F�be�~c�ͦAf޻�A���
/�8R3"IT4#��I�����9M�>u���.��:J嶀ݳp��$6��'�,��4���[^�`b�f�g� `�Y�q�r�<\_9[� ��KD�&ט��k��*��pŻE���4jf�U��ʞ���b!Gtp	����=���&g����%���'5�V���k���x�_�B.}�~�ö�\PL���K1�g����|�6k�����J,�w?'�XSm��,n[.�-�ޕ�@��H�U��چD���D��-�x-�|t�K 6��[OР`���ӓa�SB7��~��]��������t�>e��~>���(�����Em�a�\�Sp��&A�C/_�sq�m۸�P0<�Z�I�o����x;C�R(i�ST3r�㟦�� ���C�/x��c�z�B$[d���{S���&�b�O*�m�C�Ba�%�F=~ꯅ�/������]�{Um �z��E�7T]$�/��H����`>�D�3���<�j�񿺩3��9N�4���\"Iؠ������=���$�� =J��Y��c�ZdR�:X��`�	tl�����<�mj�'_��
>H8��$�0���'K�<w��%�8�~"N�a���';rL#C0a �<_�8��(���3u�N�O��)1a.�*���.�W��u�E{�j�Έ\`�z�|�,!�}9�L��@ۜx��$�+�/Z7q��P<���mn�=eoq�Ƣ�5����˷/��Q	��y4�b-țV��3T�+FI�tɼ4�N�b�W�Po �I	~�Ys��sm��8>-"�@�+=n��+"��`��5�#4�zM�%�~8`�%`�N�D���/�n=��%X�k����ȓuh{���D�:����[B��K�]��}���O?�t�A��x���tݴc
T��"��zy��,�l��'J����������(�)�C���^��Y}��V�� �V)aS��8���80&�#c�(J��B�@�T�-�9\��7R��\$���UU��E��u�r&�s����" ���) ]z����,o�¢��#J��╻����I��N��>�`�F�	氕)r��N��m:ݽ��8�z�g�@�4�;(�F�����L4�U�/8�=G��A�	���Qb�U�y���&�R�5���B��6��P���tN�}\W`윜3�rb���*�����:���YE�j�c��GK�e��Ȕ�K¿S~r+���zj�R��СVL���|>���k������XVu�6&�Ύ��3t�����N9��)�9<�K�+!(��(-�ޱ[��}��'���.kpR���&?bY��x��������+��w��g�l�RMk|�i�d9Qf0Z��)����H9Ab=5ҟ7-�u��靰�9���<�z�L�;��e���D��ޤB�'��O� �}־��o	@y���g�yY+��[6;��YN�z���?�_"L��^��<����q��,�)�4ZmL%�M�U��[��lSr�2bS�$�����u�ıS��G	��a��C����~�.[�3��HTP�5�&Q�\k�TE��r-�k�z�{#
�t$QO�BG�����ԍ'R7�.��esp5���u�X.�?aI��+�O�Z�O9������<e�1�@������W��s�	ݯ'�tP�=�&�{�;�]T�E��Y�&ژ����E��-���,*�8P�.S�Ё�w����s�\R��'�}pXr� b�?��8�Y��ڢ�of�.��0C>pƤ$=�0=���<���S�¤l�_���<��3Q���L�Q�S�]��cB06������;����F%�����7�K��M������~���M0W{�ͨ\��/J�����o���y����r$'2�8>��	K>��
����2�A=>�������.����ƀ����^u��Su�\����0'�����@��m��p �_|�Hɉ%v�;By� ���	��`�%�C��Wut�PG�}�kM��O�͉y�R^�޶���!R?�K����H��"a}�X�n��֌V��c�V�>+��8o�&?�qC���xVisM۔-o�����Φ����|妰TRˋ�;��ۂ��;�:%~6Fh�����$v���N��Ͽ>L̈́4��uՀ���gJ�~ �h
�K�?�ܱ��h� �~��2����	���D�^U�l�9~��|���"�����ӛH H���Y���$Moͅ��+y�'x��K쵋���a��S�~��:�Ƞb_ݷ 4��H�'\�l�[�G(�7��a8���y�[q}�i@*�F^�.����R�>J+���M���}1�0ҧ�����e"-]�z��`_�r����>"�b�?�:4���~x�Ǥ�d�j!*~���V���zᴀ���zNT���6hҚ�Fp�� �I��-�H[͈~dO�ǎ�P�K1��}��6-��1�p��0��¸Z�^C�5?E�5���B*�k�w�5��.�rn�P�����o�{����DΠ����vMT�Χ� 7�� 3FdX�yj4 �^�4xSd2�k&BȪfo.p�.�����Wr���Gr5Bl�ߎ^�� ���,\�؈c@�p���2x	���D�E���C���')�c�K�f��^PU��W>�Y>������6u��;δp�+��sD�������U���<��G�;}���RߐB`E�Fƿ�x�dN	�@Z�y§�D��apՙr"Y.��cI����3�˳����Ɛ^U�w�͕ި�c��z����3��/��犤6C����a�NҀ ����E�&�G�S=�V�\�$���Q*,�)��c���=P�@d���O7Z_�HM80��zH8��S�Y��	�77OJ�*K;�\ ��Z�)5�a�&��w�<3�GP��+?Ϭ�<�@��L��=	,��y��_C��s�C�;j�/�u��X����T��[GѦ9��e3�<R�`�X�kW*t�Z�^R
s�&��ϣ�*`�a��Ӻ���1����?�ݧ�?��e�B��A-�w��8|�D�/@B!��W��,ipު,��	�5��%���|RG��n������g~c�`r�Ka?Cՠ�\n�Ɵ˦;�[�x�Ⱥj�O�nѨ�N#�%�O��1��&�ìj<��#7��Zx  �G����Q�	�`QN�W�^�Y4@���u�|�!�Oټ�zQKϬ��!-@3ЋjдMK���Y�	�C��N>q�\���|��Ƌ�U�f'OT����}2�j��u`��{�E�ƌ��PQ�C8)W(c��̹Ho�F��цP�,��#�n��c�yѬ�����k6����b�gEj2=�$f��?]�����ᮛt��K~�kj��zF�ƿ�$�@����)!��)������En��x��I ��7��+MsjN�tK �Ԛ�NBp8��{�o"�����6'3�^�t���
�����x��g����Y^sOC�c��DTs�mI�Id�t��R׵��͵V/�%��>�7�k.c��%6~o���,�`����ȆG�������1�l�O��.�P���uD(�2� ?���%�qG~��YJWq�7���l�W�E��L��[O��gE_�m�?slٻ���.a�����x1IW����0X)�V6==�[kp�i�TO|9���E���+��NU(&\�H�Zqx�=D
\?6�У�>�׼@YƁ�ރ6|�4�e�Hr;2�r�d�5���2�Ț[0�jaK�Xk۫��,��T�(��r\�}���uݮv���СƣyZ�
G"�rE��܁q�z��z	�O�MN��=NcEcrbi���d�tz F�$�̟��;|�W��B&R�T@��M�:�_��O�6f�󺌝��-�mI�����y�Ӯ�KFSXVv�]��E�� BM'_q�����I���EB*p����W���T���1�u9i
�8 |�o�T&��0i�.��1??$ 6��>S�2��uą	�S�)>��Q}���J;x���Û ��a��z��57cU��FV�]��O��쳽�]�JX4��C�UX/Y��p��%d�G/Ԕ�;d��N`|ܖ^Ͽw����atV.T��;
z����y^.�t1��Y
�:&XL$��P��S(�� ^`���u=?�&%r�.�d�-e<��mQ�h�ke�۳s�R�������<�[-��U=�T��6����?�7+g�=m�`VSf6A��0�P��7���:͠�-;�i��
�&���I7�~��6$����$���Q�f�a��B�l;{֟tUT����[�����d[C��u`}��d���*�wr|�D�ݞ���	NZZ;ϊ�q7���y�1E��vX�ˊ�h�^g��33�cۀ�)˲yA�;���'�*�,{H{炿�n��h��Y�����ϟS�J�� ���T���_��ݟq�)ß�殮�����ê����ܷ�d�܌�J~]�/Y�8bar�L?��64��ah�c �h��!x��R�v�s/'Wgx���x����S�t ��z���f����Ɣ+ƺ�R�:4@�$�Ǹ��]�.+��W�Z߇��5�!�ڄJ��ፙ�
%���.(�Gh7l]�5n+�@�+�A�L���hX�<!F��ِ�I�B���5�2�	*Bűa��.8��v �HV�6��V����1����~2D�˂�$]t�Í�IF�~^tBOZ(צ��c�9�^i~hm�a�h�ͫ��0�&�5�p��!����7q kz�~*�;.�&����{�_�s�؊o������1&x	�z��Ֆ�?v?�)�&�����8M���a��Ϻgo�?A��4��F2E!X�����.�.�C7��'uʵ9;�#�s|x�]y�����?q��^�^�Ŝj�N��Z�p=���8�� �
�,�!�k�uh 6��tF�u�&*(����,K1E�8���`htɵJ�\Q�P �4��{t;��ꟌqZnT���ǡoT��ykM���y�f"E��v�ַߕi_D+s6d�w OA�`vz9e^���g�8��%Bhϝr���-�_[�o��]H~�)�˦n�d7��4El���M������R����^�~4����Y�;�c���������B�������C|�?�G]�܊F�2�.��A[X�3�}��G9�E�gǛԒ�7G�M��t.B�O\R&4ݟ4���]�'9���[����R�;�T��{����6hxrkwPx����nL�Ҙ�Gd�c[�r���P���Oz��3�=(/��;�Cvň��M���d3`b�a�Y�����ә�l��3�2�V�QaK��ǎ����9�S. ���`���H-�V�)�!����%�|<c� �̛�m�΍ǣV�מ�<�-C��
9 ��˹�XA���u��O�O;�;�t���*=�x��������,>V�Ǝ;��apr��niL�����[����>�ޫs}D��i���|.u�-��g���E;[���}� �SsG�fg�g�q1�<9ew���O*�H���\�"�E��F��
d1/��^�^�;�5�7�z#��3]����7��%%O�tV��o##S�Y��4��,�0@����G)����ǃ����M��#�����)�e'�y��K}>va���lTF��;`�fƲD��@sU�>I��U+��]��{�j�l����^�V3��˨n�X&��n�a?W�/��"q5��r&W�HyH)����1F���3����e@���@�u��#<��vJE H�"b� |��{���4ۈ�#﫺 D��uc3Iu/Yk������.�W�Tf/�(��+9Au�X�����j��IM|�`Q�O"���-��'��9��q�v���o�!V'cMyU�,a�J��$<�31�� �#c8�6�9����FG�����0W�Ϡo�Z���om���@4� �ؿ��^�[��YҀ*nEg&� 5i� ����.��s�[�u���C�<�������F�  �!��7Q�5?Iul��0$U4���_�e)9��¡Џ��� ��-��~ZZ�ǌU�;���!""��h
&�S�f��H��z�R���F	�@��w�2%����\W�o�X$���Lr�w��Z"	&#�H�}6�=
��3�/�#R?_��{����oc!�-�&q���EFS�@0Z䕥�#��,MR��?�x��)�C���Z���rm�zX� �sW�\;˞-�cm$���ǋ����9��5xB����������\x{K
�i7��Qr3��z�lG�*Nб�L�]D;`��0�}��BI�"��:GWC�L~�ʽ���k�|p.�d�^�V���_r���/�@/������ ���a�h�-�'O�l��1֏p�/[-&~^@���H��Rcː���F�[�����'�?�W��A~F�\L�2F�FULC��Fy�l��8��p�Iŉ��(�y43��_�'���_'�J��"�Bi)s�]^��1��o�� ��Q�B"߹Z_{(g�{U�K��z�f��x$fXre�����W|�4��WT����ƽ4�LC��p�s�A���=z5��pK������րF�0A�t`тO�QB
�TUk�|v����vp�ͱ`�B*$	���3��ЦMX��;T;*[�l��J@ �R��>��<�z��/�s^k�֭�,�6zs����?�K��:�����i;��ءV|�yCV>�R�Y��hq��Al=`ZG�W�@.�+����u_��^B[M��xǬm7²;]GCc>i(v�uz�)�5+�_��
�Q��~��rs �z�@֬���DE�
�W�������kz�c}��#:[Qig��B�q���f���lw�cY�P�.9r����W�)�o0����?��mA�D���7X5���Z��2
|�n�g�5�[i�P�f��A���Y��qz�_1�(�����R�Q�#'.Y_Ǒ,�� ^�G�߂C�q��Q�)�W3�3QZF�����ot��+��o�P�������D�zk|P}�n�12��M)�f�������6��x�,���֜/���Vw�X�#b���&����:>~�Ku����x������_�1h`W ,i��+N|�2
w�5��k�f�pS�&kGt=�����+jg6/���aK
=�l+�bʼ�1�i���3�XψG�\Vh�+�{��c�ה��Jv��*�*W,��Hn�/X��,��~��xV�#���v����F��]
�)��w�Y[
�(w(Xj��"����w,5��r,�1k��$ni��'��L�D�щ�?��6퇡M3�Rn��oҌx3�rژ�c������������6Y�� �9A?ͺ	�m�%MD�G��o���z:f�W��r�΁|�w�ڲ�O��F�^O$;^�-��w����;A�>2`�>���TYU^DV���e�s��7<Ŵy�C����1�^&�\��m��E[���4%0+�b6��c��'l�>[�[ѫ���XS"��HZ�w���#uG.�^qJ�� ���[Hx��$טb��4��]�Ճ�eMb�?�{�УX�]U9�d2�X�;�*L>���]�,t���3��/o�����~s�K�/���yw�n3�IH�Q�o�D��2�:�ܯҏ�8L���d#$����Vh �G�Z������A�c	#�ulU�v�y��ƙ���͍IT��A�t햢^&	,�T����@ElJ� ��	�]�X�~���B�}�ړR}���HП=3v����9Z_3U��d,Vz�ٿKr���b�������j��IU[3��Ur���[�r�	ް�����1q�Y���z߫��%����S:�[ޠ�XC�[�ό>�	�d����!���H!�Cİ�0�ѳC���������Y^r[�fΆ?�_&�b���'{z�;�mp�^)ktw� ̴��S�1��Ɓ<�7�C�^��H�2T��:�����Ӧ�~�,�+R��ɕ�,�K EH['�$ՅY�m���m�,���������w��oO�~��t zf�t����N��q"��*lD��ͧɔ�e��_���K{�̚��<q�M0f�w�����@J*�:�1ڵR�j���M��l���O���Ox�f��V@^���$ns�w)��~&7�Q3�m�r:!�p3E��||�Y�{�_G/����6���̸�;֧������v����ʚ]:���}h|5;��&Qk�Z"n���c�c����(���7�ך*����� �G�F��S���09�Ae%-{|9�����O�L���4����qK���E?'�=� �[��Ր��s�d��sV�L�DM��h�_��'���ru^����^�2D������}�t�� ��M=J�\�p*���X���cA�b��b#���6�����X����#�Ra�����C��t�R�e�L��E	�LJ���vI�><_�#�rF�;�_T�3p0�O�3ab��#�!�+��g �����y>�Cc�&�4j#}=�{�-�AY��!3���ZÚ�Q��Xeɲ�瞙��#
�g����FZ��؁�J���X�Nd^�j��M��+��rB� �Qh���pˆ+E'* 5����=��d2}$�rL� D�D�?>�(�����%Q��v�Ae�d{h��F+���Dg)���|��k�ؿ�o�|��?4	)��I��ui�b��k<4q�$��۳|���TD�VE ����SZ��1��K7�F/�s0��v'�WfK��4��琏y
Q򦎛��eH{�{��� �X�/�Ǆ�4��ʷT^�ωņ��[����}�S��H�š��V6��!'ab�\!��5��T���xn�'��U^E�ʏ*�\�s��	�Jm�!�c	�&�'b>�����c��b�CGR_�ꌞ+c��G�B�Q"�)�"(&1B��Fh��*��g����h�T�O��Y����|k~�5|C+�J����}~_FI��)7S
0Mu�VC��	o�B�$�y�>���H�5}�J�����_x�P���YA��3�+�4��\�˦$Oղ��c�k2�;�W�u0+�@[|<� ��z]�T�y4�C�����eE�˶��Rq�歕��3�Py���G	��{�V���.���=�dXTd3���|������%�:�k�u��d�Y�g��f �������*�����xt:��j?�vR��5�U.&dVg�I��O�cA��?��;�ѡn_�1��w����@=.�����0ݴ�@ɂ��R�i�b�-硌�jv�ڑ�Ŭ��0f��KT��	@~�'E	-�暠e�������l��Ȇ���pf�~9-5��7�{��[A�)��3��6l���5���B�d�O-��9���
�H�*Cdm�ka+����wqʪ�Gv)�8�.ao�Ʈ�-��[��q���7;�����ZR6�_�1�����^����&��a�S����43����)�i�+:)�F�vI�	3Ǐ@��.�-x��E1��s�[-c�W-#� |��e���R4�S�9 �.K�+��Փ��vX��ϙ����}����ܟ�>�t �Ć���Ժ�@�M�CG���V�xg`�3y�N�b�L�/��Z�%�5����ڝ���֯p�{�t)BlC����"��(�����M��%g����f�^�>��������dU��%urT�!�x%ZNq�����k@V��g���&6_�t@���H�������=��FD�[��{*��^2�^mOF����-&X�r����໺%��*��~�U��Қ]�х��F�
|Q����t�Ro��;۲�:'�wd������G���#�����w%���R�s�UL�^6��ܰ҅ߦ!���f._��\`��8Vo�F�٥���: ������G
6��rY8:3W���N�T��N �<��o�O�x�ze���t�{��K��'_z�"3ԧ/m���� 5��� ��4�q{{��v݈I���x�#�nN���B0�
��Օ�!yՐ���D!��7?j���䞋���drU
}¯�u������5:��F��ӵz�l��ǲ�k��:�\D��<VO7CL��¹�� l���`�2�6VB(9Z�O{������D��5Ҭ�Jf����A��Y�B%�jklB'����5��?aBk�ǘ��6l�,zpM�[���ky�A���z� �r���Z��>9���e5/��!����w���1�]0��UM��z����M��.����v�M�EGK�=�)����������b�y��d�ar|y��9�ڲ���a+����Lv���(� �� '�Qޢ����^�'/���=���@��s����;���O�a]�N����va�%d�ss�Ro^ (�r?��Q�#9/b��;�2g�K��6�$Q0��\�J�!;�>57�.!,f�E��3�NL�@lM��}�n��s�I\ ��t��+c>�Fj���XCN*��;���{�{�5XD.�}�K�����,��������t#haf�vw�,/|����J)����@�*���㠏�,� D�0 �Wi��d���DXuG��WTxK�����43t���� ��)�f���Sg�!�:���ӛ����R��3Z�@��k�4��,�?re��ݎ��R(f�qhi��ӊ���+��ظ��S�@Y�J�1��o�̴�WeQj�C�'	aM����γ��d�pm��F���j�ߚ���2�,��d1n��& ��t}��9`�^6Mm��vT	C��0��o��~��Ŧ8�+�B�� �[�[�3B~͎N��	{١u��u�:ϙv�GW����&����A�=����u�X�A=GD���#���R���s����+[�;�l>/y��F7��F�m/���X�t�k�¤%U���d�K`!C��������r�1#'zq�y�Wy��p�rR=����TE��f?��?M��&A�-��RіbP{3]X����'��ޱ�=?�?>���s;��s��@�+[��']v|�2�Ć���Jy�A��{��0SGsQe$G��'G�C�0�=��׳�0����Z��\�5<���9�,�'Q��N, Yt^�C3u��^��3����󎻖{�=�"!��j��S�����V�?<�7�,J�혟���%U'�����=���n��ȪL���Wh)a$�����X9 T��Ae5��'�$7F��[3�é=�JO��C�|ӥ�?7z�J�n�I�1��̿Ңګh�x A� �u���R7/�ʶ���߻4{�𵨛90,L`^��T���%�q�� �{�S�����	���~��r�(�y�BD��(�z�R�F�1g\:wXt��k:_38�h��g���$m+/��V+{}�_�	`�`4n�k]����[\��M�ǧCOuP���/��nwJ�0!�*wtid�a�$5@�J;&b-�g�v_��AD���@�I֊k��y����K�Nb�T��iZ�V	D�!�v@P��RV��c{: ��G�ZͲ[.��ᝤF!<[�<H��N�c7���P��?�X�/^r>�K$�B�Z<���LzQz�-&�����~ӀI� �B�l�%Sӌ�����O�v�N����Sz���,>ŪO�>H^\
����Z��=j��7>L`��2�.ÜE0T����J*W�kF����m&�̖wo싓�v���ju�)���	�\�;�wR�y�l���ؑ���"tj;#��,��,P���������ذ�����cѬ,�D�;E'|݁q����jg�G�B�p=yԊ��z�
��Y�ˁgs_ZmJVLxJ�d�is����47�L�Ic�ObS��z���|?ᄍ��2��N�̮��o�U)�Pq���6G�~^�Y�R�P�8��<)LP0X�#�m*��3X��A;$#��\�Pp�F��}�<��@�X�u2]��dXM��؄s@������9��TT�S`R���{+��Z������%3��V��t�M� ĳY~9�1�����8���A��~?�J�:�6ab��}D|�C5%�ă���7�*�E(9���_M2ܭH�;աg�)(���w�`�_��~N�,�`Z�����Z-���+��;��Z7��q�}���؊�'����P`�o�X�r�a	i�ѩ�-�Aq���p�q�6�U�1��{2�K��Uw����w#D�d�ͦ����sq��ģ�چA��7�� |�����L��&We��qg:�3�D�Lk�;.I�D�G�D�J�W�+��7W����i�qRy�@ TXbmm��ɷ�"�����NE@�s+Q8���pڬ��1��D[��hU;����(�p�M�/1���2�����>;FJ�}��b?��yc�C��v���s@%rG����+��өd�e������_KE��9����N7lɝ2��V`U.��*M�K�ik�����'ہʖOc9�U`h�V�L�ſ����X��i@��{X�Q�M�T����:q׆ꮄ�y��gUKׅXV��a���+"�z��z�]VO�ϰ<�L<.�I��̇C�MeXj��.���Z�Gi��A�ákم��¥�s�s��f <&d�g�ˆ��'�+=��^���:2�S��� e��ѿ�G!�{M�D�>�x��W��V^;h��N�)��?���E��;�ᳰ�q�Wl��X��P�8�̰�A����Ć&/Ũ�>�c� SlSΧ�E���53�}�}3�?��_�"L[e�tk�f��yO<ʥ<7�� 4�b�Rl�*�J ��x��,��-�o��q·ݗh-�b��(��$���1M���A�R���?ǚH���-�h�9,�ÖCY�蝁N���z�z\<�����6V���ߖ�d��9�Ȗ]�e�\�OQ2lp���$�z�^M��0���c�AVz��/_��Ľ�x�/"eٞ�w���`��<�4�}c��
JJ(D��X>�Nr��e���۽j��"��]��!�B@',�g�V87_�"l	܁}�i,�'�A�0,R��JZ3��!��SpP#���[��r�W���@�����v9�-�_
>�>$�2�A�`� H���f9*`�bFT��tg�9�G��t{�l�;����,�\�g���r�n�d�;��-A)K��g������f~�F���	�I�yp�?1_$dy���y�+�$�^n��w�7��������֦�����#�KǙ� ��� �cE������F�HM#�!�}[��EɖM3��O�V����qJ[���d_��S`'��2����e�vZ�b�t$�# �+t؏U�0�{�i� �{�Z\	����?Б�-�
��i��W��xu'e�R�/�5Q�Gq4c���7z���V�C�m�(r�{��ݧ��Ia���"�I����i_�� $V�����Lc�!=�ޗ	�Kl�r��~�邎��@AV�r�~Y���.���mz'�2pb��V`O8����?q���=߰��g&Ȉ�fx͈��pO��5�ܕ;��{�+�UB����cr �˞��\%�;��Y��v���(��6pu-�vK"��(�\ ]лex/�F>,4�^'���4nz�6X��E2ۆ=eR jz���$�.G;�7M:���5�?�����w
��*�X������G�+��	�&Ѧ�6V�L��!��Ȩ�9Jߡ+(lԊH,�
��q���@C���3΋3~�=��ԙ�R���M[�_Bř��r�o:\z��]�ӳ@=�9�������]�*�P>3ӺC"���Lkޭ!�eՕ�FVX4��V��>r���t[
��bWmY�0<oQ'�{��5�b��
s�vMLbdt�e���ן5�R8^*b�$�|��7�R�˴�Sg��֞�#��fCu�E���X����헰@�����Lz&#$y��F��83aj/�8%>T�.]�@�eF8q<�8��w��e�g��(R`�v���V��g���@�U���A����������Un���A3���>]���έ#J~�6K/� �^�c����4�w�x�Y����5�h#�b,�(6�	����6
��¹u�B�g+4��W���ֹ�84��2�@T
��n���y�j:B`K�����,	I��ia�/�w�d� ��鄷�E��2h����{���^a�[�	�ݧK6�s�߬��_6�
�b
3���F"���/G>��ɪ��X����l4�r����*n�F�!܁�`/Mwfl�K�|D��Uv�}�7���]�O��Ξ�"�=7���4t�?SWeo��:+8��"W6w��Z�����Il��n�Y4�Di�O �Ԯ��6�H ��a�Y��@�k���҂���jr/x(�>16�����,�6?�xƴ�������7C2C���{�s�,����zu��쯼'�S\���ŭP�7� �ú\)���1Ǿ�%4l������hb��Gr`�Cj¬�o�x�=�x^}s^jc�� �}*_�����m���׿��ח�y܀W���%D�z��CN��<�N&��WeӲ���Ը�R\!����c�$���:�������E��}a�E��yi�����W�zR�]~A'���}�n/��:;do�V��M�V �48�_��O����l�䳙���k�V�/~"\	��ъ���q���J�ע���۳U7�;��Z0�VoA�<mJ_�'{9)c�Zp�E�s�^ڔ'��;|�:E���������9pseb���I��c@�1z
�Ѹӿޫ5T̞��i��q�/��'��m�1
�r��=XA=��0����k~N����2�7S;�q~Tu�gQ�W��g��#���k��Ԋi��È���΋�$�o��bO��
.������'8��^FӶ�3ɗ(��dT�� �F�7�����P��=M>�N�x�n�-A�tE 9ܬ�F`�� +������(�����J����0�/�����^�����FvP�{Z,�+>�F�ܩu�<����Kp)���`n\I�z7v,��*�((0�go�)!JS�S�n!�H���K��䂯�"�Z�:`I���&�T5���z>���WN��M-��?­�X(���Y�k-��뇊�'��rg�q�Z䊾��`s��;/��Usֿp~��|�F�X��1 L��]�R_MIh0�'���??��vq�T܅�A�ө?C��2�$��4U��?W�R�E(_�CXw����L%t5��o�d�u>T�Q�猔��E�������F0���].���~+s�ܒ�bdl|�P�R�&h���F�@<��C����+�X�U��Y�]���7v��<в`b7R�K��"�R� ����nAڲK#��&Oc�,C%(|0;������'����v!��"���i~�+/Mk\+m�$�P���G��̦��Y��o�����xn����'�	*��nME��_e��7^
�g �v\�:S*ju%�?���IM��V��&s>q��2ĥ�"hm���̂�n���ރ��Y�h��뽲R��fcVX��b���Y.m�݄���:ʾ�^��y�{'ŕ#�!��X$S��vte�n��*&���w���d�gg�F�0GjC�pd$������-�7�mR���;�;�U�Rl�|i8Eh?��7>"�~nj4~�O���B ��ꉤ�z��������ka���,n�$$Ct��E��=A�SF�BPj/I����}��Y�%���!����޾�����w6�H�F��G��M�9
��FW(�w�u�K�]u�:ɖy�;�P��Z ���L�B�ه�p�~���T���܄̹0^���NXs�-��8����>c�Aw�׷���j�$�t��᧐���<��J8PrQ]����#S<�N��۪⠅]�������F_��r~��(B����n�o���f��+�8��~| ��@ĥn �L�y�s�W,7�_T�t�]����#y���[ꭘ �ۜ��B�	e��������b{�����Q�p5�~Smn�3�x*�+�����[�Z��R4!�V��g�d;� �ѣ�ާ�����Cl�K��Z��3��˘��7b{��ЯE:ִ?���Q��O(��0�Cd����X`�t2�JP�"CQ>��#�,����PY_�M��qo��~�(�� [��	�d�-�~��7�u�$��."ߛu4|TvbS��7z˜jf�'��t)&������)g���z�!v���$�g�����,�ŗAUilN�)�ݾRw�x�3"y�y$PB�����yT��i���� ��$[B��K�/��M䅔)t{6XE�2C8 \��L��W��=�*���3&����R_(S��Q2�����'������PP6��+��&�蟐M��Ƅ@�RR��1٣RԉN���4+d�6l"��1��� ԓ�M�G�����Z��q+}*+���7�����aA�(��Z�g?h��aݴ~-m����8�Z	yeW$���a
�jA�0?�M(6�?�,���>Rշ\�E�SW�̠ٟ+U�<��C僘�l�������$U����@S��"�-w��JLR,���|�'���ݴ�O�DB�d;����ڀ���';��O��!�h�	�jJ�SF� A���� �-г@���LB�7�r��V�h������9;��i�Gȝ�٩e�㽛���s_������T�� ���8��Ct}'Y�c�,�:G�%~(`�Y��X�7B�8	�h�=�i KжWx�O�N���'�I-a��oH�8���Y>3v�*��̓!�Yd�����lƯw�ӗ4ƃP�ʾ���Z��tT��Ȫ|Z'�Fװ�٨��Һ���U�l���Ƞ��c92v�.J�lfN��JH0�?�og�Ҋᠱ�O^ͨ���mҵ��\�D����^��0E݆Zʻj	Տ|��**/�<��u��y׀��4����q*9A�u�Ȳ��M_�����Dmz`ņB��j�5�n�H���g�X���E¾����Rf�E��97�⃚G���\�4�qT3�I�O����G}`u�v`�Yﲴ���|sﺍ�-�GYd'��R��	�h�|��bE�I8��~�a��dORnP�ovॳ9d6�߾�H�D����J�=��&՚����<��z����"�\�N�#[O�Kޤ(o�Di�1�<��dN��B�[�#�y��.)���Q���.�Ü��ݶנU�=�� �����&sh�+��z%%�@{F�WP��@��f�� &���Tp��	/������/�l�N���IB�b �0/�h5��_.� ��V�-!o0S���zĞ2g��͓�o�����4����6z�&=��ȏ������hSM�$�����8�~m��-���ʻ�4�v5�B��G���R}��S��E^+�՘�v`���W���_��T.ʬ..c�� T&j�'��ߘZThr�/��M�e���8�&�K7��0��N�6�������Zc?JAw���]BR�~�����V4|-�#@��7*�&�W�k�Zk/wǤ,��C��>Lv�5����g�V���$�D܎�_��Zΐ%�/%�u���l�:h+�������J�Eqx.�&�?����,}�T��N���+����cv,�߆}�z���Qb��U<3[Ӫ 	g�� 2���.��"ҫ<�xd���Y����H�F� �y�=�E�6�k�]��H���2���5d�3���u��y�� S��cz�^ȸ���?�=�y�� 2�>!�69����K#�N�?�i�ӭ1
�F4���3�W��>yLs
,X��2�0jcDϏcI�#G�v�#k����L� ����ǸI�uOߊ�֌�{���L*T��G
c엾g��~vC�B���L�]ru��w�c�ޚr3YȮ��@� (�\ֶ�alR��=z}6���!��4�Ȫ����Pkr�A�<�x9�����(@��k3�������/��$=���r+vB�%���S-bs��4�-�x坒�8(��.�Ĳ�A�$d���vnb�)U"	8���N~�	(��R�`���"�jHE�ԭo�����~Z�2�T����P���l������н=��˱�Q�Ĉ�ht� ���d�P��_���ftO��I�ͪT�D[��1��F�G��s������*Ho<jw��=�<F�z����E6�*�ƽ1���ygӎ3�6 �B]�ڲ������*4u)���B����H�viQ^F�B.+S��e�I��o֙[ʼ!u������U�އި��{��͊���� �ѽY�����(k�U��J?�Z�`�zBVg8����&!��ƫ�U����?^�9Z�2N�2�&���3F�O6��$(��O�-��F�F�;?F@�>�g��>8b��,�������#¤��bݚr����U��>��T�XY:�_G���/?�&(sEe���(3��J����p�	զ�k6M��ӽ"
�<�BLZ�c�'o������1�1s���]��ܩ5���4�V��i��gn0Ѫ�<3�~E""5�wk�����f�Z�{�L�}����Q��T7��8(
l���/����[��G���!q�����3m��/V
�W��d�m-�5�R7��������<Hd�6r�չ�.tA���O�2��r���Pईf�������G/��.Ո�2����J�=Rx��D8g��`)�ՏV�R��3.��\0�m��ܗ/}��Oe��\S������M���F�aTN��\��S�)��9�E����B>�]*<0�O>M��Ct�F�vլ�{��Y����6�&L'+cegU��̬����.Ep$�6`N��}��]aԓ��yǛ���w�;��<����X\<m�Q�o��{�q�:���_@}z���I�0D[��\�E>���#X���{/��|��8����>�'P���G���|�5Y�����7�$
�0([b	�y������3�=专��b���LZ��0�f,�`���N�
���3X�v��ݏk��O�}��d�zY�ģ�@�H=#7�*��E��Vކ������ }/��X�I�����4���D�������m͂��#y�?��_��+7t	�;_��R�rd	"�Ǯ���T���7�p����&��t6�!Ѻj�KdK�N��ȇf�x��&H^$2Pi�l'L|=:�>xq�[�,�Ǟ6ܻ��X�7HxDV�Xv���z��
p�0���n��@AB)�kr��}����G�����^��Fw�'���w���U^��z�:!1�1�F���U����-w0�^�9fH���ș�2�5�vqI(�nʴ� ��3�j$ʼ��8����(7Q:_�Fxt�#I�˱�7��~��3�}��f����7������SDo���o�i�b@�ps���^.r탵6
F�'�]������N�-2c�W9�ЁO�b���l�R�'���p�d5�؆�vơrE�Q����I?]� xh�y�=k<�lJQ���Cl��_]%��q��j�Y��dy����X�`.�mS��tL���U�m�������XW���)xQs��L(��{�?��Gm&�aȎ���L581���[� 74�������E�i�/.4�O�� ����Z��(ު%s��ԗmdx�&�ߨ�zN��"3������k+�rx6��h�cOXe�>� �1�d- �@���佗�%	Cw�,v���[(�����������b�I��mv�v�9�U:�@��㨾C����u��h���!��y��?�'�EM�������/Y��7�_6ā�;��\�ӏi�����E���.���S�}t�[���Mӻ�YJ8rW��dp|�E\Y@N"P��p ��V\[g�'�U��O꺴���-ϱ��L�0��ɣ�4X�&�v d��?wC�[ua��\G��]�������1�jw��  �;r61qP�[2j q�,^����,�������@RC67����!��?������p��yCwJ*#|;�ɟ�?\�\ϝ���#Z���&��(���*�p}R���]܍C�?�o��{j�;&��'�=���c`&f�h������($�ē�_��⮕��|e<�3!Vf\7C�ޭ�����j�����)����-�@��ԥ,�,N4��X�<���ks]��&`pV�f���HDf��A���8�t}���A�������)l�@�/�jH��uOObP�`a�'��eq�[s=�T�p�W���р��0�_�����0�ہg�U��A�.�\��,%J�<�&��j	��V�I��p4�`��ʸ欵��{�Q��7 Է�����ں�nҷ�C{�
)i�q��聯��NU�s��*����	>���&�& ].�y��=�r���Q���}������0!SN������PF�JZ5[s��	quƢ�����M�s5�K}��	$W�t���x�d哝�ThF@]�Y�K�e	��M凲No5л� H8��������P� �C�����Ch6��b���EE���&������m\�!l�w.��V*�W/�o���~��@�Nm]�#��%�,�B�˺�%4�8�C�5�lr�'C.}���D�1ty`�S����l���Ri�WY\y\	
��(���B�^a�&��O%vm���q�|k����iNU�K�o���|����I��F�?�(lx��-5��0�2  ������۵���='�&3I��5Tα�oЗ���)R�d�`S��Y�b������4 ��g�\���\�d0:u���uX��[��ݟ�=Y#���h�VbFQ$���U��<�u ���O�T���w;>���Y�ݡ�4�D���7�ߊÒ{Yn}P�-%�:9j`�fy����5W�-8X� �G��ޖ�81�G䟉�3�oPx7��r���E�FB׏������GN%�L���6 '�R$z@�u4�ܨ��6��.�U~�z�4���Oa��{���V@�� h�m�������|ᶭ@y��*��o_���NRwQi�r�g? �ѿ���w���gR�����rc���]ά��2[ŏ0�֔Y0���^AQ�����f*�&��H8ԲGf䊓 J���D}�f�AZ"��(��X�.`�z��r���x�9u�J4��ӽ��E�{hV���P��S��@S��)����rf���͠�����;�����ys�e��ϟ���.
�=뗶�S�-�ͺW��쫪�������5�K�<���~�5qM��p�ͳ�[I&��S�u�T��d�?)�����4�~�Qިc�H�Y���Ym١c~�Y�u3�%UF�Q'|�$S�pGn$0ܻux������Bz;lX�k}��#z�/�uq�WZ��m�F���� ���+*
��I_��Η�d�#��A��MN8�4�a��P�� �x��z�b������O'����z�#@�
����m斗����;&D]'l��x${�����O��3�a��pu�vΠ䊑C��P�<����G�N|XZ
5��'}��v�Z���O_ҍ;ͨz�/X�G��?=i!n�K]�p�#��6!;k��ƙ�|tl�^�Gt>�������l�R�~[<T�P��k�k����w�B'e6�B{�����W���Tk��k{�%ֺu�}
�A���
��߭1�����P�0  ��]����8�LO�(�Anj��UO�����xIM���B}�<{ɢ�g��#��7��h�����׿w���c^(􆔥G
z���9ツ��I�U1��7�����"_=�BŇ
��qt��Ǧͺb�E�����w��&�1*jë��"EB��η�AX�O^�:�.��7Qi_W��<DS�#T+]��e�k���2�p�*)t7X��W����iZ� (�u+��������5��_z�u'F�b!@1.VD�
]�մ�,�D,��;[�aMMꗤZ��ʐx��1��fLF����Gn����CA3a.zz�Kj�JJ��Q����
 �8���ʃ�̾��9�*�ǢFP�1����!6�-�J���{��O�C�:��1��y��K�q���=��.C7��n3KTp��B�(����.��8N���U�Ev���$As.�k�XG�4G��e6��:(6\4M=�����|�b	�?�&aSK<�S������6#��Z�`x�K\��2}�؄g����L�qn�Rla�a��T���;����g�V}C*�s������Sy�lǲk�3p��	?�S�a3��x&��5�cx��5(4�/)���?+PgV)��)MJZ)�q�H���S}5��)Sn�N�]]M3+���<�]�(x���F�Ϥ 1�!�䛗�SD@% :�d6O�xt�N	��Y�v���#5��<��_ސ�p����.�c&Nm3�9��$�
��oPW���6x2,���	|��E��N�\�y`9C8�̱`k+��rv={��Z&ç"���8�,N�/�9�:�/V@?�N��sœ�u�s*yd�κ7��z�ǲRH�1���F�-���;r	#�v��C��D�Kͦ�qԞ��+5x�2���v���;3.�:[(��v��O�2��ݼ�Nb|��v�t�><��dT��#Dº	SGx��,�n}�����´C.N6�Q/��,�=}�ǩ76������Mp�5�Y�Bg�R,�S��%���Bb�����E�θ���\z���ܩ�7���
)�DG��'9}a��`H�� a�4 6'�g�\�I꫄O6H+��~����N�� ��Ca���� �^fn�{r�7��uCu�|`���5󣒱*���2@�h>�D��u�׋�h���Y��T4�T>���h��p��)��?Z@%����܀��t�VS���\Xy��,�X
��q>=7�Zi��ɏ�g���Dy�|�����t�O:�n]tOH[ӏ$k��ޓv�p0s��>��a)��]#�q)}*��J�����y�?��)	Yq#gJ&k��}�����	Mqݗ��~�ޝ�@���ن���ΦP��p,Ϋ��d����ƶBR���%����y:iC��<�O���g!6�� q��	�k</ʈ*s7qD�Ls�J}����s�Q�r'�>�@IX�ݏc�jzb#{�Q"U}���0A�t�4���=��2@���f=��=��[��#�-IS�v����qK�����$��I�M�A�7Q�L |2B��1�
 ̙$g-RF�&lP$���ԭ�[�M_u-����/G*{�u���z�zr�+]v�>R�+�Q�q������0��ro(_��L]΄�+��40
I8�zG �|�i~���/����J�{"_I�/�s�:��Յ��N�0ƶ�w��Uk!+@�#�B�Ԧڟ��a�=I�i�̨>��F�_7�xZ���ȒR�!#��6���B.�u��a�!�)l��g@�����&,=u1�����������ȡ��#��{U��[��aW��m�*+�2��WE~�A�u��@rIʃZ=���(���'�̑�̒��Ǆ��^�E��G�s�xΆ�c��;ѬPs\e B�my���_��i�Ԩ��+v��;�)��H�^:�ʫiZ߯�Z!�-)V�;mb�`?g��Y~�����fQ��$o�)��8�V���O	TK��#��d-U��W/$}���b�3{��Hb��?�����	�K��lg��4��ޖ�@��_�RCja=�~�i�[jѫL碒+�:� �+�z���E_۠W/�]�Xf��E���Z�͡�N�w.'��ڗm��aԥf�q#� ��вG����r����#���t�B��ȆZ����_ۖf�de�d��IZ�
1�Q�e.�� �-T������ln]�A�*�Vm�,M/�?|b��g�jlM@:-�`U���j�>�	�<�̚��pt�8։�2���ƽd��_,7�
�%�vE�<7U�����D��S~F�̆��.���z�!g�T�N��?�ӈ�|X��NG%�l�_������t��!yf��J��J�����|�E�<�Xx�Vʦ��ٛ^��֩��L�0L�wݦ�	}�!9}Q,aR��`�E��ԃub��h�;����.r
k&�N�ě����$e�G�A|5y�#I7㬨�N9`�=��,T^O
���-̬2, �)k��+;MR�;�����%'ٳX#�U�@k r��vK��������2�X�}��Q�Zhh���5ϳ�G�u�GM�B0���
;t	Hs��F��y:����q�H$�O��m�������
X:���Ԋ2��T#
tNi!�t�=m�^�r�����=4�W��o�&;��t�<b�_�<��׈hzd�m��sb���܀*��U���0����V�<j�1�e&���D�F0�ǧF�����4z��E.�m��ģ�D��wז�B2*��>E��=H*����m�<��ٶ�|����_0j=v��|a��Q��쵯���A?5xk�w��UV��m9��ZZo�>(��_6^�v��8ϊ�s�to��}@��6�@��++����g،���G{'j�{��]q��$��i&��[�K%�0I�h��O���%���ܽcӇ�-OLUIK�2M~�����D|	;�Y���D��?�����we�	�6�>�q����/ 2�y�f�=>]+���b���.��\���X�!wм�V[Y������LS��{�ɀ)����­ºaj1ϣB��Q~�������(
v~��ZTց�}2��ג�MO#�]�'[���:Jx6մBu����f%!�2��1��2��i����W���HTr)��l��X�b�h@'���7�ُ�����H}̋�6�8�F�$��!��}����fE�C�!�@��5���+]����᚟�g&�Š����%��Mpi����O�%S!�SH)׋�R��T����0t�<\=�A�����{La���g�F�dE
�D�ѳ�H��G&!�,_�L+�e��!��ş��:K	��Q��6|'�����k�T�&�/]�M������h�8���Y7�\q�`J�G�[BzA�x��+㏿?�����h,��9�RG��Z��������#��wSu��+l��w}�5�_��D�� �=��Sȡ�6��S~���P��A����5����na�X��
�ꮺ��� V�k�J�Vg�X�=���ѶϦ��̌W����9:��7�R���`*K�2�=	ϥ�Qm��lو���J>�H�)w8�#��m������ޫ��>�����Fg��9�a�D�u��kאRI�xX�ԈG͕�I�qk�h�U�n)�L���*��#�Fq��4D[�yaLT��J���|�@E83�g:Q'��{�>�H��;n�JIa�����׻r��TK��ѿ�E�8'�L
:μ�^�3���WC0<�Z�R�����/�l��!1`�o����\y�/f\6�ژt��f˽��>�)eM)iBleh~P��K����sS����K:�g8y�?�p����x��?Ϯnp����fn1w�)��U�}��c���3�E�Ԃ�qi�5X�b'b2�����?^ |4Ȁ�fe�1���
�;Zz���DVi����9�1LMW5��H���O��8>��*E:�������\Al��Z�%Q�P� ������ 醁��a����1$�n �����#ۦ��������BM�����w� ���
��k��KuQ�lJ*�����!{�?�\��y@@�t!�N19K�r��ʫ�ֺ��r�\�F�Ӏd�[��׆We�0Mp
�u�;o�8�d!X�ӿO������'��lN�f��k��`����R�4�.�GRs!@�ڀQ���_��|��n��_�E?�1ͤ���bP�e-�~����,^���P����0�{�O��*�yĖ��]YJ���GU�џ�ց��򏄔�Q�2�_[���C�tk�w�Ej�����`2��'�[g�����k�� �Y04H�S�5�n_�>�pUw#������,�SD�����l���G�B�Y'�I��C�9��!	ef'4���T9��)Th?AL[ܭ޳o��h��t8�	%�A%[�w٪Hs�"�+}׿��9�<ٰ���D��{��BU�~����u�`�4<��#�U��U��?.�8��Gg���%>��v�e��
�0���_�2��w$VA�"���|)_��Yq��-@����F��"��ʥ]��?��s*	�����6S~˛gP#��2V���{W���s�L�y�C�W�پK=���>Ck�m�v]/�u>P��<F�3�F�b��s2�E)�9���<& �O�e���V6!x8'U0���ID��t�d�����������O"�h	��~'m�/����k���> C���WB�������x��d'���Ѷ�=�9�Ɲ|�=�9}���28-���̇���PN���O\l�0bc2�iS��ќL�,si��;ɀ��5�	��e���/���=�,1�-�̈��.�b��w<�O/������y��ƒ�������V�1�v�]�l�	�-����9�d��Mn��u8P�\�����^X<֢�uF��U�<��z�+�M(1A2����}�\vՙ�r�p�k�E��s�,"�i��jE�Y����X3�YV�����r U�Je���2	��m������X�d!���h�'gn�s7H�N���x�j�-xX/��V6�c���=�Yąe���E��l�8�w���K�F��I�1�В`��ͦ�)��dB�]���P��ܨe̡�=e�6�D�^+ɝ��:D��톾C��>m��,�����Cp|(Ui��!�>��H�"rD^�
�VeL�u�(��H<ͽF�46��v��TYt�n�u�5�k5>r3�r!�9�P����"���|I�RI�V��UԄM�wOf�Z݉�5)k�o������}B��%:6QQ����Ou�e�g��d>�ˍ D��=5�%�n�W����:<dd�Ƥ��U�gp���~���I�1q[!��l��ja=fLb��LWz�x��BmN�=wB�o�����va��Ч]KP���P+����VOJtB	�m�&��ĥh�s����a���q��sr���A��\�ݘ5a.���	4�(F �ߐM�����ZE��T#v�"$��)�-W��7�%�ַu��u���܋��q\-ENq�fP�R�R�¢�cDjt�rWK�Qޏ�}ǁ�^x��퍑i�rK�x�VV
J�����%M������-�;��TV����%�y_Y ��Z�v�$��%���)nP,�8:�¾���(�?r<�o[�j9�v�j^��
����E�L��d6�9���&���p��kt��� ��/�������������a�"�}o �x\�|���*����~��l4m�������9< �j1�08��yO@D`��z�Q��k\3\�Φ:�y�/��x���]�P��W�� #��(�����Y�\h�=F����:�04	&r����x��������m#{QA����h|��W�/m��(0>�C޹���g+�PܹԞI����OU 4`�~k��P|�ؿ�R)Þ���/H�v.c�.�{;�h����I��]��=+IK�D�R�C��	� ��(�{#dM')(N��o�7�E%�l���f�(��3�[����dO����z�!Pl����b�o2h ��8^�P�%5��,i[�e�t���Y�V���s$y����C�(�joO)%��x�VV�â�	���� ���܇`�'�z��t-��͡y��=ڂ\�c��>���_�·�}QUj�-� ��SҼ�n��a^� �W�����>=�GӘW���Z-|��HpB�Ý'��d% 	�����.`��qY�ӥ~�B�ۧv�V/�}�HMme� �����q�NV�ux���4�z5TU!<�l���t�[^�E�;!���RjziK]�>Q���!Οr5���p���MX�;;)|dol:�|2r��'��M�%�^�Ѿ��^ΰ@0x��kD
�)x+��| �L�ϒ�"�G�6���~��p����+�@���zl���gh�at�!Z�&U��.�j{��.W�p�@�kB����H�	8�8[R_:1�Q�o�(��zizl�+��i����n�p�мT��U�>����Hq;|CZ��Ki�-���L��s�Q���w��L��Z�R��˝o����m���=����T��+M��҆��U�Ӛ�>x �}�H"�3d*���j�l���ɩ����F/X��B/���,�pf4�xe���[|e��g�Mx7�d�tl�X:EU(�+ @�=W�N�T����q�n]��5I��]���UлP���9� �F�z͌U��o{
�6����i�j�N��'��ꋕ�A��usӃ��(S���8�<�̒��
%[lu�&��1L�����b��,I� b��gQJ�FhI�-X$B9��'�"��O���o�N��F��m����[
}^5�b��`7�'�nQ�0>ӛ.������fM4��������̠ z߽���gڣ�*轡|�`@_�!�R�N�p��[ſ>lB^��������� /�Lh�;���4��k.F;�A��GwP������M;~.��u�J���B�L��8�v�?nG�2��W��JpZꟁ��d��a���_�
$r��v̆���cQ�g��=$c ��C�
Vܢ�(�9�-��a���a��Y�D�G�yp������D�Hp(h� UG�D�B�|ދ���2R��!��`8T.���xNY��4��{\��}���cl�~�̀3�=U�����*V�h�.�M�y������F����Y7R�K����l�n���ڶ�0X��$�]xFdK�}CC��k� �����@\�b��L!��ݱ���r�ߏ �	M�f��r|x�BI��}/WQ)	�l	_� l5 )Ldi���Qw�Y�-�ݸ��Ճ6���J��L��k^�p�5D���x;���V��
	�=^�~8?@I�W��+�ï:�/W�Y�gY�/�v����ƱO~g���v�~+��������Z z�,��5l��?lok�L�8��.��A:��"��;-��o
�@1Q��0�B�Z5 1�ϭ��V��z��8��ϰ把�Qʽ�@�p��3��NK�`���p��δt��S�&
_�r�p%��c�_ b�l^:�!��SI�1yV����u�ʞ�WU������=}p=�p��C.�_\����r8�^�ʒ�t�
5R֭���}7�H3�Jh��@�R�̜��2�����$�Z�v5h�(�8�?A	`��a�`����P~V����k�o��`�XM3t��c�/���6A�s��.��)�a�v�.��1A{�!�Ԙ��v�W��~����e���0զW�ġ�;�}�O��)qz-,�* u��&n�u�{dȒ8jxI��LM�^�>t�ڇ�|c��;�=|�}�0�|-%bY��a�>�B�^l?�:��� R�f�&�} ��;��R1��hB��;LK���X�NQ�)��L'<��M�}��������]cs���ֺ@�|�$b~�`q�}��wL�Y["9�ϓ��vZPq��>��b&�3���xK�i��;�:�}��/��P����6|W(�h��IEޣ[G���m�2�9=H����Ȩ���pY��?��Ln�ztE�7��75�z�DW�C���ofc��h��t�r)����~?��0qF��x�k"��Cz���e�"�H��#�f�o�:K
���o.9�.��i�죡�p��EP�Ϭ��R�X�C-���7� �)�P�X�o�M��Bbq�eDh o�/­�j�o�*��HVԄÞەLp�ټ���m�\��a�Tx���;[��?�;K�Ƿ�zp%+��q"&<�7$� �bvn&u��`M�����[�]J="$�$sՃ)݊[��p~ɹ��ae>����a_��&�f6,ğö�u��D#�4��|��?��"�
�3�iu�����:ˮ}����&;F�5���Hw�Oh �輕؂Ʃ�l�[;�X}��,r����s<:tzpO�3�	��]`�.\Þpi���}	ܔQPJ"�I����A��9s�Q�����nU>�?�p>�YŖT�һ��Pd��rw��u����%���LN<c<U�9M��v}P[ 'o�]��蕔G<|�+�|�ڥ������23:8������>c���m�U X�y@����MZK��>�dmJIvi�db�W�PsA�T4þIY��V��Z�`�����R'����4��'���r�&�.
̡�6u�_�`MȞg-�)�Y�>������R5'0�`eɄ�GPBTM���M�Y�;�meJ�' H�[-�JDV&�����J�L^�~csLwk^]_t��35�G��c.uc[*�j��pK�`C5���5�*�Jy�ig(�q��REc�٬]�K�n��4��ˑ -�%4Jl����>�[���Id���S���`��ଈ�Q��o����S�+3S��:�}	���_�of�ek�	ָD�t�#$O�q��jWg'�� �E��&�k�BzTN�s�����@�[��zJ��_Ρ��� �e����⳻��W}�78O�D܍��`�߄��[ek�Rby�.g��"X�� [U-aO�+���BV2$@^Ӆ��*p��!R{��'W6)Ji 6c�^�^�Nد��c8a\0(tW]+P���3�i���2M�kEU\>L��&��R��K
�I���c+*J�����.���GV�x�L>�����%�RyOSbAE��Z��W��!�^3o�rL�I���"���L���>1��y|h��p�k|V/�U� �NJś���}>��s��:��M�f�f�;��<�ʧ��5m�������;��;$G��<0e&�0`��/o~>���� �x<5�ёz��վG�6�����r�U��]��z�7Kr��x�>\P�|�[(��~���[�����``o/+�hN���t���%Ud4�L:K,p159��d��<F�|7b�w���v���s���������{���j(Wk4���� yp�� c����80-��� ݘ���W�o�n���3�9�i9C�z�@5�c▯P��R(�ӵ<�g?"Ӊq����e�w�%VNVi)�����9fKe���H8���C�G�>e���F��ZQ���x�-5ö�y��%BS�~�i�P��O׮�R�ݣ�Љ�=z�o��-����*�e��e�s��*�9��U�0��ԟL��7�{/�v]����r������{+Ä@���q�A��^WV��-lt�[Lc'�m
�L-`f��I�=���/�o�>;����C?CZ������SS�8E�
^,�����8�<]@&�m��M�l�a,�zct��+�L�L������j���MeVM��[���;�6��O�
~Z�'F}�/K�bm�Cn���ୟ��{A�2߫<��� f���&V����F ���H	���ָ�nz-� Lh)dм����^��O�y� m?!B֒˟{n~$tvs;�k�ꙝ8h[��ܕRI{"�X#�	H�:kX�֓���]Z��+ASO3��p�S���0�w(R����1?� 7ݿw�d��M��e�"j.���$�i� �*�\bU�Ÿ�2�藢22�N�uJ�v�z���r�t-Hn�/�I�vu_Ū��Ώ���C� ϳ��ΡϜ(nxa�P_�au�=��1����d\�ӈaoJ�Βc���=+��z���;���:��O�0d�)g�)]=���e��$[U�A>��m���Φq��=��l9+ ��({o��������|� p��~���}+����b%�󢬴�������/76��"0'^���oH}oa%�����5aq��:����ܪv����"0A�{�Z�r%���e�/y�>	���[������(�1YxՓ��]������3�lҊ�����d����AaLv�̾��
�D�5å,�y�?�0K'X�T^6s4�춢�:�5)���vi�A�G��j�8޿���0���9l0=��iAy֯�b�9�����y���Ƨĕ���p��v��}�r���������C6�<[������ks��c���D#��/\�wf��v�O�����a���W��a
¼�+�)�����;�/�-�eQᤲ��t�w�+*�(�}�z0"Z.n�GG�!վ�����z�4���wǁ����$�[�#hc�_rP��Z�R�I�>��k��5���N��T��ı���OYU�5u1x\�*��	��ߺ�
�E8��A��Oܰ�sE�D�[�͈�6Ə�4���j�EEؙ���E�v�/���C����G���=���&�ʧ�u�QeXv�����m7sf���,�Y�����b�É�>�N��_ A��8̘V��!�W�Y0���(�����zMl�b/��L+4Y�GW�"S�0E6�X����U���|�ju���E
~��Y�Z��
�Ǌed풬SA�� �%ܺ�>�7���bO���Yh{I�_le@!Ţ�˻�s�ܲ�OcC��g�C�Ǻr@\!<J���Ra���c�2��e콚�T3����o�Lx��]���T�a�CA�j*2>��[XaX`��J�]�g�*c�f3�++���VG#kW�7\��qC�?"�wȥG�^�}%WL����>z���6{I���hknw�	�������L�n�7IY��+��U�`�0y�7Oh�s�*7�L������o^]\��\ ;d�1���֞>$���Ty�X��:滕2Y�
T$���Be)X9�I,�q����W��_>�/��,���81�t~K�T���]ׂ!��aB��T  u���"9a�o��H.��g��B!��¬�72Ǳ��q�$�=�;�[O��W�0c�+�v��R�8eJ8k땙��%l��LR��V��ӧJ��tW��}"�~�S��O�5�KMou���� &�X�r`u%�֜2�(��eв�+��j��zM�	ǩ���<����woI,��$�6#�s�*�z�p���/<T�Jѿ��&����s��]�mV��`��4|3�2�E�/,]th(��o9F�8�ȕ�n�RG�" %����	g�DB�ɭr���9="ܬ�@N�o�����jcw����ҀT�c����4��Z���X�.��w��nI������@ �	��H&�ܘB�'}Y��)���Ѣ�XL�3i�W���{�e��O,e��s&��g9���ǵ��ɭ�����mD8��Й9��G��kto"LI}�	t�W��z��U6��s[a��{��>���8�m��@ݸv�󇐒���H����}���ni�i�����WuXH���}õK$%����%�t�J�Zվ�?�?���ڃ��zg�P��ؙ�=/z������}��yqxd�2��%�{�,X�q��Rm�L�2���힅�T�PLj�
�{��N���X�!�OԐ���w�7���׎¬`�?��v�'�J;�ɺ2�wuM��u����X�Ba*�-|��Epq��4���=˳in�:����9��<���f�{����z�M�S�b���k�2t
�L���SGݝ+`�["KOȉ�$P��Z��sfϖ4��0��c�ro>W$���8�� κ�8�V����R�Ǹ�oK>�$j��.X�j��i�q��'��v�M����On�i�7L���e=��1��y�S.���Oиx�)GQ�t���KƴB ~ŀ	˒ ��̖�k�L�l�i@L	{�Z�C�vt{��@����6�� )R�~��%f/E��=�-1O�+��ą+�Z��,�1������Qb��P:#<]��O ��S���s(I3Ox�e�R�U}2��s���=I�j�$r}~�גE̚~�5�/��c�OIx��nZ����n�X���:|�h��BDY?���J��fN>F��r�s�["�,�_B�Ʒ�eU�n��̾�1���>�Sн��)��}"�lk3�N�ǳ��%�y:"�p֙��|3&Pu�a��f?
`딋dJ��~� :BP7z��O���/|o�`�|��f�m�	T��
5,z���ĥ{zt��i�(;ƽ=&��V�7}�$�9��DtmV�Lf����N@�r���	x��I&��?��a��<1:��1>&]�q�O�uckx�+����)���j�fH�� �`�#ᔼ���[NT�x�b��E�h»���|��>Bɻ�W`Q � =b�onE�|��s&��+X�%+bY@�Ҽ�����+<��0s���=-�kF����("����`r�B�F�������߹�aXo�Doz���qh����}Y@�5����`H!P>���C�|\[�;�I�U21�Bc���'|����}��)u@�iLI���ʡ���L�S��z�A=:�;͡�%�$2θIً�:pY>�}��S^Ӫ��@�VKh�]�d��0a��z�lg[#3�ަ.��T���ׂ����|0�{���Ԭ(��;B`��t����%WUw��c�k �O���pӜ�6�x�#�>�dV�G����f&�ysrM'��9�|����׸�� ��-�s������'���8Tf��s�8c'z�I����z`ɋ{}"�3lM*�=��4�+l�X�k����'�[2|��R��R�4Dxe��j\'�����q����-���X��	�㩙��5�׎S�AΉ	���^��Z,�5�3�*���,��
y8��5�VC䜴:�g��߳p֐���ۉ��P����H�5*�ᥝ�72�����E��Xy�3z�+�̶��KO���E{��6��=�r'S��U"ݩ��W��"�����z�g+_���j�~����JVz���vU��+�3����|�\JË�?��V��$ ���yٜC1u���Tf0C��ҮCL|&�D����친y�F\�$���0�Èz�,MŔM����*��N#s!ƻ'���DLI�d�:c�1	[�๔�(3�>9{in��~�����m`�5�q�1A�z胝4*���in$l@���g&���QWx�o�3~m@�n��`c�Kx�6��j{�O�4L�����]dE�=�R�QOs=�%�av�x<�@�m�(�9Vz(� ��ݢ�F��Q��.�H��π����%av�߁����ga:����ƃcAt�R���cm<�4W��%��V�^�@W9S2I:���1�a���3@��k�뀶��+�~�G ��l.�Js���TgN��ay+�C��`� ���a�l��:��:�h����$P�0�_��1Fu}b� Y�GF���x�����i?�a��(GJ�g�~��qSwu���MR�zr���%��������F�����8�9�.����9�ܥ���J�A��:�H] *:4���֔h���V�R^�Ud^���L�3���P髖m�ص�_R7
�q���@%����p�+�7.(��&�8�y����R�J�����YOP�{im8�l�`+���`��~�#��S�t��0��q�������yѨUޣ���[٤5cL`VX_BC$s�0 y�Մ�s`���;j��\��XG�w�'�E>�]