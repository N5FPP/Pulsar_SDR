��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��e�ik3�������w$����g|��J^]ؽ�2h ^A ���b�Io�C3���;]=+A��$�w7\�5ap����~�{}k�|0�.-a=�=d[?��;�SN9[�8޹�h���7�un�đ�ה�5.�=�*�g_Q�p�`v�� ���o��pm��<غ��J'+�ձ��ǚ+�����Q�[��^��Eӽ���~Â	�*  5���9ig�P�_�c�@̑�M�2p!2�-�n���o����ss�k�"\>��ǲ���1�[A;�5��wU����h��p���8�$ְ��To���C^�+R�c[eثݕջ��d)�S��h�n_e���5�h�݁~_Z�Ij-�ox�=��L*}!?��U����$�ح��˹T�m@�k;Fᒦ�������܀F^J[�h۷S��!����BWW& ��OorYz*����"k�&�}�	��o��/�h@�퍾��
>&�ŪA?Y��(e���)�P���������h}FwY���2R�\ʎ?$�����Q,�%m�1�n�z�q�K!���ׄ=����@����v'W/��en��'  j�[�F�� ��K�V'.���A���I��G��x|�c�e�ҐǍ7B�q���<��}�K�B�̣rr�&�Q��0��9G���J,������������P���0A4�(��K1*�A�ҽ��hw�$$�m=@ʊcJ0aq��d)m 3�_��HE\�K���t�;d�'���"�=� �y�d
��t�Ci;-���H��$�'�����3?���� ���ǂh#0�A�I��]�O����4q2��y>�ܨIn)8z8����������W�BᏳD�G(b�O��M��������%:��-i�X&N	?s����S�|�"e�0t��x�E3^v�<���U��A�!nh������w���h_ݫx���it9a�:-�Uf�����}�0՗G���M�<.�/��Cn�A�$^>!�*o�6p3��
 ��a�b�s�f�O���ip2kx�:��5��PT�ܞu��G���1.�S6��5a>��"��8���e3��kF�qx9+K
_���z>gh��^!�&��D��ɛP��˥3�Y:K�v��2žCD�9nHiw��?诋F�@c�f(�C�N��s�?���ʿ��x
���@6���������F��~w��:ٕ0�^ǆ�s�m^ڨ�"`aIW(M��r�������<㓩x���*0�C�0���Ӵ_=gb+�2�Kn��}�+I�3�m:�N��1���o��YԦ�Y��=�����(����}�����R��k?�6����RX��݌�P���3wv�њ���"�t�؋\̝����U���pr�����:�/��U��&�;�E.ٶl�S�񇰬}����`)|];�`��1��K���9�Z�GO׮4���6��"qx� �}kԪ�����d���Ȯq;�U[kW�g��m�������ĿB�n���k]�q�����$�����hC��I�v�-�u�Ԓ��� ,�Q���jr��	$7! ���*��f�$���;�N�-�h��]u��E1/�j}�v�,p0� �88�\���9~��#I��!��k/�n�֤�����2��5* ��{[4h����
�rMj��~��/!�Qv�]�J^�;9��;������:
�����ˎ��r��c�s���c�� 4?��.�0R����~��J��](h@�ɒ(���ۨ��AQ?�Ok�f^�#��Uf���[���E�N�%���~���vW�tmIk�r]���d4�ȵQ
\�$�K?�ctv��9#�M=�٥L}�i(�d��(�c����d^]������ݨ1�F� L�5����%��
��gCqY�In��T	ĘA��L�����t�f%a .���R#�3UvirK�v�d�I�4��1\�n/��~���p���RW[@�7<`�Au�z��;@$�/�j���v��h�rUm��P$Ed�c ����9�����#�2�Umte��؛GĜ�orCpF��6��n<x6ʮ�T}���aD�q�5=#2����Q�ddp$�x"�3]�- �Bg��6%��#,_Y�儔X����m������#���}m؎��f�
�����sYOa�(��k!~���	]vz�[h��j3�Fx�/#����4��ԥ�t����"��`���� �G������,�r��ǹ6b
G�u����{m�qt�4-���J������|t�-@�~k���X���i��{�#�0{ƃ��1�`���U@���r|I�șb��]����?N��M�a������;pc}t��l[����N�dB%����&Ơ�g��g��>S��DV�Ƥi>�yժ��yyK�2tE���o�h�N��L`kN���B(=�%ܝ7��������M�d���}�*��O�%i�qa�;�4j�@q�T9wA�v#A��2<���@�����{_�6f�A�4�r�-�$�:���" ��������U�K������������є�MX����:<@C��#]O����`7�L�">Q��$����F��-3�O'%�Ď`NBPЂ5��8�[�o��/$�Z���N��u~I����&H�K��%��h\�ӞS>}�����H[��N"]��WqQ�u�z9U̯x.ȌT�v�s��%���z���%�x����_�Ev/P����BPY����a��
F%��Y��|�v�F#^�f���sk�Lw@6����Z�}���t�pG)I�{e</*���r����2
'��q;�)i�lq?��Llc���>g),͎L��fG�Խ�� 8;����:5�2�����Y��B�A�.�'c(W�n�/��.o
�G���S)��+�Y�j����Uc���>�s�Ci�X��j{�
��С��ݩTv���2~K�4�0�,��A%Vi�ϊ�\L�cC��5���P8;���u��VrBJ r!q*Q�ҁ�c��B�,O�(QQr�>
�$��?��)f�l��١����!6E* �1��Ke":)�� �|�j��)�-z�{��4d��Q6'�"٨�:�8��2`�;M编7�=sfG:W"]9�;�1�!�So6,�ܷ	�y�QRn�Ttk5��j� G>�ti���{�!ȧb`�ᚎ�A�ѓ^�#�	�e'��i,�^�8�O��.���sԈ�"�hZ����4�nm��(Q��KL7/YV�t.t����Ӧ6�^#��S�'�����apVD��L�J�7��=��=볩��P�F�Ti{�Y�G��2�J�W��$W(�5q����Hxt���pV����S��׭<04�r���ӊA\z��f&Ts��C��^��1;�J�.e��w�1�	Z��9�����(�Y�Q �1�1��B����B"[�D�K�M�b��(�z�����p�rm$��ɦ@C���5(�~z��xf�3���ศA|3�}A|U��>��2�²'7�i��U�����hg����z���יͬ�����w3r|?b��ګ��z�<�;'�����>;7��@&rn���\;=L�#:.lW�n��g�32{�;z�>I/�z-E:��8~�0&������5�(��6���9�偨�0'9Sl���4�JJ:�l�a4xxX��Mxo�Ӄ���/|��t��E�1u])D����؂3�cw��+�;8��?m5_�f�E�Y�� L��r�*�9��K|��?�8*��RYa���\��$��y�6
�3q }>e�`��J��#m�H�=^qe�����% �^�74�K�Y�r9n,-i/���`=���?N�
�o����cW�A���N���R6�Y�&������!5 h��*؁���q��A�vt��W�t=��  ���t�vٳfO������-�\;B��h�T��*��]�i����ɦ����X��B�O�U�궝FZg9�������~-U�_��WМtz�̹�y��D���&�_���Y�z����*���Հ�ג"�*�R��~3���;(��?g�J3��'�[� ۴wJ�4�]�V��۲��I�����Ĳ��A ��IA �A���(�"�Zu��`�8>2���[��.;�֭�H�v�\w4DR�x��^C�6�>�iV���,�$��A=8f�G.�8������Üo��J��Z����ˇ����pmYq�{�W[x�a�,C��xc�ă���E����wC���d���]B���9M��C������ºǜH_\aXc�V���A%'�u-��{��-U�J�S��C����|�&dI��њ'����(��a)�id��~��*�c� �4#�̋5PUM�T�$?z��X&|4Vd C��ԕ�;ӽ6ײ ʷ&ҕw;�O��'4-I��8��ɋh�������A�۝ْĀ��b�_���м|!&61w�Q���o-����`1�F&!��.�3a�
7g;�~e7B��sϐ��e���PL|�h�e�]9�dN��h�fL��(dv��]�U5VH��qF���jK�ļB*b���9_�k����{ײp��Me�^��ه&�����Wq��	���ތ�$��V;)���������e�syb��xm?8� Y\CW��^L�=�~���v��\�y��"��S�|F��.����8�m�zI�W�
��U��Y��T�X�ru�S�ت�&k���<`5*>��/��p�p���H7����C%Ƞ��u�iq��z��s׏x�`�t6\ONHH��},&j��=[ӯ~��l�혻E���}Z���g.!�=�ƾ}4q�%�Sk�4�4/�<0-�W�Y�S9��!�\Z>�"8�̴M���LI�q�?
�����c�z��v�Q\�a�*�y�9-�ZA�e�#ϊ)-�_��4���a)P�&aͼSY�C��-���t�;]���FG��������u�?�yߎGN.D��&;�Ƕ�,�P���U9Cb�Q�3yU1�ο�y�t��G��'짞�Hg�3�ll���~��9�l.���.]�+WִŹII2�o��m�^�sV�|3P������H�����T{w"Ƒ�)%�!�lYeq��j�J������C�9t�F���䍃�KіO�d��jt"��$��R�/���xaF�$��m�Ą���>R{!os�41���^�O���I�Q�*�q�:59t麃XC�.��W|c�"J]j 0����Z��G&0���?5��	�e�g]�tY�����g��S�åư���P'��.ώw��4�Ҍ��*Oltr+��0�;F�<���`ݴ)��!�("���������ծ���٣�^>���x�	��>h����ݙK�����q�$���JY��\��#��G��G��#�"}����Ps������s��%F��'�K55���?���?��-A�V�U1�4U�������[�?�2|�T��t�+؛?]���\�є�� f��,hk��RM�R'�l+�>��1Z�g�r{f�0pʇ~�z�����VBk>�4lC��o��x?p
�oP��"
�B��aN`�ޑ���i�r3��p��j���h�� WRρ�����,�`�X���n)��؀,!,szEg��ڷ�k�_���L�
,�bzs�+���u8K��bJүQ՚��6��	���$R®��|%u� ����E ��d螭dG��O��&1��Jv���oU��&���K�R&�Y�W��e|�+�!��7����yo8x�3��Bc�7���٭��	kY^���_�VyQ ��#�'[����F`�F~��V�B�ea��0Y�쁪�9:4e)aޣ/_-����*���'y�iVP�3�WngfQ\6E�������
�,�r��B~���H��@�͌�m>�g�s:�Ix�+PQl*��iD�<NMG�^_�B���@(���
�@5W�ͭ;|��o� ˡ��<�k�%U!tT�~��
!����zq=X�Y�zϡF�Y�W�]Ø;�I�Z�*����,�Τ�B	�X���;�,3����J�G��������!m��h4��lM�J��
�E�Ͷ�MSy,7$�W�q�hѕY�J�%��(j���2��.�B�h!!�Z|ð���y�=R2鶿��M��e����#?�_M��K#(�_ł?MI@��ś�`?w���@2����^�
���L����$S�Ӵ1�aX����w���nD�y�5���+L�Kx���iP���W�S [�Z%�w�&���=��!�g�IdF�5;?�N�ߘT�c���o��fE��O0�f�+('���a4I1
r�3���?~uԃ�+q�Z��z��7%���!c*8냡��\XV��
���W������Y�R	^��Ĕ��~ě�x�So!F)��.��eo�Mqx��B�"�ǖ-��k���Pq5�`�F<�\���_�F0��I����9�i�OS���	�Zx�S!R./G	�]�����K��4_`��<�)�m�-D�o�y�@m-�0H�+�.!�]����<~�[j��*ѳ�`�kwt(��\/;�K���C���&���J�UG:$
ZF��?Uh�C<!|o���4�T}�C�;Dq��9�����;`F�'�h��zA���4
<��F�
��!Kٻ��So��P;�lQ)��}JWF��KX�$����T�{��lҳ�����Š׫Y��z}�5���T�����K��&��3V��e����?V�|���<���&K�W��v�i|�M:���̈́гt�JR�%�I�E*�*P��Iˈ��鹿�1(U��~�{��������cׂ��g��^뗘s;���̧��j���+n ��<}r'�sJ�4��v��.'n�x���,�y��1���Z|�k=����L�Z��:��t<!�.�W��W�!̛���?���u�8��5����1�Z��M5Т
�C��E�ng4�w�T@@lxM
�,%��6�bFF�,�߽_Yr�k-܅���n�[��`�O!q�U����k=��kZ� {C[�BUgnЙ�G�-o��3��)d�ₑ��f�����3�F�J��ጫ�F��~�]a�5��� 4bR�B����f/�������2ʣ�J�r4�	B֝����2q t9�z�E δ*���R~�5�k���G
�X́��U�U��b���=��	p$GXT�i�f<-H.�.�!���F�x�ԧ�7չ}�d�OI&�<�#�Ce�	���_�+Ɗ�[�g��(�p�R�e�?�x�=����BkFs,\��"*Pޥt�La���-����3@�S��cOjA�����
{O�t�!�=��|U�od�s�	��gٸ���H]����~{�O��5��䩀�$R�QsѶP�<��׵��6��;��x<��,�x˝�T��ɨw:���7�2oX���f��0�Lv�7��pU��1k����>+�V�;�@�|A���]κ?Oi��L���A�~�9q��ƎL����`�	<>+&;rm�A�BS��>�c�O�=�9�y|�w#�*G�\X�L̬b�R�����Z�=_Ù��a��J��1����і��V���4����6���أ������)9��xۇ�D��ub�wū���u]4�4����-�F���W��F"�"�2���Gl˥���3NF�K��s�.�G��<�m��b �Qo6=E��_;���C/�Us�c�,�W�j)��ɭ��&��*Ô[��P�l���?��!�TvLo��%$��+���eY2�U�.j�z�XA:ĭ�mp�����t��M�F�{��Q�)Z��O!|��+*O�y%-/6�����B;�R����-��w�!��� �y��R�����v-7��_$i��M���2��^��>��k���Ԃ���]Q[ĤR@F��j>�f��3Z�y6�����Ⱦ�u%�uM�	xr'HJ�u�`6��~I�[�E~�f�1����/�|�}Wq�G�Dݸ�(�G� XW���Z�`,uoBe~'�5��f�	+7��3P�H�����َ��t���&��$�;K�h?>{��E�##A�*�ħ677ڬ�L�"^�OH\:��%M`��4rԥ�u_m�"�1s`!~\��%��g��$�%=e@�t���l#�rS�����jY�=�c<}F�vqP���q��bK���&E	�d���"�Nw��p4B��*��
(���慗+�NU;�G7���3b^�)�L�K������� �b���>���N�Z�=���������0v>*�W���:������UV���7R�.%�8D�}>hԺ\���A�m�O�(F���ᠦm�����O�63UŨy��~y2C�(8������Q�kky��>u�}9s���*)�b����;��Au�������z;(F,R��nS�4۟������8\���:	L�|*�ܵ?s�˕(��Ϩw1��o��QdPu����DϞ�tے�4O���7�ad��[��1��^��N&�#nY�w��i!5�W�G����=5p<�u����Z��qƙ�4!H�'+�<��� �ƿ�`T��U�t�Wx璂r�
����u��e%����p����⤿�1w���wDY�O