��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+4ڑxſƆe�Q��fHv+�+Pn_<�x��Ԉ��5H��k�ځ��*����ʻ?Q[vhŜ��yA�B����3P� ��"����
--(a���@�_�#�D�pz�
�n�ˋ��窣��W�Jn�=�|�"~=8U���&�#ƿ��Ҟ��=Mx
���>Q9�9�
�Z�-��yA\$;�c����v#<�X��v�l�O��%�I7Ϩ��<O��2��6ol�y�#�e3"���Q���L]�̯���v�L����z�<"kw��23(?�8Ԓ2�v��WV���x}\}��y��F��ř��<M_�+�w��Z$�ş"f�%�P�ΪhG���%	�)�ź�Q�1c�Ȫ�ށ}7@[Y].�@���T=�5�(3��u_^E<U���v2�2���Dn3���˃�4�3�2{��k�Ĵ��i�F!���N�?ʭg�8�r�UO�s��!I�@_��_LKI�}��m�����z�n�)��Hs��1e�p:���ps93�Yjdִ*!���O[�l�7Wf�F����@�����O�.�yģ�EP�W����|�Qw�����}�˵0�\�2"-��v:��q��0ϺV�"%���w���'�-r�SEkr>��lz7z|kV�P��#��9�)<�mM��ޥ]�����l{���m!��iܬv�v�� j
��疸�6�Z��HW��;ѯ־,��FN�n��d��Nb}]��J���vE"����1,�>|�\��xb��;7��=_�e�/�ї�����VXI�9#�Q�s��` ��Ԭ3ƶ/C
�R<�)R�ѣ�d �T��ry%����q�(푀���D��Ǆ#`&�#p�-���t�)���BW�4�G���v� �6��R\�I���𗠫6@�aL�����6#F����e��EocO��ר�$��-��ܧ$�}��@kI�>���>֙���Gul�}�ſ�?[�?����5�8��m�S�F��$vZ�j����݂����h��-$X(���[9;XȞ�<�.�>o�\+�Q�2o &��m�K���QQ������������{D����ƊVf0l/�lq�3q�8膆74`��e�c������bDF�.k�lS�MU��:�)c0�(%����A��* V�]���i2��G��f\�{�"ZF�n7����2�P� (b�9��z9��EZ�>F�����"�a� [��q	��o<=�	zLV�y��X5��3"��4s��������!W���,9
�M�B�U��z��m�=6L�;��
E��?�)�v�oo��aK��TIjx�9�_j+����}��^�̻i�#����{��Mk�p�}���O���������Vg;�>��?�0�K>���-��ٰ_\ؐ��������M�F�'�.���?���U���7�@��T���È�I%�8���4�
~S����#��"�݄T�'ur�҅+��Hs<�q;��P���x�|#�2Q���7S����a��
]�Wv5sf�4�[���	c�ʐ�������	���9�P����	Ʀk�K3�D��%e�>o�蒟fx�Q+̿�o��Ti_ft!8�5s�s���bI���㉻���S��9��K�<�9���D����uUmaO�'}��:+�:�%��֫X�=�+"��0�p�a��f'�U�G��܅C�B�I��'�X[x�}7�����I��?U���I}��4�8!�O4��R'����i�k�}�:>� '�p�U�(��y۾9��R�T����J/_�l�'է'�9��Q�[3<�(��hN{{Y��k�~��t�/ss������m2w<e3�%�r׵�0������r�/<�
,G�n�Xv����X
6ZrC��p\LB�(���CɆ�]���\�D�i
A���'dY���Q������DZ=o�t��c�j�Ж?j3:�`F*YPD�0^�0��k0�
Y<��p�P^�2����Xw�0QN֔�3�xV��257�i�g6&ʈ�̿BG�8���J����3rmaי�o*4:��WZ붊k�i��/�:�}��)̱������V�W#�w-����i n�g̘�w��-Ǫp�,:���`�V��R�5�4ǁdr�������͹x��޻1�JO&�<��[p(�y˙Im&0@C���	sۊ
�MH�n�%�/��Э ����gO:CV�&�#[��5vU4� ���� ]~�B�%`���Y��=���Y���c�So�jC?�lcbu�d��\-�Gto��oY��{��E��'{��j~��boLO������p>_0���ةP V��Cg�uu���=��~�=^WSt��-EUI���]N�����_� p��?��`�PU��]�8[�!�=6��҉���v.x���y�T�Έ��he��J���0C@{��QV=N�Wf�7OܠW�K��9bl���Ⱳ�5?��\�����uG��Mz!)��[7-�@69^�J�+�.3ɘ��B�g�/	5�?�#�v�k��Mʕz�L�A�c�(�,�펻��#]�4�.*���f&��u���M�ԥ�\�	?�G "wXp��Mb�wI=��{$�X�zT� ��m���ri���-~}�C�W?s;����x��-/�k���iX?u�;�M�����I9�y��E�b8S��L`���u�G�UD]Dz��+pǛ��W��uQ��Ǻ�v���Fx��?�(��/dE;h�9���aN��H�*h��1E����*t ��舁��ª3<��R�<!�