��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VYkM�#j>cR�	��~����-�A�l�����59�3�֘���߹DP��Z^�g�Ӝz�>�t��� l��0��ᖤ��R��v�q����ôW��%�A�4(�;M��b��N��)�����r񶛜{h,��8�z6s6v�п�^0lR})�V��+����*!32��!a'N�	���	98��$@�����{}��̨�S�G6p��(`>O5T��zI7
�����)2u,Qs�a	��$ %�7��H6;�mi�W�&��w����~G�r���!�;ԵcV����+�ļ�(p�~�&�0^]P��>N� ��q���]#��zj������V���H��g��SzQY|se̮���=Y&���ߊ lH�� 3�&���j��]�0'�ԝ.lui)�`F\�����{gn	eOҊ����͜��4mv#�\$n#�޺���R�OE��)����5�Q�,�v���qa,��x����Wmn(������,IJo#�~{����&X�o�u����Lf.�W��3t4�/x+�S�*ja�`e`�gB�&K�|�t���m�ˋ\���ڃ%��f�4
+�K����)G�hz��X�����@�Z�1~����(��T��r"gr���d��X	µ;�C�|b�[�]�N&׆ޖ6�X��M��Un����"+:����u��-�_�V�0�����9�mU{�P� �1��^��`��`��Xڶ�S���v�=�ޛ>��|_��:T�bJ �K����G�h��r7�윏=�}��Y=kצa(��C0�T0�5E��Jo����jE�����0����0F�����6[�U�3+M��r���(�1����E�]��#ڸ���{fO�l�yh~L�����KFg$����3"�������T۹�=#���d�}e��Oa$r�i��>Vf����d�r�*���=�b+
��T��U	N��_Z+x�����)9�J��ܭ� $Mq�x�a
�-�8kxm@�oc�G�K��A6M$��Co�.�Z����ykr����0�ڂ���V�8bE���'AM�o���+>�Ԉ��N2j�������R����+�5���\���Q���t�@PW��!a��.k�{Tcj�{��?#����[P���x_�J�Ka��|�
��e(Ë���v4�K'�Y�@ue��sq��8OG�e������� n�ښ�d�'�"C=��g�c��E5a�stdQ[O���`�����F�X5���9#^!t��|
���Z"{6m�(��n��bٻ8���K�N�u~�{pL��20��XkO�ߓqۊ�.�w�b�����W���e��<���]�%��RbA@#k����4r�����C6���K��(G�/]XPG#�,*��<��T����m ,�tK��23��T��5Ć��a�M#[��,1�Ձ2m��I��*�Y��Α�W�OH�������@�)hԂ��a2f����E��@�ҿ�3�@e̯��C=�%�Y'Iqi��X���(X^��@�1�կ.wm�����V�������.�N�;�ViB�6�>B���ìYH5��,Wa~��
h���r.vPg@�m|��9���,��x�J�Q��r�׵�H����X�S�z)��U1�3�X�&Q������ş�R�]U+ �''i� ou
�&C}�k��Щ�,�I>GO�a��#�]�(#�fa�.��y$���D_@�'�Ig��3B)�%�� �a6`ʖ�W	�J[A��oS�3�4�H�^0��N���ֻk�a9
����>���MQ���Dbqp��-*K+��$�O(yR��t�"O�*i�1��<�4Gi�u�B��艏�3m �/��� �K���2����H�:³��b0W�bӒ��/ ��[�+����ɴ�20�rN#Y������}���j1��3��M���ڬ����:[>$Z�Z+��2�Yyx�d�w��nZAP�_!sVm�r��� ^��Dr6�%
���\�k˱K�d�
3�fT��1Kw����a!��;��N����rD��&t}��Lm�������:V��a�����4����%�I]ȵ>�����$�\�2O�"���8��eĥ����T xiŨ2!,gsz:�u5���ٛ�!���8�wp���r�e.2"�&۷U��!S��q5d�8c󭟳�S)�H=�$X4�_R��g�VQd�&��l�V�Aq:�*�C(�E;������H�ZZ[�z�Zl�q�:3i���D��Ap�y����O-�a�dI�� �_z�|�8��Bh���X�9��M	��������1ͬ_`���Z��Ľ�o������ �"�X:�[{��64E٦����k
��b+��E��G�j�Z��/[`nx����jtҴ�姨:����<Pҝ�ݛ��Z��O���?CG�J 	FCTG����]pg��}�V�QL�H̆���:�G3^�;<ԔȠu��}"�8�Ro#c�g��,���df�4�Z�L�ZE��R���܌�p���(�NΰFW�~�¤���	����#-Uû��n��H�o[��|��V�h����[����q�!报���C����iY.�7\`(a�|�VJ��e'����f�O�ˤ_�ѣ?��u�O��`��O���l
n8�D3W�kD��t(�����F��kK���gN�c��d���Z5�
�� ��(_C�86E_�U�H$��GWA�gk��6gQ�����;Ugu�Ǡ���Ў�c��c�7�L��y���8P���Oɕc_��y�:��1�����o��2�Ea�d�T�23�Ԫ�c5���N�P�n�z�i۽�+6�L@ 2��b7D(xql��"
t�7��I�`c��V^��Dˁ!~my��?�����cf��X�������;��n�����RN�y��M�c-��~Zt�Y�T����������371Z�]���.��Mz�{a��F�깐u��z��&4ֲr���G��W�0��Q�i+<�j˔r�"[^\E��%���`	��>:�&�b��kv��TtӪ�L�aQ��L�y�(%�� ��zչ�/�y��㇚�Q&��"S��.�X��l,>ӽ;�b��f���U��� �Ui�c@��Pf�z�|���O�������ȕIFU_�bnX�{��SkJ�2"�o����)b'�0ь��Š������3�IvT��bq�p���� ҩ��ɏ�g��/}��"���7�����sR�Ӈ��?'��*�_3	�3�5��J�<W��x�������O$<�Y;	jF�j�#-1
�\*��7�h��w�z(-`Ӎc�tZz�ȹWƼ��~����vH Pяj�U뢷��Ǡ�։a[Ǝ�I*H���tIϴ��-�>kI�!���d�D��=Wi\�'�Գ�w�����������	!�e��I7_�̓.�����L��L�����P5s�[E	,i�U�4 �j�;�V%��E4D]��;2�8Z���y�?q"���s3�uA/��/�C��-�l�d����X�	��ttz��_}���n������$b��ߢ̕�?��=E�[ѾQ�׸�sYֽ�g�Ud��`�G*�-�Q�P&�'k6�bJ�o���Bת�`gy]&7+f6%Df����ґKA�дL�B���� ��}���C���mˍ��Z����,�=��K��V�^o�H^�%�m�)�	Ł�c�����'�'r��,K_>�gfM*�C�� �����0M���[�;��X���r<�>��\���5`UK�B�&[�T��A�c�A����ԁ���=,�)Ha?�枔�y|�
�~�x]�c��8lZf�{�ڔ*�yl�|&�Fhyb��aL�/Jd��t�*�#�? O�ag[*`-|��H��#��Tr�ϒ"�w��S�W�F��R
'K��Q ɤ�WE) �Hk� Ѐn�G�ϊ�ߤ�v�>��E���tty�I�)��%�ȍ� ���%��V܊u��ݻY	��ҽ��j���}�n�#��[�ϥ�����GS�p��D��ځ��6L�J,��f�����x���AN)��P��+���ǅZȃ�lW�b"��B=���n���B:^�j����qog����3�1����2Y���]�/�a��j{4%��V5e�/o��n?G�|�<h.G�r#���L&"͐��u��1\#�M&��Ϝ.� ��|�	-�����Y=Ȥ݈�3
�8�I���	�3bFèc2�7c�Su�.�.hzs�U�/� ��~v�l:l6z�%Au%����M��r�g�=�ƾҽt�KA,��䙁����8��z��f�*SԒf��&�]���
#Zh~1��}��|����!P�KC֓pJ�����I���v)3$�pt��e<�i�:��k������8������<Y���K�����x�=p|0�%�)C�y�L��y���4\���M篽�����
;f�jz
"���ꩬ��ޙ���4��GЈ�+�x8�J�.����~H8��p������j�����bV��?�	j�����N"I�w/�����&4�M<�����}�a�C��Kn�[�%A�
aJ��[НPwY<֠���/�;)�5s�OJ��=�H
����~ؙ�o;���H���:�������.���.�$�N�#��VVE�:��T'I�Z΢`��Tr��mQ�t|*� ���yB� Xujr���I��4����m	o�j��{A^O�Sj��J�� �BﵢOu��׾��L�J(/��2��D�4���ޒ��>	5�#��s|��!f��.Ȃ���������L׷��˙�>������ -��P`��2C��I%= }ލ��V� Sx�a��P(��4�e�d��ꡈ5�$9hw���T�$gP�%\�jƋܦ��w��@��:�SGf�6�"�1cZ7�f.W��|�xԕ������*M¢7�}mDRnf�i[�g�/���i����M�ƭ��b�:
�aP�Q�M�3����b��£�^4}��+@���C3�>�m9�d]�U�l�5�̼_�k���/*&!av���P
���?� g�TG9���b7k[x��_���deD�f|��uQ��$ß4��
�� E�e���������B,@RHzŬh^��(�p���(lJZ����GÛ�7{�2w�=;��[��|�dC����!!8����Կ�:�JT�����ςg��N؏D��]/u
����\��5��?տ��wh�s$�>�象�gf�"�n� �ؑ݋�TEJ8��?w�h��Jy��m���An���<4� �<�����l=�p+��,���R!�}F��e�R٣�I%![�_���%Acj�i^��aԦ:�o�T��$ �:9��L"Y��1�T��YU?x���f�'n��-tA�!3ƪ����+ �íc�
@,j�κ&W�b���Ԡb�x��˨��镁���QL��w��J��"�M|��`h˶v�A.T�؀�(���@�s L5-X�Jw�/��-�'u4N��T����g���ڧ;�|+2;s��y���a� ���o4��m�Hy�hw�dr�G`:�F�q�w�>��vب0킽<c�TΡ�k��;�w@���4�B�f�ޥ0ѥ���H���.�lJ5��Qk{�|fU_����>�ͬ���m�M��B��>�}2��=�c1�������]���4�C�w�. MJ$7!(�8�eX��I3!�ö	�T�N���ec�.��ˊ��?�-J�"U����]쀹ĂH��Na-�U��)vy���1�D*�B'��,��F�g�W�$T������(lvɐ�\z>����������{>�"ݔ[r�q��*�U�	,�T���$Nĺ�m��� ���������<��	9Du���b���Yu9�Vj�������^�Ʉ�>Qri\R�5(Z'�&	-��t�~Dc�#i�=�˂;t��xw�U�M��s~�Ԧt]��+��Po�n���_�v��Ёq��@
���6�e��7�܁��$�n��3|�%ӘD�[�~̓&�j�����:B�/�u' ^Ƙ�q���@�כDun-����=��!�zp�Y�����(��m)�����V(���Ĵ��N���#_��D?��?I-�c*�|�3ɲ3�2���M��tsKC������ed�}�촐vnt�H�1si;��ma�z����&��]�GB?MJ;C*(���[�8�G$�X`��Ng��n��G�^�yP�l�J���[մ��Q��5�f��|��pb9�J��ǋ��T.������N�Ѻ���KU(�U)�����$ܵ=e�%�8�n�X��G�&a�~�S���eU��g��0ʫZ�����y�ܡj�AXI�C����� 9�n�/m��4+E�]@��,҃��L���D%x#;���kRzd�0���=6sc,�FX�F�`)>��t�v���o0�5(�{�J5d8�H~L�zID�,�_�T�wo�|j-�x
{g��0T�F�'�����8���O�����1��
m�����6���oimy�
&(�\0�����8���Y�����(��'D�!�ksY��*�U����+�
�~�<���D�V+ۺ#��˟��{�B5������� � 鱿��í�9��u^!�Q��5�o�gBQ�3,��	*0��"CwU�3���OEN�hu\�&��*5�2�Ȭ�\��Z�Ax����Y�:��Ӻ�Z�9"�v�=����4MJ�a�MW����p�*$�������Y�U���7�&ľ��2���Ӻd��-�7b��]~��js~KnW,0����k[0i
i�RE�#��^��ȗ��BVc�(=GD����;VY�X�f� �~Wl���	�;�@n �L��$o�A�F��n��+{���H0�����pi�\T�ݧ�_Ў���o�e3�E-mep'�a�Ge�_��~�#�}�]���N���|<��3��?-�g�W�_��)M[]���·)�����NZ=�i��\7����±���:��%8�*}cvM��!q|�Pn1b3�8[H��Mb@N�GFjz��
cD款B�u�sM(,1��[�a��. +�Dñ�6��ԏqL�0���*�d�VΦ�1����) �Z�5�O,fzM"\~���]\-K����'r�*�z�-Tnz��Q�4��u���c	U���ƝW�=�Aeֺ���>d��9�3�)�˖�}�p�:���2A��W.J(�y,�c�K�ْ�ڤ��DPz���AH�;^{�F�\�R%��ELُ�19_FKwSf�<O�����uu�z�6!##y����p5�g4b5��S#������\)**�KyҸ�p����:�W�]��=X��9�zc�� ��S�ŴT.�2�r�����a>?堮!E��D��<@��f2̯��������?�o�w����d��Ņ=~ן��\���L"p�6}�s���SMz��L�n��i�C"]����_-��5���j��ڮk�����A�$r7���9�nA�`m��s��C�K� �,Ji�Tf�J_Lܡ�na�ٸm#�j[q�k�f�G�Xz.���_1a�לO��lv	6���J���d}���U�aw	\4��%*w��-sCxUw�^��]�3h��QsŎF?�E�<�!9�$X`���0�&�(ʦa�|/w��D^�~�|,�>��2�X�:�M��z�h#d�J>�ma\�PƫҳE���X��e$`f��]�^�5��G���Q�נͤ��4�fQd����|����j������|#o�L���?�JB�T0`�q��qx���G������8���ҔEF���[�.�+3����Vz���9�>hhɇ��G?9��Gٲ1�e*6`Öx����E)	(��a�j�{���A��<
���БyCI@�M� �
w{]Wc�b�	�ͥ�/x�;^��ݱEF�3�(��m�����0�W�7�� '�b�dY\�y��J�/�Hp4��|fǾP��S+�7�6�D=�A�q�f�U������Y	>�*����F��P�,��h.����D*�ܟ*�.�/��  z��
�	{�rZ��BX�qc���H;�p%��7cɚ%JWY�K�Fc��ZF��O����D�`+qHlcQ媕U	�G@� ���V�p�+�����zG��ف��w��T�ܨ(	#�]j:K��~X	rm�`(�љ��C��Q;�8�[獹=�S�Zz]:�l
�3n_@��w]��i]x��4���j�t�
r��6c�Iyx��m�iwqO �A��L���pqm���|>�R����sy1u���	K�>$gw�'��>1����t��{S�+򗝜�{aPǄV��R𸚢�}�.��`����ü�ÁL��B��1�w'�M��M�s7#VȀ�H:��7m�zږ�ݯ���nm2��N&���ɺ�jj��3'.��� Dp�iC���)w�Ԇ���A� �"�|	43�\{�2���v}�>P��A��'ڰR(9�KG+6�5'�^~)��%�J)�wG�$;��9�ui�`��\��:������rb��@�;WsBz��U3�o��]\UV�޹f� �M��g�w�QT�&|3����n�	�D�@Y���+�t8(�J}ΙD-p�"XR���Z���G�)W>y�)&���z*X�2>�b���a�O��*�<<�ӥ�R����`��+��T&����G]���'�o�b��j���N� %`�O�T��|D] ��cw�G�@='��F���/]6��/����
�ԄǆZv�SD�ӆ�`��&�e�l�.�<���jT���ݷڐ���mI�L���yܸ�Ǹ*~��G�t�D?�dD�EKd~��,��z͗(�R�)��Lͪ������'�߱�ʖ_�J�������W|�h$8�V1�{RiŤ{}� ����ةl/Q�I/1�W9__,i���{xF�3җmWM�@!3<p�۵�X#�ԍNjUn��Q�IW.L~nD����>�֓���Ľ�b��H�T�S��҄��Z�}!?�(��yVѤ�Hr�=���w��%��)C`z|f�gG������Ɓ��#��lni�@<�#�;�BhI3]���8�ڒ�+W85�?ԫ4i<1"�a%�2	�q ��L�)�"؛)8��h�Z{��HO���I�c����	3ĸ>D-#���T������8[�V�!��{LgՐ��Y��Np��a��Ar'���slZ����x����@"Pf�*���뙂8M�i:,ç8��y�1q�f�����XJW�pD� ��"��A�?�n/ .	���G����i愳H�9y���#|��+�$dtGXN��r�w�yua�����}��$�Xĸ��vF�:b{�i8_��B�L 8�we]�g�zi(�qSbZ�>D2�'\QC����lh~����O��
?��E�~)���3Ih�%)\��-��$;�;`�c�c�	K)iS��h8�s�� �d.0�������hoTt0{�۞>���u��D�e��}*���Ap�*e�_��*Ȏ�sY>�ڹG�F���r�RT)/w\�ۺ	��2	������p-��7�����{[���T�-�k�X�M�M'�!��-ȫ����]_�kŉ���Cy�=(��}΁��{z���ko�=𶽨X�]���V�7�`��ii(��vt����Ǟ�r�,xLL ;���ɏYӛЍJ>����B���ˑ�b�����b{��S�$�O�G��*��9���[OӍ���-"�YB�q\���i%2��`}��j��w�-��1�PY��.��2�����I<�6D�zyYa�� �d�I+
�5��J�KȦY��Z�(�'6XI�Du�y�X�^[
��<#^A���������_4C����&΢~�{	�lR���q��h�.�/�{i�/yG�m=�E\FP�D�O��#@I7��%����J����ieF@�{aj΁h�����6Y�×�`���	��T �ˁ Mx�Di1f$;��㞗T�B1����G�M ���r�&� )�y�:0��eA�gt� �,�S�M�=�M �Sp8�%&!Bh�/�K��ɸ��g;={�=�^Wk �Ȳ7����J�*Ut�6&@�����<�f��b���<O���k�D�����{Y�)��=�PU@��Bm��� �/�?\R�aZf�6nz\]m�e��:��X1�����������Gsa��23��&�+#�0})B���>�a��FY�xu��w�H��xX��U���<�?T�.(<�2������V���$�LC0�6y�|�qBB�,�>R�!��)�_��n@m^Q*���#pu�+\H��S�.��k8>_��6�J��u���_]q(�c=;���:k��Z��JT���#�}�H��m�3\7悧�Sv�����y� �p|פ �N꟦�a��m)�vN	a������_\UB.ႠIne�O>c�7�.������U	���o�}��̙���4ӖN�Fp'D>�2�W	�EZU���a���#��5��/��,��
cvRs� �}Es��
v�OB���K�	��5�
3B�����h�jh�>�nR�/[:�׉�]����a5�	)�
	'>4CO���,����[}K�è#��hq��/�8��d�;�H�"M����"ͧ6-�!X��+;����u\�.���E#Q]�n��L�{#mYs��:�T��3��БL�D�zl�j�<�����lH^Vwz��D�e�@D����F���X�j��A1�*ӟ��A_AHOl�O��X�*;�xr�]�_��%�(n�E�1��*�SsA��E��W�
���	_,��6��@.� �(��J/y�K��D
�,�U�"���I�Ci�ȒV�z�*��=
����3��}el��A��f��m�]�Ii�Ch��NFpB�~}�P~����w1RB$��&�|z���sg�.���M]�cN��0�d�!�Hn��&h����P���=@�ĜG�?�?r�ʙF���m��b��F4 �d��@�p����N��ѱEqg�����rǌ{��/�yꗚ����#O1戎�c����.��d���5���@�Mpk�~��Lz�2E�zW�>�q����Q��L�d�ci�����X��9
��Զ��qԽ�/�ĺA3)O1mC�}�k���U�+]``lm�����WC�f-���YγD����-.D3�2Q�DK(�io����u`�e���r���I	i���7���P�
�i�ޟGZ��bV=6�r����b$P� n��b���`B�(C�/8��"2���Шm�= ����z�7���HѩL�0���b >!���?���ڐQ��xأp�b�|�լ�(����sX1��͵�:�n���'r�^o<�!4��U�^G��e��ߔzN�\W
��B"��{�q�X�)uteD��{�(塨sZ�ln�"�6@�K4���iT�0_u���'��$0�-��9)�'ڔ��ϲ��q[�
?�W�b*�Yxu���t���m���TKZ�E_"�|�vn�[d��:�X�&�;e�9)�Den�"5G	�����Ni^��u)��"�I�Q��9t��]�b0�尛�e�(5� �'E�\lk��!�-l�|̅�&�����-�����<І���mfh<��'���)BD�� �΂��u��>S(��l���Z�QP���q�o�H�9,1�
���S����!n7|��$n5�Gu%���PF4g�<��,j�Cm�>���N��(�h��;�sQF�$���đ�^�ڢ����Y���tc�����(�D5���m�eE�����8�ҀM���B�:k!ڊ{\�]�[J9���_�zȻR.��$��S�k����`CZc�I�$o�F�oS��ag�Nf�e��|����6K�H�~�y��k�?��G'՚q�E-@x��$,��B���/]�(�s�A�YDX�1���ޔ@Ć��K�m�d>��O��>@Ƥ<-[C5��>�',PvN8|X�}�
۝k�z�R]��ۧ�ߦ�����j�E�I,e|l��@�.!pY��sȷ��|��*�A��X9S�C؊�N�͝�@;�Rȅ��Ž���o��^NLvO�nO�b�#<Ǜ[�f$'�T�|�<�\�܎9ߎ����q?0@��������Xc�%�Ծ�M7��7RZ�
���Ec���W"�s)�a��ޝu�Bi�k _�`c�#����!�:���K�܉�/��� T0�+�yѶ��C���@���д	����:Z]��*���a����d�E��Աl�h�`�z=��"AU��1T��P�e������ڡM��bA��Q2>Ɉ���g3u�A�����װԘ.��]< p�@��~��=�g?��X��?�˹I�y�mT�l���ߐt��	�ĆLEPD��G���qIt���iJ$)Fo6�'�yg栳T����$�s����%�P�r(xb�������R;�����iE�%��䕲�x���3��C$����ꗿ7Ö�>F�
{f�x'�o�)w9+H(X�@�W�f�5t��&������i	���'F��AAP�+�m���MnOJ�%{�
��L|$��[fۭ�݅�gE(��~���ftR����M�6�*W��C���7=C~O��Ř�{ �r��gNPOp�N�c�m�T�&H�@����g�#Ñ�Zת�`Fb���W���(!9��W��P��ԯ8�ޏ4\F:`ڈ�7�2߻�Pj���G�	R�њi�h&I��!��V&K���"iӚL��=I!��v��&Ϥ'�Ub<֮{Oj��OĔSj�����W�Â�<&��sQ�_�Nҷ|&/{�
��#���[s�ĩ�1z6t�$�tP����:��ݗ�1�����Ne��(/���A.�5gt�@�[���2����8R�N�Е"[1��Q�od��p
4B8ׄs甸�8�SS��8���b͞E�AP�cq��K��Q\��� �p��0km��SA�ZW���?���JhK��\5�|�n\H.\�&3����w���\�*�OZ�/>4�E��з�M� ��x6_��ؕ:$�4��0;�m��+�R�A��ڢ(T;X8����櫣�D�Z��B����r�b5~��󂍊��9��N�#j�y|}\����^�&HQp��٘p�xJ�Y���/��N˭��5��W���B�D��~-��R��-��Y���p"t��苆�.��x<��h�}��L��u��)��5���~�g���Uno���_��fwa�?	;��{cVV-�Z�M�o M�vGu�i�Y(�ɲ���*����E�=3p
OE7�-4 g�n`Z���ë� ���MU�����z������u�1�EL�J�$?�A�R���~ !Km,M0�In}l�ۄ�X��=;��Hv���my�4|²�eB�v󵑠����)BT#����q`ٶ���WF��wҍفL��]��p�O͸����/��7������z�W{���+��	���F�j��2TJT_�W8�X��� ��6ɓ�]�������3dP�>�B��:ğ��JGK?#@t�>��ۛj��2��/��RUK:�����[;X贑Π ]�ټ��__�d1���h�0 � iY�MA�0�`�=�9���"���Y˟��3tC]*�מ#W�!��Ӱ��za�yJ�F��y]z����o�ǋD1K�o���U�&bp����]0/���Q6~�7\�4���s(��y>FC���s��,	G ��	/[$ ~Ήx��Ȯs����E5��h����R��"o[���Qv����dY��8�r�T>�ή�����/z��~�%�X�û�����{V^P�p�s©�WDJ߽��������L�����ջ��D>u�0[�e������a_(=��U�u�x���+��
l>\��i�M�����tY8��+5���\`�Rmu�db����|���=�����@�cKV���Oo�'�1�RM՗��H���p���������4�5�P>ݳ
��O��=/f���7�Y����`j�js�{�`q<�ڄ2�$��{fգ�\씀:���>�L���ǌ���֬^Zg�}o\t�$�嫎!5Z̲UO)NĤ���y
QW��߾�~|Jy`���_�g�r���ЍոΥ��f����A|м��>#,6m���c��iŜ�U�:�	q6 ���K'�I�v��t"!*���௹�=������N�]�w��0!za	�z�rY�N�6�FJFI^g��1;�@��NW- ŝ�dD
�T���m�\;?���_`��~B	�L���OFb���)�	k��K�SNʡ xJ�?�aO���u�
�R��z�C�N$��(��2�z��_&DLAG�!h29*���F����I���7]n�7|�q�4�3�P� Jjh�� 6p��Р�FL�Ե#�����P��'�3*UF!��bW��"����ǖ_~7���lx(��w�����%q]��}��@�Q4�²���B��U���ӭ�5I���H�t�����S�Ͷ˂�.���=;�0U�C��Z(���ۊ븺��:u?Z!����oӾ�\��D�5���f����џ>,.^��
l~F�����l~׹��+�=cEf��P�UHt���/кa�8���}��ݧ\�A x�%%��'��O]����`�ȵ���xy>0Ϗ�R߿��dy��=���bti��*96�Ӏ�64��y<�`E�ͬaLD��DG��_��ٷ��'�2��wXP33t��WRl�m6����{�AA�ʀ);���!�K)��ED�����Ş)&$glt��{*���g��=+��e�1��M~��7�[��H��\�덲��Л��d�We8+�1��U����ǐ�d���cSS�G��dosw���;�sK�<�q�?!�)����{��x/��f7��7-�� �]��~�G�L|�\�F:|�e�����4^�o.Ɛ����Op1D,o�������M�$��L�/oJX>��=��O�k�>:�����c9�Vq���>�д�t;��[��S�����A���_�PyiNT�_��	�����5T���2x{���C\�1U�^f���Z�Ѭ�v�?)kp�ON��2��U�=���֣�������3:�D&�4���iy�2���g��pǷ���ȧQ�a1��q��˙l�(A��\V�*��������� ���T���N�m�nŋ(4��pwͶ�-{h	���M��{^*��{�^
�L�o�%�_��K�����f`ǟa�U�)맴N�SD]y�%���@ s��~Pj�ᔫ��"���U5'	�$Z%��Z��G�T�L��#�M!6�D�}�e"Y��[�ex`���y�����6
��.b��2={�[v7Uن�N ��A���õ�x{�9��<3�� 酱��H���E��{�*��o*���R��d�N���%�ڥ!����Q���̹�llhg��`MY>D�d�����h@�V��缳�VY��A�0�G�Ν�l#4gb~˯���DF^t��65�Z���>�Wi�թ��j��|��7^-�N7�[���c�{�	8u�(j���'���'�R���%�^���iB@`,�Q� ��v���h����$�1���h���a�fU+�np�(ĺ�| U����~c�fŉ����͑R�oi��K'�ɭ��Q 1�g#s'Ve�ۢHqU������r�[���bG�$?�d�R�����.�`X����8{�yPp�b?�p]0g?��&��j	6��R�@ɐiSq�a�v�.�mm���I�\����2���w��X�5���Bj�R�P�~D�����Ru��L3ߍ�A2������`��k���v��F�!罬t'�����lX�Vh�+}����|��)З���wW�-C����/��*2D,�~�Y<�f�����Xd�A�Y��^�]�QрIQ�̍0Qώ�?�ڤ��r���"�iR��"&�H�J����ܳ�o���+�첡� ���(�N8W��Խ��s�B�[�mK	�S4�l�6���Q1�L�l�Z  �Ɍ_I<#+�Z��������J�+Pn�ih�#<pt;�g]���R8r΂�SF�(O$Ծ!��������m��'DTh�(A- ٹS����
	��Sl�t#E ��Us��)6��Wg��`|�Y�l.�h��g�ϙ�1�E/ռy /I0�LUZz��:�\�*�N�g����Ň�����j�j��F�ޤ�R�d�3�̨Jݢv��{_�j�%��E#)UP@]��l�w����浠z�o�R�{qsxU�a�5�Q��b��y_��.,8E�P��Õ������d��?���芎 �@�����%�$Z#ǝ���^�2�6�5�"r3,��=�@~q� �o<�[֣ÅѢ$�Aw�_�G�yB��c���"q��ҍ��j�[��r	2P�A(T�����H���
]t~�?� F_��}ĩ> C�9DRC-�@�Tky���-�dn�H��c�=���"�J����U�.Hm���ᥚq���z� ��K
��GPdm#9E��4_y4�QX���]��Fxq�2�tv��g{
�Sn����b�G���!<���ܟ�h�Q�Q�3��af��~�����1�)��Ɖ�R�:,=�ge�O���V�ý2^.'�������� ��k�2!�#�ڣ�� _ww��E)�b���,b6|7Ŕ�xג�-W�~�9�!�ٛ�:��X�6���eSǁ�v-*�P'�g�A@� �^@����Q�vyij1�%���������)�ŷ� ��SR�]�J���c���ʔRm<�C�(g>O����-ȳ�NS��Jjc<ò��4��C�@��7CË)�]����Scqt�,-$����e�Nn�V��hx��?��s]�#��s�w�Xe#�����g�(�xp^�P�	�c�v�t�ꢶct�Q�0}q��aJy���;:� �IOb>������MX{�� �h��]ԋ��0F�6���P���OR�nT���g�F�'�2�$� t^`�3g����XYN����;5��������� ��/�F���\o�MjaD�J��VG��sC�u�Ekf��B6&�z=�m���+g�u!J��ɫ����������~����>�nST�u�Y�?%s�jLَ!Z7/�7Q�`�?S��$>a�Ī���U#T����*�DT0��V���0li&YG����V��r�bpƊ�i���_��g���$̷L�h����4�P�m�>�m�����Y�/�E�NCL0M@<�J�q�8�/w��]ܼ	V8?�Ca�@v鋊��Vܤ~�t�ڦ0�ͯ\��=�e��,�����eR�{�-�~�ڝ�e�5�_�%	��5I�{�w��N.��Be�?��/�vjp)2�9��\F����ċ�N��s����:�z���rg�!]�ta���i^�$J'�{�p��B����������6�,A�&,�{/���-�c��g�f�����O�����\���ɹ�=$5�v=���.���'4�	M�ը�0a���.�+�˲�n2Z�~�`AG�||�����l��@|P�el�X�	c��3��F�Q�Bg�P�b"m����*�ps;�RW�ۗ���`����r����C�Qg]���ǭ�w�����{Θ��@��檃�٢�jW�ٔ����?��Z��A���� ᎚?�9u��--][2�XN0��N4��bL�9�w07����!��+"q;U���F�+�,T$��}�ڂ'E _ȝ㠐g]���0�1p_g\B���ۜ���l613l����"=]�7(�[��[V���D�p/��\��^ʲ�X��D����]� ����R_��3１�\\k,��7(Θ�����P�q���5?���UsJ��Z!�^1���_��ɣU������EK�٪j$�}k�}���i�
�/j�=OT��5��ov8��L:�^i�1�ˀ�w���'�u�Ү��-{vg�9��,��w����a�Ƀ�ZW_Z˪U�q>�|��R�l��}e��$P���Wt��-
Py��	�	���i.���[0�{,>Rdu�j�v�	�4^�E{H`\3��V���ϟ���BN��fs­6��^P4�a
,���׽�5������]j�Y��5.���$�nMV����G�~xS�����F̊��N�\�g�t��5U.���t'����@ιd����-��u>˗d����&�� ��@�2�N���Pw>3f�̏?���*CY�K=�@`V���|��r�m���bz�v�U�xZ����*���9���SwCx����nQ�-��QUm2��2���V���e*�j�Fú
Y.BV�YH�oz�}&����ۗ��&�񬺅kKc��X+��e턛h�%�KF�hla�Ӡ��f^�$Hg�� W+Y
�uB�6�	�+�4�-�b^����Z�'�O ( ��<�&�dD�=udL�g=�$����x_�Ԅ9;�ء�@�υ�X�7�9�[���8??9R�g�}�gW�#&&�� [�^y;Dײ<yc�bگ�M��]��d��������屸+�Bu�$<n)8b��zQ|*mj�q+�= �R�ՕO���.'fK�8N��%����#� <�o@h#m�y��@y)��F��L9�C3�	�iH?i��6���K����34ua,v���2�hv��I\}��Q�F���O�l�U�/.�z�t�t�n(fS���klc�L�=?����m��b_Y>�P�z�0�-�l|E1��#��/Ah���M�I
0P��+3s�W��U�|d�t�U�ͬ��irc ~-�J`�J��&-J�N����wf��S�A8���R M��x���H)�D�}��kʤ�.{/-�X�z��͜sz�����Yx�\��:a7�Ue@�O�ϭ�V�+���rL<��RWX!�A7�A��3��5I#�2$2����!��ٮDz��X�=����(5�����&M!s�D�|�8�w*b����y�}�-e.�P����A)���h�iF���|��&�Ї�)rF�ȃw��H$�mo�M��?5kꞣ�ψ=$�tν��G���~��p�xz��Mꇰ�^|,���	�*���'47h�8g⣑t�z@HPɺN t�'�����Z�U ;��9v`��19O}���L\�ѿ�T:�Y�{�M�e`�T!�C��� ���&k[@����h�����dsc좩��u~�pؠ����֦-�����c��M��$����0jDּ
 �E,}�ǡ	��ҋ�Ì,�e��8^�wiDy�R���`c� ӨY�<���� J�VD�x��79�6� cbU�<��h�k��Kc�P/$Ye8-�}�+C�<�?T!�w��Ea�Z������y��ö�I����J+���r�a��H8�4���(�-�b�WA�X��ηqo$>{�������#��=��Ag3���eB�� Rݢ���\Υ��n��M5`��� ;YУϥ�X9�.m#���~줧ΧAk9,����T�����e L7�rc�$	V�PS�\ʣ�l1L���vS��&�渕�(�sr�n"JI[s{Ԑ�t��;m��W��i^n��]:�B��j��x��	vx:9��ʂ�\(m>�R��wk�|��Xz�+C'5'�V�g*�ba=k�8�+Ƽ��1�9�;(N8<���G$�WQ��H���
�}f������@�O�0mE����>~G��WCw \s��+�
(�o�(>K,�@�pW�d�z�p���	����/:&��X(�-��|�a�χiN��ܦ������N�7��j��q5,�o�������eߊ41�n#�Io��������|���ngm��S`e��Ӈ Q��/31�f˃�O���61�<�e��-�ȹ�� �W�?���sh��ix9����L�b����4�q����cw�p�����7ߥ���ѫA�R������aajL�<-�/jq�	Ӯ�=U;z?Q�_�K��R
���r:휞�/G��Svi�>�p��������j�h1i��j�\w��VT<���p�%F�u`F��H&1ΧHE���v���� �rJm��AI5�%�Wlj�290>lv|��͙��Z.�w�H�I�e]�ǐ��� ~](H�$G˫�}h�D�����q��y���:'4hB7%8bzT
�}��<=��T�k�}��+i�e���m��:b������g o����*x�0ED7Ȳ\u�20m��'n���-A�K>xtQ��v~�Nq���&/o�z�kw�\/V�^aH��Ϡ��ԩ]��2e�#?��j���t����7CuF���elf����$�!�7�_.�����&����T�<�6�9̏�ҬǍ�����c�2��
^�r27�������dQ��,�	�}(��8�uղ�������%R���fT���9��e Q!�u}d������#(���s�F�!�k��Q�O��k���+~��h4���|p�Y ��l�9��?�|�;5E���e���>��<�������7�6MD�O��e���|
�`
�gB3��������o$��5�S����� ��?P1 &���}6lM�-�h���� �[=��f���r��D�jD ��ʜ�}8V��R~#*/���*�:#��ߕYD>i�M  ��.����,�W=�ɦ	BN�쵊F�: �������L�[���\YTʧ�� ������kXo�ү_n�S����������{�G7%��ZS:9UF��Pʐ*>��Ru#��^B�W�
�sq�ˋ��.����NP�70�۠�V�&��'�έ�6�}z�%���b���R(ἆ����s�:g���x�-+"����G}|B�hŖ|����n�&�s��
���d^��\A�?&�Ur��Y�R.��)��%��zͿ��j�.?J�� �}��`�.��<V?�杞d�7��Ű.�㓌�@����,�2:Q�B0f/3=������?v(0n��nS��o+k9�t�v���9�$�fjm��h�)���t����f��"�r���3���e�vV�]X�H��ͤ����KA����7g�-�e�����֏���ݝާpv������#b��
�a�c�qթ�}©�a`�Z�?J.a��4�����sx�O�_�s��c���3�\����I�1w�LÛ>�6�Hbl?�Bo�hQ��a�,�l��J��-^�j@�VW���WFh P��Q��N���v�d�������<A�`ґ K�֧K Js�^"D�zM�@�u�h1f��̝�)n�NY����7v�cJ����*�r��)Mzєj�D�tw����:��t�Ɣ8��{��*���%��e �F�J��Eo7��ʦ�8mv�m���uL#�Y�8�$ӶY.��3Q�w�0�.����je�c� 5�Ӏ�i��KKN�U'Z% �����8����@E��|���U���wEj<�.H7ȹ�0�
�ś��h�;a��	�L��?���l�z�^3M�u����b�?�l��'OA�N�-06�ܴg�;���<���;^�U�Y�G�3�yBc�q^��� ����E^�B�|6a�D�S��h����B�������$�H��?����O�v-᭺�'�(z�Q������2�����w���-I��*�k��l�r����e�?����o���>YbE��˓��I��H*�	̈́bW.�_�?��5J����[#�pن�r��gL��M�
��U�mbh���|��K6m�(W���d��!��(G]4*�/f�ڭW��X��R\ڂLB��Ժ��1�9%ua�*k��^h ����¹���{B��-�t)�;2"��ݿ�NB�45 `��4��d7�&۶h�V߱�%YG��&�(�EjYuƣ�?K2�g��֡�?z�@�ʹ�v|EIֲ(�������!{��{`�TĄ�ҩ#�ƃh`l�򇤧��b��~��m�,`█H��:��Ȕ�1G���.�׀��x��c�"�{K�SG~.W��=*��l�Vr�~,�mE!{��j���|��$Q(��)%��"����6e1> ��6���{gw�x�/��h��Ì~q[����B�gO���x���s�$�݄d�f�!3�{*�t<pj�q�T���=�8v�Lw1,z�@�jB���ͤ��(4�J'��ew��{��󸩠5�0�`P@�p�����rHc)�tj��;㛻fI$>��!B@[��AW��kj���l-B���,P+)w�o�� 0����M�C>��ɾ��e�$�-�;��4"��{��wI/����h�yT����Rh���\X���KY%��D@J�U�<ҿP�T|4�  QW��$,�C��Rj�[�J�h7r{�{�	�W�<?H"B�m����@�M�'���	�SB�>�,-h&��Y�Y6{V3�~A�ml�	Hl�Z�'���j���+����v��<�f|�E�9��s8�s�]P��y��SU��XC�K�.��:X������ANLg~N�S�3� Ri��(z��<Z�9��}�6�<nϼ�bp'?�GF�Q�,v���aHwk�(��&Q��J�>����d�����Q:����/EL�ҧ�1C���U"�q�Е$/K��zu	��R)O ����b�-G0Pԏ�܎pC�\�`!R��~�G�s�RJ�zt��:����^�%�Ş�jS6�^r��;?-+Lb�����U�!$P��$xv�	�ng.��/�xflD���Re�b�7�{��v�F n6�`3�F�97͒��~}G����ADj0`K�{��1��=�YZ�@�"�C�5h��A���I��䂩������'���x'�6��Qkp ����{]�J�i������p[|h�v����2�\�Ý���ɔR��H�F��p8�6���MK\��m�l��(T�2�/�Ͱ�ˈM��ʹmO/ż��^����
�M:s����(�Lh�qc3�*~O2�2py��Q0��#�+��GY�D�@�V��~:ۺv|��?>�i�� 1���%Ҭ������e(��eOf�!�{h���*V��ć�Y����[�uLa%u�n�\z.��ܳjN;����<))FY�Z]4��ݝ��.�εFĆ�A��&�
��8e{���[4m��.��m�(<g�Х�1��=�Pd�ʅ�r�ꮏ�DQ�FÛ�J��#�c�%
]5b}Z�M%�MZ ����T�msHşG3h���ѥ﫟��������X˭�It1B���_7{äK��K6>7�QJ�Pr�����$3#_>��]{��bv*�f[SGZ�\�r��j;G=��7��k���@�Ό�����&2�u�~p|���������[��_+�&���D���}��c06���w�v \�� _�a[��=�*�`�0���<�9��:}�Ń������6�!ؤe��9�Q�ƊM�`�j@/�*�$T�E���E�K�Y
�_�^�a	9�2"y�S��#۳TOL��/j�Xt�Z8�/x����|5	��:�Yi"���U��u�̘b��Cm0Ms� ������y��4�y_G���t����s���-���N��l6�(p���6S+_�����}�/�jV3�[
7��3J��\4v�Q��vo�p�dL��7;A��{J�?�����>Ixb��
#���&�j��Bn��@N��뚂.=\1�W��)��)⌠>�f��1����-V�
����q*Y��r��h�vai0���He�g^���.��R�#�VR[TFQ�,�h���T���G�m�	e�3VS	�{��v�ힵ�ؙze�W�.�#Wzz#��!X���m�X�6*�[P'�7T�C�d���(�����w��\�fA�S��w�4���&&���!̬��h����)$��=U/�6R�S�O��|�=��kG9�v�n�#\*4\Ҿ�~���!���ë�RY��E�}��~G���:v�A\Je���z_����|�K�7}�#u�y�֥|kbx�x����9��ّ�'x�)j�,�oFz�*�p��;�R�\�e��P����1t?h��.:
��#�x�3�,Cx+���#�Ux-�ي�.9�n:����2`0�9�x;)k|&U��"���6��D�褖���
�s�f*Ň�B*�pٞ0d>J,�(��V2w��ez�(��N���>di�S{�mݫ��7�M�9,��.����݅�� H{�6uԖZ1[�.pHό�:�ځ��z@���eg�Ԕ.E^��*'��FT��P�GWxZ��@�0S��	��0"�dS�
�)\�]3���w���}�@�#,�����+��1K����u���Ws���*��C�⥅.>��yw �H���������_�t�k$���Ɩ�@9އ�`/�s�/�zȿuM�8'���Al�5�ݻ��*�ɾІ�Cs�ܣ�DJ6�3�)�S�Eo��tkSa`9Ųi^���V����\��#�f��y�.(�S ���X��`R�`	���*S>{6�������L��;��-�:�Ð:��3��׈7�M��W�H�z/���;�;e��@�:B�� �8��z�e<���~sWƴM,��n�y���2�.ÉL��9l�fX�ݠV��J?�����."�1�F6�]s];(La�����e�<ۻ�6��9�Z?&q�	n��m�C��Cd�.Gn��A�πmd�S������'}5�����:8L�Dbe#�{A�WD���G�^/���`������ �a&�G�|� ��"��.W��V���ϦEɆ$�;*>"�����;Ɉsn��Es�I75㦻4����7Tw^��;K�iX�V?̉X�b�tN:�F,�(~���'���	>_��&����������D�I�#x��*d��"֦� kaԼJ`�i�����z��Ju�n�R�%��	j���W�!࠻�x��VS�����f-��yi4KY)�EL2�c�ĸ�ۿ4�Q'�)�����l�E��I��J�C$=eъ�I%���d@	Y���*'��k���q7Z�4�-;��rM�;��5�����4�^��*B;O�ǛI2�X4��� �C��sN�Z�C�J�S"gaH��81���u�׆�pi���El2�F�|����+P?�;;�>���C�f����ЁO�$.��6��C��?R�b�W����x�i�Ft6�9X.� ��K���9��8��"g���;�&D���yJ�Ǽ�y�GE�]�ZHA$D���60��5]B�.�t֗�.6�E�p�P[EK����CU��6��b�Eu���I�Knk��y��:�S��EՆ�6�REn�B���w7�d�����U?e�Q�4āiηs3u�g0d��D��I���?�	;����*��#6��/��(C�Gu����AxI���'?'�JG$��ۣ0cLI��RI"}��d�Y�'t��(�TG\Í��9%��@<\���5�:���~�%m��צ��)Z_9 V������6f���pPb�<��pZџXv��M���$&팦l4J����%0KS���)� -������4���sN]�P(��T��ȷn%i���zK t"w������_�S��~N-�w>p:�~M������j�1������.��K�1�������c"4���^�Ħ�Yp+��&��	�(�ăʈ�@N�AM� )k�����r �8V�k��BTm����أp�f#*�ӫ��#_�I@�k���"&Qd��n~z]P"A�x7f: �C4^�S���5=C-@g�P3l�~�Å��h��z>��I�`����Z����?o�NG�A�U����T;�/Y|�"���#9i��L�X͐#Q0<�I���W�Mt��>�v|����L���|���!Kf�>p��aR {�߮?1��(+� x���B���+/2N��7��}{һSȭ���?���B�|�\�e%�����s�&L�W��\���z�� �IX��.��_a��ا�+H��"�O	JgQ�Cǔ��+ ���.�v�Fb J�+�����b�-�>��n.gq�難���˶
�"OK�;��r��������_��c���t^�2}���w���m,>t�����V�v�f�d���f|tf���m�M���`��O�k��@��8�c��n�,Z�G�d����d���	��4y	�v_�J�7�b�a5	�O�;"tF��单(�Ϩ�o��ڊt7\��x��ہ� T_te�N����+��:�dX����"b�״��/�8d�Ok�����4����}U�r@s�u���{	D�[���<엨1U� �ǫ{fQ^pJg}�lh(���vȑ�ϑԇ�>����&_��J)��p]��@xՈ�K�Ϻlz[9�ȯZM�5"7�;ĕ>B���,��)a|�
'�p� <:�Y5�A�`��92�`lX�!a#��K��>Q�u�Y*���dM�66}��\�$���6<����)� I(��[Y�D>�^�~ԡ��pŝQ�Ą���ct�2C4�{���u�9�(mZ�F��̉��N�p�DԘ��
����w�.&��:^�/�h�!q�b��ؾW���������'�`�aW����S�4�A����/�:
���}'�N+㣿����Ѻ�{��tiȐ�)�$�ɭA�d/8�/�D{˳*�լ�K~<z++rY	�x�˥J�G�*~ R�qk�v���;E��
�f�o��'�1�=)�Ԫo������L`Z�?� ��v^� h]m.�L����^`A��}���l.n*w]��<T����U`�p�@F��H7��*,���6��������&��N~�����{�f+R���SeV0k3�6$�����3�K��A�Nѝ�E�j�I���y��T.f�,�=���X{Z�	'��cry�f4�6���2 ���mrD�g�v���� 4���?�\F�df����x>�O�Ȁ{x��(�A�8_�a�a���xs�r���O�)z4�~�I��!*�=��.��-]�ЬN�+ٚ6!��#��;B��9B�B���2ͤ'�8�fɠ(Z6$D�=�x }��ǡS[ob�}�B���PX�t���d��6��t2�%M��,�
���E��p��ӓ�:�����/�e�n%y'�a9���Ӳ�>j�z�M)�g�6_>�7&�}��02�W��	*�`q��8F�<��}�P���;��x��!�W)��Z4�]��6�;�"��X�8x�M��Y�k�i]f+���~��_��HfI