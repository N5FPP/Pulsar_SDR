��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@���$U[H_#�/8�y��,��F��`G�m6f�f�aiI`������tC����dl���=eZ��^�٭����B�FYĸX�G�����݁�]}~�s�cC�_ �c��2)����$�a<��d�6�q��tӏ�ˡ\s�$�L���Ÿ|^*��g�@U�*2�X���2��^�:9��D<��;�h��É}����a$;��몬g��>��W��iv���o�ăN�G\\�[�4�������W4xl��0�;O���V^��@��l5f+��\�&�7F�CqϮ�Y"�� C�T���/��Ƹg"���l ����~G�_y�kIe�+E�9�>Ǹ=�oWS�|���WV��P����������L��΋I2�G�r	y�i&�l��vЦ5�o�#����T�WrkV#��+�ڛ����C��ɀeG31>�����k�\�%�̶�@J�%A-�@�'2�}�0�΋ha���RN;zy�Q}N��5Z��}L���Z��¼�1<}M�����g�) $�8��Ρ�g���}E����G�@).�b���L��<�1�~:�~"�S��Y�p*-��^(Yj�����k��=98VK�ϲ�=�Zhy��� �#��_���c���~���YƯXrh"� Sao�%��Ƭ�;���cE��:�<:���6��E����Mr`2C���L�g.�T�"/)(dAX �B\\�xG�� ����	��r=�ى��x�⿐�z{�&��!�$�ȠC���}���?pEp�����p���р�e��Tu�M�@(���v6�ɥ.D�{(��Ķ)B0�h.ˢ�ا--��I�OtQ��I�ǧ�b:�ot����'�� �AvY��ɲ��c�Q��h�v�z�Fo�6$�ǧA��h�;�X��?F�4�E���j���X�Qd�i�� �C���¤T&=Ò�z#������z?��:�]q����Qw�۠Z�]�i*v{�-��JL초�+t���������?F�JF +f�鋩+s ��bg���ȬF��/�q�4����Hnl�!
�ǘ�;a�CUﶜ���|�=�eQ��:�9�?�뭥�n��IaUj�	Z��ʱ���S�n�o�86ν�nȚre!�~�Jm��F���t���W�X/B�ڼD�מA�1�N��ދ��P�L�N���U	�34���/�q�kvB���r��m�d�,}�c(�70x�!��s����	�B5-n��ռ������J�|�u3ҵ{�n�TN/	p���m�I���ב���0����y	�s"ڇӲ�!��J$�'��yΧ�9�\9+����� %¶XF�n��k���I�'+�io��{#��z�Mk��g���:,� d��G�$���ڑ��e�����T�5���hp����v��*��I�������1�S�g���My·8���؎�*��:Z�s;�J��fߔ~���� 2)n�CG_9�dn{#�^P�mw$@2 N폥ȁ�b�#�rë(��!Ȳ�J�^�@*'���u��p	do�ͮ��w�~�[�ɤV�!u�����k��g��?�K��t!!}���yk/`4j�>�6M�@�P��Oud�;����}Y0-T�E�w}/i�/��tI�P�˵J����g�4B�D�װ���Ǡ�_��W��l���"q� � ��j�1�Ղ��k��.y�@a�ZbG����gf��'ҁ׬����ro�L�/��-��OwN�m�Z ^l�:��&_���y�Y��=ݎ=�`�=��<$�[i&�{��Dg�u�³�+�_r�����T=��q1��4�C)���]�̦�
,�Q�!��e�������T[����Ր=�v�#E}ٝ�Y�A��u3�Z�O�f`���B�a+����r+BE]½ko��7����k����;�v���o�H���7/���*I3a����{�1�~[y�'�������^�õQc�u��_<��?�-*z>����zu��[b���Ghb��m.��@�k�w30�Xg�rI��:��&mT���\K.kBNέ��N�l�����`����ǿ�Up�`ި�H�P_�(��s�ãW)����Ӌ!�I3=�HnC�a���U�CeU��WvƝ�@�i��4����"wlu~���<�G�'�x��R�u�Njy?ݿ�nnd93�5�Z���V���W���"(1��y�G�fJ�4$`Sz���@��U˯[F�L� �"��vrE�*��3{����!����:ǈ����3{I�z@نp���=(p�!���c�d�	$v j	IL��.�e��qZ)OR.Z0���L>du�۠�BwZ�� i��
xۯŸÑش7���Ͽv��R��\i�9�
�9���,��k�!Ԙ[���O,%i
�KXs7���۪�#@����?�A�1�b/��+�SG�I��"�%�ǳ���4;FE�2�]ʳ���9��qƧ���ӌuD�H�To�b�\�_�\Bv-�� $�k�I��:u \�7���h�����;��]���SR	=�Mg������7�T@�B��2���h*��ګR�8U 'z3�K�Z��`(I��F��o��X�Jd�����k����ˎ�_N>��/�~����	�JH�xB�.mBOkr��7
d���x�)o�u�ʯ��ƿw�e�,�l��s�lj `PQ�_�:W8v���{ȝ�����S���0��s�K�Wվ�N<H�Z��۴栜OS�_T��֦2�P`�o]�IqX�����D���V{ت�:I�fЎJۜ�X�_�%f�\����(+�͵�%2����1./�:��I:NG�W'����d&	�rx1kM��.��j�A���.��	Q�:�KSIu�@e���(]�s�a�ܔ�')�@�^�J��V��
 g�#�A�6"Ax��0<�*�d�$�:c�@��s�� ]@Dk��ӂ��(�ّ��B���H�)�ۡ������
�V�}���!]}.T�#/��R6���%<W~Ql���`	.15���*˩2r��<��}$���s���Tx,�)L���\���'�v��nEq�ؗ�b��q��t_Ö	h�?���CnSסf-�|��_B����/�t�&��N҄����(�|+(���;����q��R���i�R���j�T��JG��|?��
�/5���$�>h^�PI�#�����4��I{�]%C�fHϾ4u�7n?���{on/��*�D�s7�����*���ts������<W	����cG�1�(�nL��4�~�cM&:���X;+��l���7#E��A}�e���>s
0�t��dǉ_й��~0w.�/; f��B��IĪ`[Mwah��`O	=����c˘Y��@������{����ORz�C���m���~��b9@�����s�3�ϔ���d�dܞ��{g04Y��+z����	�������� ��`��]�)}�ْ������%U�Pi�Y�ۓ2��U]�N:ѮP?3�W�.� ֺ`��I4E�y7t4 5���W	 B�Bw`FzG�}�����j�{��Ҭ�WQr���K:?��5����R��������aC�,n=;~��}9�YP �wI#[�qI/*n	B����[����S��v IiN/7�~ZOÍ�w�uW��L8y�eJ�8�f�����Q}z�<�~��I	�u�!cy���@������j�oj�3�>:�)ox���Ǻ"��u�bq��`ΧN����w���Q��l#%vd4�{)pM:�v�O6{X�j�v��=ZS�Ǯ4��E�|�{�}����4�0B_��gg*�hԌ�u������U�h���+h�����v��#y�+F�ي��Y�MG/��Ax��ȶ�
���G��2�rw�a�|�r�ڗ��I�Xh�}��=�� �J�Yr�M����2�����Q� ��z��=�U	0B�?�Z���Z4*³:����`2c�u�K�VL/
uI� ��c�󃋝8a%���*��'}&m�:��1�����G�`P��#AxK`�pb��
������^�B`ֺ��~�bR��I|.+~�\J�j�d��|�w�Dd��:|k�H��ui�,čG�����a����o�	uP�$�N�� [�pKT�)�NeZ5�WC� U5�FG�5����O�ņ9�S"zW����P��vL#H�YkA�(ӷ���eQǓ��n�I1�G�lL���$V��ިBH-z�k�͹�o�y�;�lW��C	\��̩μ�I� MR�L·w>�m540ymw��M�W��#nn���?%Ȉ�Z]\�K�����7�?�#��U^�WeX���`E�Xb7�6ڃ�cS1����6�vHv:<�;c�i���G���\����}X��wА�L����Ԉ�r)niT�&����j[B��H_B}�D���d�q��<=3�����.��)�b��0�����A��˥cLλ�'|Z�Z��b����!1���^�~��a��28��Fst¯���qe��,�8���JH�ha(/c��!))��R*�>�g{�>�Ά��u�?���7+W��ȡ�Ϩ�HE!��y2@��)�[�z*XM�V��n���=?D����4��N����&W!T�<�&��"����$��k�O�d��'�9�7�\�6�tr}�x!�E-A�
^�������!�7�(T%�%����.0C�F@ZD�8��s����~���2��!��e���^�C,^Ts��ֻ�d���^C5q��n��PՃ�# �� �n�ٱ��@Vx�Ӣ,���)>-
>�Ɛ1"8�(���˺�@d�����r��?oN|�$�RI�5�(�](J��l)Ɠ�D�#Ѭ[> ]�l��<��ɘ�M e�i
�e��������t;+H���4|]Em8]L���)ʮ�Z�>�.6��1�΃�V�p�� x�~�;��q��aSyk�B�Df�L֟!��kcx��W�ȕv͒ڮ����D��q�DvA�����kOO#0��}H8���L��#���N�^��X��_!��O8hn������=��:dL�ʳ�*;K�R�^^�}�1�&�v�爇!n�1SY�{�x����ǻy�aX�'�>��9�UQKU��7H8X?)ΫF��v�=mA~� �n�-�F	=~�1L��ݬ|�k~%i�g���/*f:�0�f�^k�ω-Ӑ��P�[����\l�ٖ��Eܚ��F�e=�zvM)�Ƈ��tZ���O|3���=!D&l�;>eo��$?|�3z�q�"��ԟ�Tq�t�	�������������ۏ�(�,Y>a��
%��N���E����U 3���J�$�Ii�s/6x6e�h>{�T�����r+�K<ggbD����\��Ξ�5�E/=��s��{�7�ٓ�F�ʽVa�/��x�k?�,P�����{J��IJ�l���0�w#-��&��J���3\�d7@-�!�7�=�b�3�ꛐ��2ŋ1��������ے�L67�7���m�WJ���)������|��Q?�7�#b)4�+�+�U	� UYFH��j��śy�2$"j�d��Q����Rp�	uh�Z1}rZb<��Pg�՗=��́�`m��J��]�����A�RH�a����Б<������<�$ص�#,�{�xC��s�!J�,3X�F���q+u=ؠ�9 ��c7��be��n�J=�Q���]�q�45N<y����X�q��}�K����J��I�xR��J,n��q�X>���,"�c��5�ϴ�����8s�.}ڋ2~ �