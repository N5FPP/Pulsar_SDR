��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4dտf+����ؐ��7&Qa�z���m�ࠧ��3`����8s�@M�4�s~��B��h����&����YND��b��1Ü�(_^�[: Е'�GK���c����i�};<���k�.j1���a�����e}�PN��_�8���>=6�eK/L(�#�S0��C?v�>�-}闌�=��b�7��-6��ָ�	���8/8bWbR�рI�5�� �!VX�`�H��-jw�_�W �T�2��@�w�E�ў����q��Jx*YiEW�f�<�P^���hሔ]�:&"u�Xg�ծP��齖zd���u`�l6d�zh�L�Z�͙���z)���i2NR��uoݕ�W�y�U3)}�C����7�g��H+�X��6��e�f
��,���@2��v>P�ۉ+�\��@v��$%]�+�����M#��.-6`�F�ǹ���X�=m2����v�]���[�_>Z#�2�VLXW9�{���6j���r<w5 ���h�^���O4��0�;rw0�1Hb�&�q�	@�ˉ�9Ȧ��|b�pJr��^X�]�dG��)����<��"߹H#0�.b!�ޏ�
1ir�g}��u�L��Ӆ2.zb��pY�݁%��`���>��}���.�#3�e�(���*���Ѫ�����6j�S�&��vv�3���J���F�h;{#���ql���[*������b��:xh^"/��D�����3S (�G�xC��èv/�n�b����W�|V�,�\C�%������1%�,�Y���T3�W5u��J����ډ�E�&��z�
K�� -�8b�\�T�0&��*�Nk2�N�0��M:�;z�bӾ�|����-��փ=���[����(drl��B#�#��%J
�ͯ5ׅK՛�Pe�/^2�'^25�Xs��6�1�:��8	��ex\�Q�m5�oL�gzK��P/X΢F��~�z��c	y)�:�9�-������#<a�x�XⲒ$�3؂�9�����he��di^h�8����S�3�����2��xko����}����& 1,�������mM�XW�M����G�,�fMA8s��LQ$d�?���p��#P�t�e�a{��6��PD]weh�0�*Ӻ����6_FĜ�X��#`�oV��V�+�����B�tC��x�#�KT��A��a��N�Sn:G�M�9��M�}'�bK#Gv��3a�H,)�m�H��+}^@�0ߞ+b�w$�~V����]�zh_�K�	шt1�T�ӭ���O�?̱�;'љh'%F������m������c��煶�{9��~x�R[ℑƍp<����+!4^��Jy��}
���B��(�dv��3�$P�TT0�pAh�{���V��Ov�W�C��Bu��AH��l��pE�'���+�^�'8U���=3B�̓�_��q��%ef�\S�yb�8��HQ�4,��B��KI�f*@8~��8%ɧX_@��~˘�Ej �﷫(�-����_o~T�su�/3�Hez��p���U��p�X�َ��g����w�����6�NlP�n��v���_�Y�����3�d��I��r5�k��	�J�
��OkA�EU)1�= �h���a]fY����\�zS�ƯW]���c8��Op?��3	I#�k8�_]���*3����X���%ya��:W�'�d9�ً�����lu�蘤 �9]�a�WC&n�N��$�M;�@��bw���$��̣s> �e�ԥ�\�+�k��B��`E���V����`R�ᒊC�r��}��< n��[�Pm�z&o�5a�'V��,��/o�kgh��;N�V�U,gc�m�_N��u���w�,�yG���ۿLd���sL�����/�W2!p���_��i?K?.��0_����\�L��'����i4�ҳf#�[]4ܙ�s]�U$��/GZ
 \?|��V��ԏ��9׽�I��w�&\���*K-E@��9}�9ުU�\V�W�{c��h9F�m�·"\2�sPY��8�|����q�� ����v���O���0;��JɩDqwTo�c&�z�̓��ۡд�x�L] D�7^��O�/M�B�z�4��f��� ��2�����p0�<� ެu�7��oSx�s=h�OZd��QF�)��y�{����Àeb�Z%�����������r�nl,�(DN�f٨O�IJM�Da��	��0Rk�d�n�2����~ �)��J�^��܏O	��qI���E2T'^�]qQ����Ѻ�� 4$�7����x�O҇<�eC{W���A���h#x�ު�d�4��7�h��T���z.%=��p,Ysa��J1�-���g��'0r��,P{�((£�DD;Ƣ�;��=�K�'5���<�e�3��*�������U�=O���:�ha�Ց��}�0�I�k����e�hc�@�كT�s�8���S<���5i���v:Ŷ�`X�3�20��� [�,l	��+u�0yi��re��B�tom����|���˯�Þ�����/�	y��$�q�ŭHE:���[~��\�up��؛č}:��&����`������_�3��`'�w}pY�6�M������6�B5D+�\k�v��f��`�$*�|Z��7	���=ߑ~�3��- ,7�|�~�i�Bd��JTE�dJmb+����lX�b����)Dz֒0S�g����;�P^D��_�F�, ��V�d����T�ʕ����籔H@���h�Z&�r�x*M'0Md�-���K���� �`q!��B�w��3���0�k��9�� � =bgJ셈a\��`a@Rӆh���fb�*��#9Պ��Z�^?Lc��/������ܞ�)���6�$a�/w���	]tP��i�wr_�H+P�#�9:?/��C"����-��{�t��KX�2Kh!��x)���u���k<R3�"B;��"������q�\�\�ܶ	V�6�T��=+������e�h�@z��E�$XT*%
I=���zJ|�!�L��w�b��ŁN)Α凙��Y������Z��?]XN�1.���	�lF�=�³�"��:�=��8A��#�t�"_��EG��<{Q��]O<����h���-TG�=�{vUn�G��cy�T�;�e.c��J'/�3�����W0��Q'Ӥ^�j	����O�+�?��u��}
�us�ޣ��Q��3���L�I���P���h�ȳ�T��u�r�H.�(�WShXy�����_�Zs���se,��AP�YM]�M�8��1N��Da�俔��E���@,���U����t�X��m�H�Q�`�Ѱ��
ǒ�_R���9Y��d�S�W��|u�r��GlJ�D�/�Z�I�Wv W�2�=�����m�o�- ���G�����Ƕ ���0,��;V��KJ��GI���Ë}-�$��ӑ���h��ct��u̔gi��H�i����M��&Ե7r���;dӬ�C��#'�]�Jae��{R�9�����t��k��y��%��w9����v|�h	��+���X_���@ڻ��#�5X��ԓ�㾶�;Q4ͬ�Կ�F��D#���/.�0[��*ƣ:�Zt��R��r�'J������atP�l x��8��c�5 ��iH�|GUr�9ɚ���2��a��4gp����0�(��{`"	��l�C��n��R��V݉UZ&l$Um��!%�"��m���X�����O�~а�D�U���LEgH}44�a�Q�ik	�!Z,�H�4��,�ტlP�� ��HK���hJ��΋pVP�J	��#�����y�)C�3mK��>E�����>�`C��'�(���=����h'}&�Tc��O7�]�F\�?,5/���.xi���"�D�:��m���uT����$�z�+���)����oS#o��1��h�x\���"�=�̜�d����;*����5?I&IW-]���|�e�B[A+i��Mz� ��&���l��+���n�N2���O�x;Wi���k��9s�}��D@/����V�h\qc�L!����z���W1�(���*˗oLY�Fb�i���Bゲ<�G}W;�M+���R�[�Z�N�B���z�=�#��&���@ʳq�$������|�v����Fa���$M��i�ww��^r���x�ź�n���s �{�R^�.{M���I�h�D���?�Q��L+��A��r,�(N��y�
h�� ��h3�z�S���8+V��&mƪ��^Mwfl�~�g�W>&�&���!��y�#-nBC��������D��#��ko�ԂK���!�~�f�s�r���b�7�^�4QVb��,x-o:B(C0�~�����P�z������#���bA 2�?矨s��Ѽ�譹>5�cy况���)Qs1~�=��\u�Ǎ!��;b{��Q 2W���A�[<��z�!{Bk���1�d.R�*-��C�j泴���߃����u�T�r��A��_0�Y�[�	�Q�B��T��+����
�Y�"��J���|��