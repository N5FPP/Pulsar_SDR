��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�����"WYj����i� �N�7A!�@<e�]ң�;��5D�監p�.� ^+��Rk0;Õ\z�7PF���p�e��	��j�kdD/���1M���(���T�e+qr)zD���FWkV��������\���mk�*
`�R���	j�' �� m�cD���9:�DhT]�����۶�����i����ޙ%��d7ܷ��	�:���U��(�����#���wv�pFc�o�m?���<�δ�7P����( ��(�����1���o.O����BE�l�pSX�m����
'j�ߑ?�a\����3!���Dꁖ�0������zܨ3�")s3G��>em�~������X��5��������h��&J\�%Q��JvB�YJf,k���k[`u�&�#N���Z%���[�+LP Y���c�I���qt�U|a�e�@�Ȝ�J�J9��1G?&��Q�}��ۊ"I��f� ��h�A�P�T� 6q>�Յ��? #��<-�Rx�L���?e�����Ǚq���M�V���ܸb�Ӏq̗,�'��B�v"�g����;��'Kf�ɴ�$E�*@�?Cp\���<�	�U�I���@�X§!�Ċ/?C�j�ҿ��ҁ�Q�*
�j��Ԟ[�Wlh�.t�%�0�ue�Ӭ���[8�>Y�#�݃-!ET����]8y�&lD`N{�D4�g4v���.G)��ՖJ��3��R�!r&�Ful�C����Ɍ&����Xhd�Q�ܾ��Uo��I��l�F+����٢4�%��Z���t�܋��2�>�V�>י���74�K��T8h9>n0�5���I�tȾV�Z̔�'Z+�[t�D��|y�L���v�w�/��Q�ѩ?GL�G��.�{��M�Z��ޒ�,\����{_|�L�~z�R��ڗ���2<�
��m�	��šN@�d~ִ?Ƌ��AѧgN x�����(sx]��E���V�}p���Ϋ�����?��.+��A�u���-o��E��}��W����C�2�c�)CZ5�iQ��Ҝ\sI� M�?@[�[����o��-���9_j���򌔐�� ����z$(�|����ֆD�,2�)���
YOp�=m�_Xy��o���؉�1���U]@������*���D'�S�T��J��N�X,"�%�HvdG?<�/vX�ַ�l�sj�g�� uo�-�v�Ȕ2Jw�<x�Q�qoC[ˡ���\܎I���?g�͗q��X҄6�O�g ��k��]�֌\͕�kq�c���C�%RM��4��h�����/2'<�Z���}>���h���^���_"�hC�[f�����z��<N��W����-C;��1y|1o�"b�;:O�ùҢI6����'\�2�'6�h>�^k�`���-)a=�T>��G�p.H�'�
�P-�����+0#ۼ��`�u�ǈ��	�|������W��P�5����A�D^�Ʊ�gի�ib��s}�G�B=�F��<���V��1!�W�yn���G[N!�9��;_L��_b5�5K�'&�pn�Y�3p�.��65�.y �GJ H�v _cʃ��ȷ��3�Y!f�l�r	@*������:R��l������B���Q-�e�Ч9s�TT�6�QZ�S�����������:>�+�w�7XmS��I�5@�h��VK�����k��E��)B�(woG�!a+�ׄ}�x�NnT�v��l��ˇH�[4�!'��3?~b�� 9� ���g`.SB��"'A�I	fM��y�� WW-��ז��kB��E���}J���!��ׯ|���� �5�-n��0@�x���ٺ��c��z�+~��[�l�d��%�A�9�"�S�(U\U4�mY�_
�NG���p��1z�����6C�����<D�c�҉��}��mt�Sꘊ���[KvŗD4 ���)��z�/{�~�7 ��ޑ����*�_��N;$CC4��e-�.R�Pʵ��8�%�a��ͧ�Z�[o!��7�Lүw��?,˲�¨b����(ߠ�m2��Pl��jN;����3��h&�f���=�Y2�j_�J���!��~�wi��:p��)��S���
��
�b��׽S��@�˃gBL6U)C%�-s��O���I���܃�a�S��������}25�cyM���\��#�=��,FU���W�I&��g��v�5�}��t�95����ͧ6�11� h<<��f�N�eD[C�m��X��2q�*.�f5�_?@�D4�E���ω�ד������{�ߧ���E%�طc��/�4[���mj4\z�9����n�z_����h7B��|�9$�yTi�<�e���-xe�K!0du�i'�c<۰9��v<ƀI/wN>jemˣ��31�/��Og��t~�r{��/E�,�I2�w�M�F��9wsˢ����\�����$����� ަ���t�j�R�_Qw
;�X��Mٚ��D�WH�x�����1֣Ȭd�K��^O4$���uA�#��9�,g^+�D��hd�~5�'��0ύ�g��a��0���Y^Ⱥ5�{D
v�gD���4���dS-�L�Hw���6�;:O�\�J	*Dc��zԚX�<���G���u���D9+8�s�`FV��B�!���0z�-
Ȧ�&��_;"͐M�&9����6n�����s���3�ƀ��2=G��O�KoŜ'M����aز ��^�c��m�7M���h�1ƏV`}!��Ih
[*��88x�@����0��|�Ok>�c �� Z�8;�?�I��O��y@L�ߐ�h�D������t��\�;�&N�/�4�ڑW�[^tf-B�xw�я����I��C�;�򧸐o�F'����Btξb�ޯD=�G�@4�)��B[O����'�$�:Μ.c�� %r����"zN����a�9��1t�o�ء���t9E��`�s,�}Ы(��9�0��`��W�M.�������
��}(�}��<��#pp]�D��?��%&�g�z��.M��ˋ�iV|7&Q��Nr!C��KcFv�[��<?YqxF�<"�4�0�y���wk4l��4��6Q�H�'��=]��ō��ʌq}W	���;S��C���>�X��FvA]OZ�F��^S�d��R��������"�#�t�E�E�)�����-��)���V�9��Up��������O�9[����-$uQQa���+��e�+�!��O�}mJU�e3c�T��B�_�P�Y��B���ٟ3֋�%BN��3��������mZJ�Iڑ(�Δ�~ĝ�A�)9?�����izYm�mf�6B����/��<n�'KK&Pq�3��$#�'�`f\�����Ր�?`昈!��H+GK�d�n���cTR�/��2f�K���L84�cd�� �����oJ�ŻR��lk�Eɧ)�e���n� ���gp%^)�ա1�t�M+�w�)�)�<�{�0M��ù�rTW�lЬ�/j�����Z6:X�B��T�s�q_Ylr�JmId�[eu�
^ta_/쿳�p�������Q%-�
�����`���8�G�0���L��Z�g��T3�s���eWyG��=���'øn�I3�>��9������h��`���V䫢�B�E�Fj��\pH��f�}�����
L��°��e��Sq{��5.�)G�:��X�#�A�T?���~��/@c'Ʀ��W��ޯ� 2|����)���A%�#Z��pq�I�Ge�E���o	8maV��t�p�~l�Ż�N$���:_�ꡅ�ɻ'�v�J��4��qD1��WN�GG���Z�,�0G��*���|�~��=��L s�ok
��d~���[�Uzb&�y����g-iB�ʔ�V��{<��6��S�����A\o4�A;+1�AǗ7n��>zM~B|���e�&-���m�� i���� ���A�r~�Qc�� �.Z@�Cdd؊r�I�Y<��x��Qʾ֌v����8u��l�^��T"����S����2���BN��&�L4  �����eq (�Jւ_��*k�%*;HE�%�xnU�i��L��f����F�>�.u����n������^T=�10^���E&:@_4cu4n��2�߼��3NS�R�)��@$��p��獮��|�
���B��ǜ����B^��.�V�՝�s��35���H�"��B>�����|N����/�ϹU�F�q{\�|y��BɎ#g�X��Y���=�)�B҄��^�e�@I�4W3����͸�!'�WN�`��K��)�W+5�n�L�~��~����Ħ�D������-n���H����k��xf�x��o+^�Nt>ө�^���K���S�ҼƷ?�Y�P�UgHoK�w۷3D邱R�w1��(�2��wN���IC#�J>�r��ڬ���_�kmnt�����_ >��E�)�7�h��	w�3��YX�>ڰ�G�4P�U��E��1�O��9�R����v^~�;.��eO��J#h��oD�F�̱&Q��W���V��(rd�\B�<m��?�g�!J�v�1���wg'a��V�ٯ-r�ן���"�ֹ���AS�cJ�}��Ϲ~��,�ڜ�g��].�K5i��wO#�����r�
Fkg��SKSX�E��F1Pd�X�o/i /9�domM�cஅs<��=I�%{�0c���l�}��N�_�O٬Y`��p���G���ϔ M��j̔��ʳ��{���՞����O���|z��a0�*wz�g�A]1�n\��U���e~�&
xi�x�$t!���w�&���?���7I����
X�����X#�Lѧ�*d�+�]F	�dHHrb�熦�D�$G �G��iZ٨�f��g=�9�}«�˿�չR�����.^��G-h�u��D�3 c�	��~�+��Xz:��7�ۘ�U%�gP���_Ⱥ�W�����iEa[PRb톚S��l.���?p#�J�ܔ�4�ui�4�=Vfa���L&�`���EvhuK���*qQ�Y����ȴ��1�+RO��9�	W"��.�ECF=��E�3���`�ek
��
��,*3�'�K�!���˱����c%����h����2֜J�-�Td�c����nׅ,I #4Dh�ZG��&�)�z�L#�(�5��:t��P��P�2��"A{�ȤL�}����b�&���r�PK��ʂ�)�^g�l�}�T��O}BǡfE��ٶR���h�Z�@�{�<�g�ܼ[)N��«�C=�
4:�^V�!��.B?etx�yI\g*�I�6���F��3��ah�㉫���9|�.�H���B�A`/QB��#�T�%>���M�Y`��+yj�xF^���l;�~��,#��x��w��m�\�����ػ�P7m*��Y���O�B'�(2k���̹�Cߢ6Xd��vE
���+�F��W���Z�����!&qړj֪љ��P� �I�Z#���3�w������ ��'�,�i|+g�3�E���ͥ���1�Is�����⟂�Z9Y#�|U��S�6Y�V6�����*�\ CA�ɜ�<�11ٞh�v�4+��,�����	�>PN�9��1nE��+p3��KA:2���I�|��̱����C�KD���|U���E"RN�?Ġ|�ťg�s��i��'�|����"�h�����*��T���u�@�P��C��yL��M���'��OG+���o��A�1�-?�W]�D�ֈ2!�Y������υ}W�~-_(!P`��W�v��V2~4_a�Ǌ2�,P�j���:}�t��%ĺ�I���y7w%������i��S�T����?���Yu*`�a�(�-��P�D��҂<G���Q���m`x��t��q�Z~�'.>�� ���#��-�?�.cQΐ�V	��r�M=�5S7 ����>N݀J�zr]_ ����d����[���P�W�{A��?t�̱�¤��C8l�V�R5�ӜB���^��.����P6@�8�N�^e��s�`ʯb��h*��2.�3b��C��VE:F�[=e������5e%���ӏV>$d�����x�<rX�-H+���E��i�A�X=�˶�Jǚ�E8���Gt�Z�1���MZU�nl]�7h2�ϓ�J��X�hl*�m��>�,u��f�Q~�!��oH�%o�[#'}�{dp��P��S���L����<k�L}���#�i�m3?�o�g[û���ZOO�&�G�^5���FP�b@�Ӱ�m�C��-�w�H;h̻��i�md�wPZK�W���UGN?�Yh�׎1��m=#U��K]|��D��Z�Ll��?_'��aa��4U�T�v[D��%K�ɰ�(��6��]��I O�g�
���թ˞9]��E"c@��1F��Y��5n�<>�>y�%��N>�ҵޏB^���s���r���r�b��H����zΟ�%�O�>ʜG��P��/n��.���ڈ�;����=ӭ}�H.��|�#���j�t���næ�`e�dKu�A2R���gu)�Qet
�]tV
5�
�Z���;S�Cm?��c�$�֕����R�	�Ya�c�U�1c��"[�Yh��J�����y��.���,�TM���	Ƿ�,ȣ��F���K�wr�-������;9m�jN}�M5)��+*CPq�����$���Z��*����qOa~��P���o  ���4D�M��LYUeb-��5<�wS|��աA�g԰��vrF,A1����
����>��U'�iRu�|B���[Q��yʳ�S8��E��.V�̞�Q�L��z���Q�Oj��������m������e�����	����d����_Ȱ���oI��dk�|������@I�w���Z�J�i�p�hp�f]�uȐS�=�Q��ͽ��e����
̆������+/��]餡�����9��Y,�^��w��օ'�M*����2����蔫>^�N�A���%=t�3�1����r���&ʟP;�ʐ,�jK9�<���ޖ�"�Ȥ�
���aolM8pF�?�p�R��\�z��=�( &䑷���hbC�[�<k\�W�V����n�.~��Æ,W,2�>��
MZ�3,R��:�}-�n?"&[�+�.a�8Ñ�<:q��ݭ-[��L������g	� �C���/�@I�"�=�\�$��x��wVu�ᗵ�Q��hC[�e+��3�?5cd��N�a�g�	D6�޻_�{�gs򳹻{B��G9�h���sE�3 �V��	�Yw]w�C�5�vqHAAI�	`wr؏���Ł�ˢ%����s{ťa���d~�m{nK�(�4����׾�I��C�H4���4
,�o^3E�r@�c���5͌S-�;)e��8��~z՛�\�o>ɔ�a�?��4l?����$���S�{�74���{����Q�
h��Y�Cƪ.Ì�p>0�Um�RR&���K�-I4��v����t��^&����̯����Vܝ���D���(�w�4�@O$JF�!��9T���Y ���A1�n�?���;E0��/��lP�z3ͥ�7ww�s�_3��&�&a�Y+2VIw�TL�ؼ����Ăѓ��D\_dORq��:��~u1�B���
Xo���D�ؓ��'�7}�� ��jB�K0x��B���2\c+��$Ę�]�6�s3E�"3& �(yLK�t��ISL��)q>����p��]#���3�*�z]6zJ�H��ņ^�o�p�����or�*���OZ �	`�L����}��ڈzv��[�˄����I��΂ʶms��C���%ݪy��,�'×3�&ȿ���;f�Y�%+b�����B�䬜�2X��KU;��OT�\|���{I�֨`̝�l|3s���E���ə_�<�������h�I�~��|��x�MACF��X�d�N+)������C}��>#�[w_ #V�SI���+4U�h�3kGd�D��B���-��u6��IB�'Ve�%��W��+�����W��Nq�Ѕ�����]Y�w�	j���A���Ǜ�\��_|�x,o\̔�!��Q�����t��u����F��X��@I� ę�����W%���Ne�d9<I��D�kc�j��BG�x���=)�f�t3mݾH���hn��;�q�;B�}:j6��Z3����a���~�Df|��Cp�5-���D.:����A�/9�-L�HQ�C���U�E]���:^WXj�����~�:�M6�W��$9'��5|���@H�%A��[)�
��9�G���o���/.��]��y"���Xګ*�����Q�}H��|YA�{�n� �iU���%N�����b�l�_��0��\�,@� vp��&�,�����A_)��C<�u]��)�Zo���ӣ�;���bJ�h�����ꥩ�)A (x�G `�q�Y�$��?9o���g�4��UOC�1�ކ@\�FHzsSL�����E��U���_�V��+�V{�[B_���� n��p�p��<��Z,Q���ts�,�f��KA��Z����<�Z�we.>@��Z��ȺW�Q`�k)^v�a�w!�v;�1]�.�1�q���0��ݥ�VҘr@ 9L��I�z��֩ƮL:���s��bS�ab�R (:� �ՙ=o�y��F=
��9_38�7�k�3/�� �����{1k�Ą�"I)w H�z��ږR� �L�&��@_�N�w=��t����rƙ���h�g=Z�7�wZ-.YƂ}��������Z̡��x�+��C�k�g��o�g6HL��tɥ"�H����.�M7�hdiOE�5붧69�U/)���v̝��m�'�+y���X�����ޣ�.�{l�@{��LA�͑��н!�l���e�#���9f��Z���W�O*o5���P�@1,!99�|����2�DC�TM��"�d���bإ5u�+�l�#�ۓ�y�G$Q��q,�l}nM.����4i+�G�{��H��o�g���~���C�P��L����źH����~9`�ꉄ���Ӥ}QMws��Nx��QR��[�����a�@\.J�F4S&0��(��>Z�b]��U��N@�Y���
�C^�W�6	�nXv�.��ρ%�^�Bg]=��۪l�� (HK�(���(�%�V&���n�:H;�i+H�H���0��Ui��E|GAؙ g��Id(����)սrG����x/��J���@rჲ�$Z��D���t�`3�*J}>,�~
UNL��r~����<�R�ܫ�������耉�;����?�+�\4O>л:Om��]..�u�0ז�p�z��RmBP�RJD�<��H�"�"�rzo��t��\�4�I';����7��Y��_�����ʓ:4�dJn�V����_@�������E��`#�,�[a#&h`2�S��2	ݸ���-GR�T�E�����=�QS�QY�p��/nIT��t:����mp?����i��>�e�ؔ[m�����Y�)��w�e�a�=$c3͐���Py1��@�B��� ��S:O���r���`ׇe%��"����o$ӷ
�6	?ҳ)�n7��Q��If�R66٤�plp��p�2��	:�Tf��O�@�%{���l9��+g܃<�J���=WjE��t7���zҍ\�/ם�s�/S�6eВ����r�ٌ=�8	L�37�a��HΡc��Ss�~"G�o���>J����O�����9�"8�)+u��B��T�'�ʶ�z�5H	��?���^���v�ʣAQL[
�����'1n�܃Ř�)�5N��m� gt��+�&�I��ŏ��!Z�u��%�B}�����Bꢦ<�X�W���)v/��T-���P|��uy�/�5uM}p��a"1�]ee��e@�V��Gr7�˝�ά�ؚ�8kI.h���+����P������Y�7}Cl�4�L���"�����DFAh*���p .�E��N�@��}̌��������[6h�;�h��O#9Y���]_0]:�"b��>$B�����G�R�#��)�n>؜$%�2�Ug3>װS��ԩ"7}�}m*8�ma斝�%���P4�1	i�"�v=�o56K�6�z���e����w��s�/E焕��?� �d��EH܄[fh�:U�
�����`Y�;�1��/WJ^��ᗂ?���y�bۙ�����A���),&���*���<h�/�?��k~��"�Z��p�__�Jo��Wb��e��5�(��4��Z�sC7�o�������\lQ��qG���m�/pC����j�'�K]O������=��6^y��&�I$[l��l?�Ւ� ��,刨X@��y*�YdV���R�ζ<).g������;�A7�gɇH�׆ PC
J�%X��;���<'�
E���2c�'c	{�xf�oN��q�!~ e|,�[�"`�'��@�U��73��ٻ
	N�nC�-��3����DBx�$�o�)1r�#6$�Y�@܉ �x�N���۪�}��B��@�)qԭyz\�
�L�T�T�I�c���QQy��0i�c�y4�ćk����]���e 1O�PDX���;�h�D��b���_���%��9�u��.}܎x�ru���mq�l?�2�c����^�5��]�/�9dU�m[�r�T�����w�d��t�Kk��1^yu�Tؑ�hM9b!�2;���y��ׯ����r���P�ƲI�&뿅�,�(+��w*T��?Р(4�ժ-�k�+uOФCh�رֹ��R{c.���֣`��tp��ԡ��{�тl%���|�P$���s\b�و�#��=����a	�_߹m�`s��|� 9�R�?*I��A�P�|Y�}�[r��R�=���<���_^ې/�L��lZ����;nub�W��3�-�!�/8��Z���,Xg����%��!��ϖ�K�8� iQ#ko�^�y:��c�eU���7�ƕ��� ���C����ޥ#!��:��S�����S�����?N�T+j���x�~<{��#��,ʿu(r���sVH��nV{S-�B"�{e� ���g�<�/���V�e�S	jM��Y��tY=���Py�����Z�6%Kę�v>�A+7+�yD���r���8�#�T��n�N�fD4���ׂ�-s�a��K?�W|E�=/�=�H�(��J	�a��)嚝�c�i�w��,yq�Rxj���a+=�o��$qۊ�0D`+�;KO���V�,%��@M=�?�Jۛ�I�%wP��2�y��饒��qt�I������>X ����sR���WU+-8c�؄����H�9q��5�5��r?���U�)���ݸ�??m��T���۬q�2q1�;��:�9��7����=zew�\�-	����
H�H�k��WG�w��r������!v�� �*[��ۅ}��+n*�׉�?ge3U��F�((����@�~�=�{z�[���y��YP��'��N-b]0�Ip�or2��I��/_�9�jQ�
#Uh�X�Ԏ�s���Q�rc��)w��pP�Y����j��
���D������a�fY��qY�U�L�	�D%L������m�rPp�X��h�"��,�S��Q�i�ʩ��ڷjn"p'�+�#�f� �&Ia"��tb���)M�k�Rɪ��Ԫ~oC�{ ��%4�<�'�l�� �B����qR� ����0�}�^]�݆�ct�쳸�§��=��d�>�T�Z@^���#����I����Ы骩�⨖¥�,m�p�>-�b3Ϊ�0���x*`(�,v�F�F1��>�V?ZM�c��oL[	\�� L���y��2L���]k[D���+m�+���&Y�~�g[�

���l'�S���;���R�;��ȥ�fٔ��ګ,G�D��p�����q8E+U	-W���
��g�<��n�R��U����4a�F�S��[�J�i��,��D����<p�m��5��Ƣ�k��H:�"X��!s�,W���x�͊�6�K�m�kM���lL�U�폟������������-aW7�g	�YX�>�ו����5��\�9�Hr���@�h�u�If��ڝoj�P��Û���������Bk:b��+>�g�r(�e�3;�hwuS�^T�_���yS1]��b�cI�b�lք�Ҍ��r�Է��4���\9u��|�pf���ؐ�i�ʫ��a�[=����P���<��3ԍe��y�&�?��a��H�%!w*U
1*�t�뵤r�~B���HV\�jm��w�R:w;��w�-��r�x0J�ۈ�
Ī����Cܒ��$��%A�O��X����d�����	���|����+s|��jZZ�ne�w�xɡ��G���gn ,F�^l�͖4 VU$����I�n���`X7�P��#�n�Nib �L��ˠ	�k�>��w(���1�C3�Ou�M����N�5��>�h:N]?�A��2[�c�vGK[⪝(��&PQV0!�	/_EWQ2/��?��_c�Da.���ݺ ����N���ᶋ�J�a��f>���ok��:��T�koA��U͞O7@��:o_vNZr/�ۖ�'�}X�p�ƾ�/�oP��"x�w�Z����/�Ih�]���1�*�(z!l~�{�q�0��@�RE9	�˔�Z�/��^��}}�4�Ȣ��T����i���[�F�E�V�J�(�[/s�8���x�׸�$���7=O�&/�j��2��@��tH���6ɐ*��������K�A��.��-d�y�YI���b����6K�lHY����X^-u�ˢ
jZ������T'n��·�#ys-��,p,"¤�|�]%^��v��RǪ���i�!������FD@b�~T:��p�:�, ��KR`Zb� aN`>�U.�j���Z2c5=����@Ԃk{};E]��z��P� 3�	�?]���r�C�٥r�*E��k	��I}Y��{[��`V�iY�6!׀ZY	��G.�*��C/J/�΀�ǟ��a=��(�u��9EӥX����w�4(c��ĢOv��R_^��-���2ĥ�t�<6,���~x�'MyJ��	��/����ܛ���L���t�(샃=ݽ�x~�{I;�\;ޯ�1X��jC �e4�vÏ0;�+N�!�{�yY�����˩���|g�C�族I�Z	�Qu?9 ������ǎɇ#m���1"lԀ+9���FT��31Z~CD+��������w�+B�Σ�YT��'��r�?n�ʁ�}�F�A�:�]w��DWQ"�"���D�D_+�u���B�Ku%f��� !*hw�r�:�:4�*����D��G��+\��E����?�3�!c��.�l�D�~o�Go$��T���&����6�ӝn�5�lZ�f�糜�&�;��8�Wg��鼞CM%V8����|�%W��[��3�zS%�3������Y��i�<�첦�k�3�W��n�z����-�v���%�'���> :j����#�1Z�X:{#�B�'K�ᐪ�F�/�FQ����בgm�o�󪍳ɮ���o���4���:D��s�P�b���
~'� ��Y�	w�d��̴��MBJ^6|?3}R}���]��n�P����oa�WQ4��sL<����O�&.��!eՆ���S��a��w�#��`�K�[~j���<}cs�(-���79��,R�EG��7�w���D��:���W���f��aA���τ���20�Խ+�z]��X��㬢~GA���~}od�� u��|���l=Pq���| �u�AA���w�ޜ��c�b`��N3)���,re��3["ݩ=�?)4��?�����U�����C��:���bI2�?�WHXL M�j���	�L9?�o#`s�yG`p?���19�����B}q��c�Aq�9��F^�7J�6x�ڲ�Y��_RK�)�h?����ͫ#�kx������������ȹ^`ꌖ�=�����t�Q_�?%����{rU�Vᘅ��
�k����;����̡����pA�L�Wc̋'Vҟ���K�d����9/�@;���Qz��L5�X��� ���E�����W���#�}�X�Os�tĢt���x§�>�S"�ҁU#-!Һ�>W$^c�J��X]H%��`�?o����k�c���x,�Ω��ʠŁOLA��e����bdxP%��R:���߱�ݔq����fכG������%RUX�јMR��������n ]����z���|1�x���۔i<��������=�s:w1��{�
w� �f>;�ѫ��ɮ(�e�)�~�{�u�x�x`�`KT������9ԃWq�e����p�^eՎ[R��'�I�k��<�	
"�����~z��'�qV&i�cV�87���װ�P�H����?��CM�9�VZo88��}l������8vl^�Ĭ����%��l��A�4�r;��~YDS�
8�����k���������ȶ7�s6���k��lZ��p�O.�+NJ?,�b]2�`��w}z�S�3�u�1{o��f=Ъ��3B�F�>8:�U4���MÕ��AY��ڟ���U*�Oy�-{,S��Y_��e�D�e���L5���R����ER>\�|�0t��1�$�OZ��S��Z��m�S��'���9z<a���y���~ħ�.9��J����C�����Yt���X�%B���w�3��g��`9������!�_��GrY�VN�$����)�KOa�n;�1\��N���N��A�64�K�.�a�����#z�m� @y|����IO+��)��d����4f�{6��� 3}�sVv�ܡ
,�#W��g�_�3���_N'�3�Q+��C�>�&�Rnas:{CQ��=Nߚ��STW�^]�$.�s ���㏤����M�~!1ن��H���B]��஄,�.�����VΚ$��NM�ͨ�-gw@�J���jx6�3�"�D�к[Z��<W�nR�#�B~��4��@ct���84w#�!�m��9���u8>�$%/�v4� Y��_u4�86��Jb�+��ۤ�����
��9��O�2;Jɀƶ4�z����=�,S�tu�h~�5�b[�Шft������,8��t ��E}�Mw�8�<^t�)���O���=�M�)rEK�oʹk!?w��z�8V0�ΊӬ�\%�C-�-��ш��&�8!u��r�Cr-�
�1��dVWN�,�%G�?���j�-x���]��]j���t�腙a�QSf�@-n��*^5Jo���6��d8""J%��0�󯘼�w�B�v�����q+�M�A52k4�J�;��%���n���<���_�:X7] :"&l a5����)q?��魢Gb�u����[�k6g��ؚ�P**"d����,����/ɳ�͓X�V�]��O}$�6�W��6�4� ���c��m�/(����C���3�/�T�h�!8���Q�j�}��vf���4*���uFP�9�o�|g�0��L��z�;��i�_�vY�-�P������/bC�Mf�L8Q�D�������\�Ț�JC�W�nbI���p�G�t���5:Sa�s{u��ώpO!�}��\��a��\�]��X6\j��?��mqiP��\�¯I�yu&T�#H7(�>�,���c�M��#ê$C�3�`Ap������2����˗6,%BPp|��"�����O~�oЈ�f��Df��뒸�0)M�H��#�W�P���,�m�bz8a�ܦJ����gO�R PG��I-�?KŻ ����{�^o�" ˟eSKЏ�+����m
�-j�,pmJߋ��"�pʟ*M�~��	����I�o �?4�gq�� Q�����ce�b���1WyN�p[إnkǳ4��^�E�X���\�MI.��j�_��0з=>��a����5G	�A]��xU��Iag,�	�J+���
�J��2���vv� lf�)]:���]��̚wYU;\w촸�9K8��XgFjms&�\Im}��{n\eq����}�ĥwS��HWq`�KrYu����c���w��'"=��-o�-%�V�%W�pE4�Z�"�s�67�ڸ'jC[�]�GS��0��w�K6�{���y��>f,c6�ȅ�ϙ��\��3Xۻ�ާ^]��iq�5���XSE���˴M�}Z��&#z�����7ߓþN��3q���tz�=�eJ� �+~��MZ ��6��`pA�u5���)#�>���/�Oxr]��Seӆ5��'p�x �=�Vy&��Nɟ�^3��^�X�	�5a�88�/טJ�7�pT !��le�����{k��1|�4�Uw�{ w�͜�����b�P�	�)�^)��`&2�?��7�q $
�Y�g�9'w��xa��O�FbZ���7Z���V�Z�>�ɱO�n��>ݷ��^�k��_���݋A��>\>�/l��~���7]0�������(��������PR�BU^�f̧`zC���A�Ĕ�av�Z�vH+;t��� �-f�h�'�GSiȟ+}fWp�؂0�����-���7��}��b+KfZI��H6�?WmG+�$v�+�>E��}zϛV��`w�[�x�z�����5��b�!�Q�/L�s�Z����pF'��M>cE�z��U`<N_���\mG�����
�:�1��{a�R�Y���{�{��[���}�e&�s$�B��ׄ��]���6:+�u&���)�2�_^o�D^uI� �Ǣ!�3O��;㉩O��דLKN��+'3��$��H�uSWq�xx�gz"}D��ބx�0��/� ���q�z�Sfry��֜_I���u\����7�����L��ڗ�.���E`C��f���n󍳦���k���濢f;����oU�cUR�q��>��?��Or��� ��X�����C��P��A� ��O{���ձ�GP��;���%���j�?A����"ug.ޞa�Vb�5%�6X��L��XbM5qv;:�'�{Ԡ�pP�D;�NFK���I,�o��J]����j����cM�^����ۺ̳��AJ�4|����^ ױS�
Ke��Ox�<loa��Y�r��3������T�t�	T���G�9�fJ5u.���/ݧ�D�=l~�+u��}ď������cñC9�r��Zsv>�!�L�b���|̲R��?[��vy���ޛ���61�?43������>`J�]<V�*�@��/0��e_�t(_F&��8�<3�Z�yG��0��tf��,r�uƺE	C�����Y���a�&Q�]q��v �W�2�����-{��@��o&���C��3yYa����{��+�φ�d����-l�R@��-�C~/�?S���f� �y�U�FmMS�i|��y�Hg16'�H�Uu�������j�����IKj�\YG��b\E�|��ඳ�q���d���fp,Q]��5�do#�J��]�����2�q�g�_�R��B}��;������_�+���zu	�r&R��HQi��0�g��Fӯ���=�� y-tO���r"�e���64���ܯ�G��q�pn�P�TXӾ$�~�1�~T=�����P ˢ�U��p����˴��f�\�6`���;��k�Ȅ����6}�<nJB�����Oim���;.סԭ�6������y��r捉e��B��~b]�@�C��c�T���+pw4|�z��hs�������z=GI��9i�h4b9u�G��ܴS�� ���ǡ�G���pz.���D�+�S�����[#�F.��|�O��7�(��	g m��Y#��ɝ��oQ�����o+�5p93JPΚ�����/�2�K���丩�/��`���!A�I�|˖Kb�3�\S��n�z Ǝ*�R�
�G��m�A<� �^>������vbk�TY�|���G�x�,$O����'���
�]�p��`�p~���a9�K͏NQ>( �t�~��e�&K�?=O�w�$�U�֍r�j"��\g���j~�}?���6*W;� I��@�|J)�,��_�^/���!�<��M~�yH~���_.���u�K��|�$�ړb����\�9U3���A��̯�>)B�zgE��nܭ4�� h�E��&��y�-���
lm� ���ށt�p|a_��ɤeD�3Ѣ�>���:5/[5�)h���[��q�?nCd�s�'[W���J�b�3�H�ơ�!�0!�Q.W�7sN}�ܜ5U��"-;��:��� 8�o��/�#���x�W����NQ�Uv��j3��ƌIF��'�eTW{�dA�
�7�8z����1n=^�v=p.�4�^�\�J���&�Z��M���nlݺ�	���Ћߌ'b��&���=@A�$f}����e�s���g?�CC�2X/�w.�&��M������n7D�Tm��V��n:Ǭ�o1�~� �����e�:W8���H4��������fe;�^�k��yC�|��z�_�9����$��pbw�<:E@%�	ZB��f���]��� k�!Ek�{k�R>HN=L;��߱S���&.ڴm�>d�ì|~%)P��T���/@��
;���JA��˺����~j;�{��
�Ft���G��.�D��)��r�9���R����������s����մ;��`1�qE�
X��	���ش�A7�:�x�)�Ι��G��$:��^�ie�c�0`ub�~��kJ�GWW5����'�\dc�ŗ?�׾U�{�
<��R5�\��w]��A,gF�J���m���E\H��2����oy���0��CФ��dg�e	E
kw������s0�T |>Q�<��@{�M�>q�������ɵPs+�p��.��n>XY��5.Gˀ����x(6w���`d,&F��,u�� �bh�v"k�4I���}E#�(��}$���'Ʊ ����{u���)�Þ���5.)Q��A�Ks1.d���`ft;'�i�[���'�"�,�ԌJOe�L��?�P&֧���2�t�ŉ��RI����-�`kŗ;�9u��c����"�8)����6D`���^�@d��Ni�ܸ�Ky&cw�mK���0TǮ!w���QI��e����Fiֈ�S�+��g`	_��L�!?�����7����O8%ђ��� 	����8�[���	�W2�B-��uhR,�|�,e���=��%\%#Ԧ���EÔ��KP4U�!��u�ZW��Y�G�e�O�!�8�j/m�8"����-��"��3/�V}����I p#���OW�S���y.JՀ�~�S��1*�5(�\_��|�*�������\����OQf����?cd-�C$����6�ƽ3"PCC�Jo�dy�L��uw���+*ns4�'OWd�O�˟��<��է$00?ޜK��c��훵e�Z��:�]+3�=@�UN`�J �H�cHIV*{���B-�"��u��	�Ƿc����+Ԑ�-��*��D��#\ �a���C��zFW�X|>R2��
_e�JQ�F������>6Deӣ�g5B���jf(�C����sCѹ�9t��>�e�����r�0S��N%1��Po�8�m��tu�u�u�T����Z��SH]3�@O���a,*�o�-@L� �(�FQ���)9-{����h7��$*#��M���N�ĉ��^��^�A��0���n��yUjSDC.q��$��y�̺y��=�!�ɣ�|��d��Yy�;F��.�⥨�Z;E�$��S���u�Eu�ر����3DS��K�K:1ؕ1�_ia���s��2����kB+�輿�0�Ǽ�A�*x�)��B!@ϣ��ӑ��!ۣ�R�0�'"^\��.;�6׹���Kco�$"{-b����nc�9��_�����VD�CO��o�hN[Ռ�ș��A��S%�=��RV��²�z���e��ĉ��p`��]��|��)@\iq�v�А��eмM���>��5��D&�G��3��GG��Q�wS̫��&u����o�I~�I.�C����}Cc�`�n�h�?�y| �z�=�3��U#h���
8��sc{�$صk�Tg��qz�G�7٥Bsp"Ipй/��������	�)���?շ�}h��	�ޚ�l �ya��8�}�	c�Π������Ǥ��H�uz�2P;a�flj�$�q�2]\�&H��@�(b������
7�?k�����_$����"�N��i�����Ç���dJ����v�
�8����:�����J���+���x�o���ͮ*\��xީ�������s*{y�q���T�iȔ���F�������x���7_���j�C5���lo?~��Ra����LE�.'�n�a��|���m�&|`p�+��!��C��K��4Ʊ�-J#qY?92l8����G�v"%�*�m��zS��\b�?���BM�-R��d�e���z��6L�Rd�H���B9G;k�O�������1��e��PK3�v+ʬ�A��5��e
qz�O�d]�({�p������A�wW�S7`]1kڡ1��t�S���}���ȕ{[��n��[L��n ��r���)��#PTؿ?�	�υN�� JE�����P#k�y{Y'�Qs\%�{4�1X��@ŇzU6�����	�噌����TI]��I�]۝�VDG���L�]��ϕ������LJo-@ez�pW