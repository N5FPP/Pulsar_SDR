��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VYo�p���&� ���_TA�xg܇/�u�3 �^UL��ͻ�/C��M��mK�ˌ�q�cI���¢�T�}�u.MT(���PeCĸ�1���`�aJ�U��4
�:��x}PS�˨7@JA�6Z	�o&'+���ǝ��*zc��}�J�N_P�ݣ�<�,!&��oc�־fN\3@\�ώ!(�\y��g̀�x��&d�Y�+$�b(�B����$W[JޑN�~��o����,4[:�mozʅÁ�����PL���¼��UJY����(5{�)%ΔoEЗL��Ĺc�����AҀX�8*���(⟜w�L�S�@N���	q�'[��=��:���p�ÃvD�"A%>�ܙ
�v#�feķ����o���؊#���)���{�mF�쳻��vt
�������s�{���?�ҞQ&)��t�ZL�K������e���s|.hR��,� S�Z2.�9���B��%xa��޻��y�m�e���sjF�ч�|��Ǆ���Ȯ�����\��B8(8��Z�Suy���=�Ю(��C"<�Y9����`����f�����\��4�{]�l3=��۰�OFn�e��ql&�"_���ez!÷l���E�L~ෘu�<�c�DB��]n�͵qMD��ۑ�����m��<���y�2©�r�<�
�S�v})P��~�(�oH���p�������_�>�ƶc���cS:w4唻r��P�U�������PM�@-rӯ$���^�������R�L#�a��7� ���[�@������0��x��*4E�t%���5���5l��֓A���˒~��޻U��X���%��D+�S�����i�p�G�Qҕ&+9�������(��ˉ���v#��)^���|s8�$�|�?2�H��t!5w����g�S%?˟�KD�!�rz�
�H�=����JFMxo�Pq��`1�QcNc�@�W�;�ci���z�\�J-٤;�99͚��r�ç�F�p�nҗ����S@���mA��� ��0$l�X�W�����?߼^(K���pFq�)�`���U�CB�y�O.��8v�P�c�(���V�S���\I��hie��j��g Hϲ�����GB4�5S%�1k��xd������N��ڄ���^O3�j>p_q���&(4�l4����z�e}�(��5DV��]����#QÎ͡_�n��,����W����^G��pE�[�������$�ov�S�!���%��k��P�ׇ�L�ܤ��ZP�ww��S�:V��N��w����%|�V&�`�nŭBcw��a�d.zB���|*3rnd8b�,�c��%�Fo}N�E6J�f�fԱB
(v��.��B^U��=�{���ng�#�"�)�g����)�R�3�2�w�i�'�.wM�*ϟp#W>�&Q>B��ϿfW���c<�z:�G�51
و��� [NKE����/����l��f/߅��F�R6��J�c��x(�}��/?��Ќ\]�!�	z /���L�|���^���e�SݥB��ESN+���� �P�yn�����Oo�c��ٕ�\�
���-��aܷW0�����S,x؈�A?�3��o .9��' �љ��|�?:N��DA��)p:��ʗv�^��nM� m�1��IGOrb���E���@[FQh����q'�/5�C�2��pw���knе�t9�/�B�I�E���=���9�6� �ŗ����Y�Y
�ph�0��C.ڞ�>��Ͷ�K�#�1y*�R�ƛ^��1�uS��_���s�p~���_�f��?TJ��|���������=�L��YC\_J��W@��2T�7��N�N�f~�A�9)6���R�M�aD:F�Ȃ�j��=��ih�$����*f.R�	����e�-`��\�헼.����6T�����I��)wЋ�%[��Sn��%���V0��FW�CI�^BR'9'T0���V�f��4c
�����'�4��</A��a��,N��o�z�;���Dc`0R`��U{�wXa6���qDA���1{��C����Z$��y�tq���(��H8x̄��'�$ۃԻ�˴/U��w�E5Ѷ]�w�#�E���wwqmH,�y�pS�]Y���N�MT�>��8co�`M�]�)%y����;��$ ��p̺��22�9��v)�T)]�{9��ƃ{�`ni�3:�Is�� )K�Cu։	+i��=+�h7�f'~2K6���U���u�=�I����?6OI%^R����ev�:���7���M�w�C�|��/��N!��k���r���QMx,���^/�J��cMKdW]j�$r�D;��K���&D9-�*�:1~�Q)�/^��	����O��_�D>I<P�oc8���m]����ӥ�I���D5���K�M����ך�҅�� ��>Q��l�y�~D��nw�h4/&������'��(e�.U=�Sz��,b�0wm���k%Y͆���=`�3O�Wp��}+z�]A��l�����<;���4��~ c�8�������;�M���/���q';�/��ȯ�G;���jhS;`��!e���5D��Z�΃nj��5~��Lr�-�6�I����>��2��e,(�c����߯�V��8^��D8胑�>����Md@6��2�%�9�HI+_,�@]p،+=6�^`���I�`��	4���t��]�'n6bC�^N�.RЦ>8 ����$���R�n(��� �e��I��Y*7�6��Wa0�� M�G>ML�r�N�\\�X!`��i�T�#Az|F��0ΡM���Ȗ�dB�.I��~�WR��:�/�U#�>�*���[S���2�d~M`Ŭ1i8�Y���*\PxėB�C��f4O��]:��*�0J� o���Ԡ���s�U�&Q�)���7e��FU�@?��0]B�pH0w�g����mQ��-*��=���_�N��@�V�r+��,�!AF�A*=�g��S�A�����G���d��z�FO��j "����(��̋ڱ.����ػ�]� B� &ZP�JR�m>�9��$���x}U�U�����g9b{��WrG"�"�/}�lE1�I.�\�#D���F�������p�5�~ד}����+O��CnW3�6�����֐mJ����OU�v,���w	��1�!�P �-�ym/z���׳)�o�&���!��U�eW��� �\�[�]��G�}�@�ls�:�����W�Nۂ�vμ�J�h.pD�![d-!����$���_52�0���W��x^m�b�t�
C�����daM{|N Θ�߯�떒�ϋ�8s��y�>Z3:��i � ���5�B�ŗ��ʟ��Z����΀+U�-�N =��g��T-k~k�W]GI�(�ڲ�V�vvw��?�����Ꮴi?���ꮂ=f�b�� �"��w�q�`��}�l'�e�z�p3�1�!? w�����R���)6�:l3<�ѧ��*����b/�o�o ���hU���!���1+�Q��+y)���=���@�D��R�����VD��T*�(��n��L�tA~�$pGi�ߠ+©\�_o4N�h�1���)�sN��ww��O&��1>�O�9��P��,�DF��6�b������l9��C5�\������_\t"p����z���V�>Z�ߎ��s���U�K��v�����8�a3�F��˂����Ѝ�I�"jYK��Z���J1#���zH�� -��+G;���H�R|�!W�n(?2������6����$0��� �G#ĥQB �%ܩz���N�n�n���b��vOz�IY�Y\���҃�n�Ӿp�K];Z�j��[>����B{����ԫ2s�(�0STB� j����`�T:�w�-���U�ݢ;���W�ef�\D���\VET�Z�;�u�F,/��OYX�h7��`CȅC>����<�t%2Ē��Q��QX^���Mb�z>�����sHo<�@Y�M ;bP�����_򓞵����Z2jg#n@�T��d�ӗ
��.���wMꇂ����D+E��Ϫ/��Փը��[{��71(�v0I��	��S(��f��O�5ҍ?�.$�%���2C��,s�t�ؒ�	�� ��U��σWMӓ(�5��0�
�EW�l���5��7�=�}գY2����U1g�߉����Ɉ�5���*oL0�͹�i�d5�F�mx�_� 1��U�+CQ�o�J���m�#*��,ȩq�B��81�����f*"=�hxF1V����N�"sa���w�*�r��v�z>g��W"��N�1uA�f|V �82js��U��Bl�TŒX7����b���M�U�g�dGFp�Ѧ�#��ю�����\�J@�\��qrCW=��,%/��@򚚛ì�7d���Ge���4��}���dPҩ}z��wR#���p�ye�PܗQ�Op;Ǐf0Dt��+�v�z��#��
{RO��,�*
/]䫢��T'�Ȏ�M�H��?_ېg1eF�L�|,x�l
�dq�wI
*|m~��ꚍ"��
�{V�d����g�D�B�������3Zě�/S�*LK�bI�F,�^���S? :�������N�s��j^7��X�k06�&n�/9R��Y��T
�q�l�S��-���e��7�ȱ�]��_A�75u��K��=�_���W���{_�L�Qa!ٗ�W�������bVG����cH�w�2����A�`9�[��?���uIƠ�M8��4�U���ѻ-MбR#���pm	��uα�A���G�
�0�Qz�2Ϳ�ےW�����>k�U��/��� P�p�6�W�Yؙ3�q�kh�T�[�fQ��⯽Ҝ.�-��v��z����~�c=t
mL1P�S�9N>�Z���(���bvw���?��׊F@^ �}��	��K�ws�[���B��-|�DZ�y�7����+����>#�B�*ϰ��~&�KH�-��,�r�û��-���KҠs7oRz�oM\�������ah� F�\l�Y����h6摚�叒��������4����d ߯�ZHեq@�B��LڶG��+�}�Ov�&-{�1�Um��"$�@��V��j�:���ɾU���Ě�\�2k�u����(~�[h���=id`^��d'�h���zELi�p�f�d�w�zO�Z�0!n����~
�H����f��P7�1|�n���,�MO�(��f)��|8��x,P{�K,��)����@�1�]iX�T�#k�Z,^N�5NY��8e�X鶂R t�mw�B����LKc���vW��i���	Om.� �+�>�$��W�j_��"�B�^�К�l�r��J��UM�)�D�J���$C��U�rp�M�z֧~���?E��O��=٩ƅe�*%�2��-=��'�n��dL��+�@�&|6]�ۢ�a{_?k�E��.�~�<�T�����������L 2����7�=�l�l�`�;4�����#�rJ���;�Q�BB���!9���ݚ/؊�&�*� gM��"g��W�}�b/�k�m��(ğ�W�^��:tO Ǭ��ڡ����{�&\Es0����/��\�=�,�f ��
����k`:�h�<_�7��(�`4�j�7�}B1��6mh��^�xg���&Vo�C��RI��~�����L���o���Qk���@�� ܦ�����-p��rK�DK��l�޷/؇v��^1?z����h&�e�ZۿA�^��ڼ�u�o�%<���w �[<��qk�a{8��wʩ�INK<W�tc��e+�Ꙛ	<���	K1��J�O�C[_����p:U��/L+�4�6~�|S���1�[�j�U��G���{���:���1�?�O�
������W����]19t�p[��W���$��
�?q!`��i��,h���M2PpuP�xxx'�ZÏU�('�]��{�8hY�3?�ۗ��+KTQDJ���@5�{���ƭu�7)̢�Ү:�+���i�����m�����.^����ٙ�{=P���1�p��,�`�)�=�=�Pu�{��e�(X��A=�#��&�8�����(1/��uLM
��QXn�o�A���G���S<p	}$�R.fst�9jcK����˨�N��̎?���q�4���9�%hl9��:P0���U�:���!ִO�,��(�|�\�9؈��Xi��?{�IY��a��[c�I�'\��������N��D|�𿮆�JC�Q�7��u��`�guI���{���O���|%�P$}X�o�W`���ҏ�
_������%�+RO_A�(�2��P1s�e�F���>������ ²T?﬙��4-��;�pcn�$\�ysJ��t��ʕ�l5�ت0�%�ݱm�N
��l��#����]�M������%��'�Z}=��q��U?�Bu�`$��
��gVK�j��t?֮��E��m��f�+#�{�E����������\�����lۀ���\��jR�	�����6�1GxB �'Q�N'���*��x���ԔHh"��Yxn�A�Z�m�-P-��,����1�^:�s�f�>9�.a#
��ß����/��9��Sܬ�ʯ�����d��.쩰S�:����m�ȑ���iN
)���q�hMEvSl]&����V;Ҁ���4�a^�1��	��k��An#�
	�	�TˎF�������@�8�\����ӼKV�|;���#�]��eY�^�ֹ�%d�y�!L
P��[�S<0r�-�7�^7>�u�E��\	yG������KȆ5������g#�O1.&��kN�u�3�����.,�0�{av=Ͳ_���!ײ��}j�e�O�!��X�S-M	mhS�%�����y330V��R�#~DAW���R2nZ���Y�֒�@1;�y@���j$@�+�gd��b���^�Q��Df�0l���[�ME{����o��ʌQ�L©���FF�r��L�w4���9�~=���ԫ��C��0�a�����b��K^OPu��N8���]���Q/x��%,F�R)2�au�+�neqT�=�1p�YDE�r�E��jR�2v�H��vΓ¦��8]�^g��4)r�Dp�Z��h����2�؜zZ�e �ۜ*�����v�L���U6�x�÷[���{�B�c���/%�J�,+�L�b���}#�����zw��>��a�<��)#+�������e� �'�I-�|�v��=�E��D�ݴ�e�s�����P<i���~���� J�:�I��hJ���e���IDaH�Г�&����^*#�ܫ���ה��I�/��&c��dZ5,X����Ɏ��Ye��R�ZD�zZo�f�����=�@��� }��Z��E-��c0�� 3�7*TI�5�xB�7���h�)s��k΃e>prʬ�u�nE�2��_'l�}�������=��Mc��d����]��p�;6�83��:��N�B�+#�2���yCS�Y��	P����*�.��p��� ��3 -������U�3ˁ��Y ����]s�w���|&Nɸ͈K!/v��2� �FU�VI�M�����6e+u�wKp�7��5W����G��5ǩш�ݥ����r��/\nS㌥U�P�ю�bgeIl���z49jG����s��Qp}}�t=��%��*�k�搑����M�E���QG��s�	�Bvj/냢�cC�@/�.��d���ѐ��g&A(�h-���G�F4�!a��P��Ak`%υ.̹����$(ZKgE�%^��l��,��^�}^�9��@iI�P������[[�Ǒ��������e!m�f���^��mR���7��1�1��e�J&5��$u�%�^������~���.L�#F�ٛ(��t+v���В�9zͪ�7��p�=*gi
Ag[��0k��8k$%F2��
��	s�t�1���GZĥsn>ӪH�n©}�gꓷ:��'xhD�ٙ���+f�9J�2ju ,����G�����y�hǳV��D�O�D'&��(�X_j渃��eV[��Ԧk��69K.$���Wd��`�H�%+	d���%���N�'�����
��G�d|�(�c�G��a堆�ND4N;7����i�@{q�ˀ`��VvVL��+�״���Է�p8�Ԙ���hw�8]]Ǚ�4nՉ����M�';_*���2i���:��h��"t�'\�.��Z���C����R��l���&?|Is�|x�N����K���+
�
�Zy��s���c�%���)u�Cj��(��9܉�h�g��Z�X�kPt8�{'���<�4}?N��cA:�V|�����	���9�0T/Ւ�ߧo�T��k]A}D'��؊�M��'�H,�m.Dǥ�b�rʺ���b�z>l��&��@0�k���Yf�c��N9bl!.w�21�֧ԭ��"��[+���/�8@��I�}���v�As&J����c�9��tLA��H��9�Bb���Ua�vrٕٙ����'����X�A�j�EC��R=�ǋg����zP(&��Ps�D��T^����=7\�|$H/�{��;�3�qEx�F%v2��Ĥ��S�_��$�@V4���Յ\�"�oΞ5�����و�H�M�y�q�rij�]��*.`�>2C����G:���������^�aO�T`u���$�!�Y���;�RGH��W�$���]_`�P�~�`���g�������~~i�;��7;f��&n���q�!�E)k7�o	��$D 7�j�G��x���[s~�m�d�����Ҩ����Ȣ����pa�(c�{$�_�uxf𒈒�s�-Z��n�P� =FN9�l&1u�m���.�$q���s7#�9r.�0s�(s�xS��LU7K�p�ډ���&m	.:
��a.�\�O�%�q+f�;˙͈a���U�� &�%u�g]`O�$?Ց�U�j��Z��F���´޳T
A>݋������K�_�O�.�G�1DEY_����p�|
���o0�^dA:)��l�_�P�Tk2Bm2����=g� �q��.�dXq�����ŵ�_u�HNƏ���CA� 鰪im�9	5i�_�Gr��,K�sh�貗F�O�H�Ja_�F�̨n����R{�Zn�/�3zܴ�f��H�9��Ս!�n�.�>1�S� 
k�)�+�uu�4���5����9����' ���S;�6�"��xW�5:�cs��c���+_�����Lx�%��6ٙ��3Бl��UZ�ս<�yO���RV��Z���VZ<YE՘������R�V�`-��[�����k���S:�(������:e��K�G$���ܭ��>6?��r��S�� "����y���f��A���C�����n�P/-�H��<�E���b������tq�:�oN���򁣍�%|�_&����:Ka�
��:��r�I��o�*�م���%���H�g� �ǿO�i�f9��>��Nѿ(�X�?|vF/\?�+��sF9��2�$�_Y+�c�z�Jٯ#�����x������#x4��K�h3^<>�
\	���kڱ�Kw��A��`�d��f�;F���6��T�&�η^����$��9��׵�s�u,��aZ"�ű�[Y�^���m��2ּ��Ã���� ���t=�	lͥ����+�2:���'N�9pt����� 0O��_����`�yQ����߬�}�AR�N�3��QȤt�z>yđ�#,2�I�6˕Ĝl�n�]!�=d��poV�g�.�+$̈0��3x�v��\�Z�ڃ�������FM���Q���C��4N�#g>���<����a�i��T�%)��� �� ��82� $��������1�#|Q?L��h���e��_�p�.ٮ#�0�+9{��(g����_Cӆ��<.�!c���K0h�O��	U�Ί�$��	F^v/����?q�#�6��r�3��y\#eb�ǹ%*jÐA�6|\�,�)��N��z��y�S������a�Y�(�Ҹ1������agڧ�,��*��x���N2н�L��2Ȏ�D�޼H+[V'Dod(&��GF��Q|�ed�f�=�,���~r(�*�
<�/�Z����]V�� �EƬ�ݤ	^�:�uu�egϲ�^�'��͚����jš�h��h���m��K���0�WޱPlZ��MF*�uTZF�+U& ��s2=��0x@"I#����6�b��9��d{t�[e.���� �,��ֹ�@���*�~���H-�_$�4���l?�T���l�ęz�:Q�g��CP̖�z2��#"�h�s}�X��L�7%�g�������ˏ"���+%Oh��z���b��b `�zv^���Sp1L�Q~0(�:�_`��@��eC�犬y�/��