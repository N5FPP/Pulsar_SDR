��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY9?�C�><�|0v΅^�V�2W�f�y2vD�&����~I ���Qw#��2�L�ϙ�K��M��t1p�$�-���ivA�����]�خ��MHn�]�Hi��<]�v�P�X��̝��	KT�`��~��ƭ�JY��R���W�d��s��r��5M���O�����#���I��+Z�"YSȷ�H!0�"����ƷC����{���V��;G&���������Y���^A%G�r�}t�����u�m��^������*�
�1�GeF���wD��3NN�+!�B���A����c	�Zӎ9)[8��4'j�b�f-�O2&t��?vg\�i?̯�ѡ�W�	��k�����Ǩe�[����A/����L�s��d�x�^�@�-�#����f�Z <A��y`��gŲ5"��ct���i'��ҏ"WÔ\o���'�ӐK9����������+��T�a�k� 0R�jm��~�ˈ���Sc`�p�r�w{���蜆� יʅ�� ۛ�3��2i,I�~��V�{*�����|�/�~�m�Ի�8x}�qK�dߊ�DI�������0/��@�r�e�Z���ᮁ��
\���I�K)��G
l<Rk��Pb<&�M�	�c�!���@�a��o��ѩ��F_�`��.:$�0+K�`;�K��e��]2z�ᬘ��w��&���YXd����xP�+_�x�^��L�ϲ�0�A�o�.k��@�d�h�G���߹��o~Dv0	��1�cK�뷝�� {`µrN������n�s獳�����D����j��R��f��VH���'6����4�]��i^�k�1J�a E�Ԍ����3��a��
su�/��v}W��4��Ő�e����\
�X-������]FJ*h7A����!���K>���Sf/��	����y���N�����u�)R,�4��
���}���O��eJC��2+����O��^_q��Q�uOg�{�	���9��j��'�����������T�Q��$&iɻ$K��x?{ώ��ql3�*�:V:��\�d�'����=�ʮo���R���h$��O4��R��W��r����P��JH�*m���ծ�_M?Zv6i�R�0�Qַ(n���x q��.��Zź6T��R_g��JW����Q���j�g�߲P�;)H1����g!.�����O,"�6�O�6�M����j/���}���L6;��톅��e��9�`����*�@��П��mD�$J���CP���UFm�o$��=�@	�j�ڽJ�N��=��L]�W�8�Pp�1e�+�w��'�1�H�)���u�^�&���=�J
�ɸcO�)��a��H���<Z�
<�f�7~}��cT�}d7�z�́�TSP6�u�.t�o�LH-3�m8��q��:fb{;�u�@�Įq�����(�d�pZ?���_hVv�#z��Ȁ��܏�C�f�����gr/TT4��'�?ىɋ��m��œYP�_�!�5;�W��D.�bL� H��