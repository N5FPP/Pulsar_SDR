��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjfm~���*��
��3c��N����-��REK�!���tո�Up`��H�րS�E��јj��f�G�8�u�h�����8�WD{���CAJc��k^�Zi�@�MR�q�+��.ɏ�D'{��7�s��ͼ�T�Cҩ+���<K rM#42���fHK7���
�l)R_�L�Y�e<�T�NsC����|b^�P���\�)z�M{�A�,��.cE&�}v`D6��5jiy�ϙݵL`�&'�V����w��n ����g���ߊ!U�"$���39�j����{:�d�iw�ɽ�Ձ���xL>���+	�(��C�x��O�����&5eJ}&��OH���}Ah���d����{ۇ���⟰4I�L I��V����y�`�12,���{FU0�L�����mU23�hLe�9��Wa�Qp�$W��~V#@��+0;�%U�ȷ	���ہ�����V�Q��c��v�ҽIƊ=;r}�C�tS�i�Bk�c4�+~ĚeEF�`�7�e�ޮ��*�3l� r�Lӕ�|�ôQ�������~�T�����p2 �"�v��/ �P�����ҭ`�?r�<i�=DJ��cQ�,A�F�s;�!���Y�Y����쉨S�
��Ӷ!��ܥOј�b�/Ҝ�,St��}�̓o������Cj@��WQu��UЕ��r��1"oR�)�yLb<�Nb깹���w�"�$8��$�d-�f��IBu2ж�:���|@�9핇ќ@�0j�۵̨Fg���{�o���c�F�S��M�`b{��'r�?�@�O��O��z����Bn�@�t�Uv�A2�@+	7k�Ĭ�$s)�wfiN'��B?�zlW���K��]XθaA���X,��|6��ӹV�}W�	^����@w���Yb^�]�[H�q�Q���eg�$ �4>�ZF��M�ٚ?Q��� SJ\7M���C ��[$-|C$7�D�t�Şd���di�\V�o���z<G��/��Ԡ���
Z�#A���U�V��w�܎̡�d�krCBnH5��8���ǝA���g_9W��8��w��Մb�M5uv[�\�>�RSA��w��f^N�'�0N�@Vczt�z�Eo;G���{�a?��0�T��PfQ[��5���a�7ƹZI/ȃ�����	hJtvF�5�\�]I��ęz�>U�Я�fI�u�ͨ�#�x�o�a�/%~�/M?f�l�������@t� �۾���|�.3S8��hj� �a��޲���,.B�x���Or(��(?rD�Ǵ�~=sI9����TęHv�!�A�/#S҅� k��? ����Q��W�M��8����������P���Ð7J�!a� ��\~�<����?�D�ē#�m���?�*uU���=E�,X�)K�V'?��K�R	Oޘ�;�C�V;;"��Odߌg�L�/��&1~<�!N0m�s�
M�v���s%S4ra�L�h���3c�a�&"&Z,r��"Ü��u��iC�pU�v[�v�cn��.q6C�s���#��P�g��F=���u��"�T(�DT��ƍ4߅�ң�Ę�ծ���U&�d�� �BW�*�~���ϲ���}ǆ������!�t�ORq���x0S&T��
�xqnT��ud(J���[��H�PF�5.�!��F�Һ�l�8>�u��,<e>���ʺ�d�����3�|!�q?(�C�垫��SW����D��M�Ern��1d��iF��R;J}�j�L�'����Ф��4ѭ㺍��,U��|�r�I�	�ɼ�y�+�2;��P�nk��+�:��_(��	�����k\����x�\W���tOyʝ8�b�}݌O���P�PG�Ƙǋ1.�����K˙�"���"�"N��b/���!rNH��y��T@T�������_6܎'���`���:CTt�Ih�D�
����mZS���:�dfp9�V^��u�:J���p�J/_�-�R���w���?%�{*��=Y�����N�8�ϰ3!ȧ��8���9Ǒ������^h���4M�J�>q$s�G�r:�f���׆�T��z��4�QW�G�ư�g��'� a&	����ѕU��_6w�v� g�m�����bH�!�� E����B4x��#�]�CM����=�l�A;Ѯ<\��E�w֭�D�͕EG�P1��/C����ԴLYz��NR�y]���!��q��{�����Oe�3���� K@t�P���nݡ݀�UՖ��Cc�8{@g�]�_�4��s-;��Aa�g�;�������[ _�e:�̝�H���,T���H�r�jGP������ PmBٟfQ��V��ꚼ5�9Ф��;�To�$�Y�,�)aĎE?)U)�SK�C��)#�>�AM⦏]�{vE*o:��5��૒��������펤Bm�t��hk�'.B������ȣq�e�&й���*k�G�Y.� �h�B��]t(M��'IT���8��Z���l��lڋi`�`��[���j{W2�>�m-�-_��a�#�6���)>�lCë���o:��	���g�E9y2ݣ>����Q��)0������)�3���+�2�x{l؅'�'2�A��o�)�����If�Zat�yǛ6�$��Kjc���.f���8�	h���;V�W:.���\.�{�n*K�&a��uF�B�k�Eo�!]k��H7�߽m��������ח��y��`rk*;�F$m��ɇ��x�����օ*�W�r�+�����TP�sc~KS$9���n��/_�b�]��P�nl��=�FBea=��3�����㌄�X\$��? ]�y2# ���6# �:��pl��SDE6b^}�0�.�Zw�����C�s�xW�q�S7�>�5��~0��.}�k�b ���s|u��c�xǃ�p��@�m!���7���} ��-FP;7Fu}1��%�*�����϶���:͂���`E��t"�rFd^��H�[|&^�\�bҾF���ac������i;,S:G��ri�[�j�]v9Se�����bs�v2J;�r��߬Z�W}w�Φ��5|��_4���2��p��KɊ��$g�E]Вq���E]�3Z�'3�|-)�/hY�,�!�n�sH�F�G�E�g�ϭn��݄�(D͑�g��)�(07��H̴�ġ!m�j7�!l�]�	�6H�)�Iqگ5�n���ڌ��&#.��f���:B¨��v 0
:��}�-s�VC��ZԂϯ��9f#��e��ϭ5t$����hf�A�#R5����9��:�z�m�O���{�L]f�b�Z�k,jQ���{9%�4�N��b�1�D�iy���I����[��X��5gF3;������G4���L��tE�n�Ir-������kE��`�>�mW���Z�D܌����:����?@>�{,	6G�{f�I�����: �/��P�>2ڝ/�����p�ϊ�Éd&0���>q��ӛO���FʳŶ]���D?u����<ZΑ�s8i$��Z�W�3\ݪ��d�I���'�-m�fn��ƪ�`[!	3̛�ΌΊM������\�D�h`t���S-��D88����2;�X�����K5�(��J�BwU�vL_� ��g�J�����6=ɺ6!�����5�킱��00���yI_z�]���f�\�@1�$��	u�4^�9�]�ڤHo�U\GOpAs��uY�I�t`�т;�>ķi��]������f���,~-��bS��=��,~�m��eg�
�/pT�ޚI)IO��þ�t�m��	i���|$y�9���ʍ%&��r)���ko\��7�G�@z�skL��CQ�6�G>0J�}���� U�#����J�J�[{2y�D�;c��{�w�+��n�1Ƭ�"�qg�i>���i>��~��Vύĸ���GF�6}6�SPU�m��L�<�ܸAZ��8��Hm�����Mg�D���e��C��z*޸o�Z��v��݆��9hB�E�p�U̕���Teo�ޯ(�%�����q��3eW>՟_jSLP?�$	]�d�J��<'�JmԀ�4z75,�j8K_b��c���󡍱�D�ϸ�q��(g�9��㰗�!��Ce"��8�
/Hq��t�|��UhF����pϱ��Q�Zq{���r��
��Y3f6�佺a+� �P6���Ċv��*1���B|	m(\K5(@�`��CfA4�� y
k����U6Óv6J���[��{�J�O�CL~T݁�W����k�W��D�`J#
47��Z�`UJX���1��<3������	Q*ZOɄ=�|X{�wyD�6��L!~�������޷0��Z�7ĩYֲMd�{g��S�� u�5�����N�e�`J�v%4���^Vh, 6t��φ�v�R ܦ@`MΚ/m�/dJ;������:I`�"6�M��c艺fD�c�����z�����xx�۲?��6���[��w�j��2$ӹ�jb!U8Y+ۏ"�cֆ��8z�o�z�j�};O?��"7�u�W`�^��*��[�rN��c�3���Oy$!2�K���)r���\��GaT�5,#Ks65�;�7���!��)­_�)R�� ?b̤��B>e	���Ųt�E:9��E0A�O< � ��u%�r�F�_@����&9VP��,=[��d�Yy�*�s�A`L�h�!�.�(���^B&)�EIl����^J=�L��j�b��~�n�-��qD��zO��1w��8������j;���h��1�z�~�XF��T�p���)`/��H�q�J��fy9�θ���t)��-�]_�B�p��af����,��E4�[�b�
L��|�G���L��N��'�����L]���EyA���j��m}���p�\��>x�$k����w�H�8�[��BL�����]�G�hP�%�gU/�X���u��KBI�<UQ'��77��S�"+m��+so�9�����,�:�a�=�A�\ ��z����1����6���i��D\'wh��ۉ�ֱ���t�6{�C2ytTol�k��)���w?V$�W�:l�φ��:f��mAy����
Cc��6�b�B�7d�`{����W���fW��?c����E����A����b"�99O
ڶ@\f��0֜|�U-7��Haʓ�
{�
?��.�v�[�'%��0�1�ʷ�ԣ��)��Aڳ����,$�s먨�~.e����	�}P�����&����l`v���+�ʌ����3�⣤���a"���{Mޜr*���7`�E�!��&�\ܣr���r����0\*�og��1�i�W�Hʓ���ǷQG���v�X���g$4g�^I*���n�vIe�=�{1]��G�"����w\�x��14a��ef8ݣs�=�5`%-�C[�����O �&�����86ݟU�	�4]����LDN���]"2m�c�B`���H�޼g����8��� &�1��-������ٲ�l��:�N�u��b���V��i���3��Ӫ�a�R�ϿS? �����kdiY�ݦ�H�r߂m|Z��v4&�R�a����p��XK>~��GG�~y�F��!���A�uz�"l�?A� ��{s �L�7I���(�M�r�Y?U�@�W%��	zX�_e��ĕ��7�(!��q��}���nF^8�i��"0ŉU<�W"���m���Dʆ�Q�?���UɎU�a��Ob*iތ�b�k�i12�u�x��X�⁵SФV�JR��aw�FO�w�Rߋ H��oBN����kE���m�ۧ[��l-�����(W�d�������-8�� o-Q�kA%a{ѷ�Dz#Z�$�ŭ8$���2��[���{\S��D �g٧"Nc�Ѳ�}�#�0�c^�埭|��N)��ۉP35�7j̃�6�8�M&��Z��Q�����h��l?[��ǰ�д�+�Ɓ&��,�!��&3��K�,�����xhȐ�q\�g/��F�T��u�l�3��n3r��z�R���#�_�eO��̫U��J�\�R��XB��s�� m|�sA�Ċ�D����ʻ�Q	P�C�z�ppӝ�!q���o�m+�%��}��w��'�YJ���'�����G�yd7�X ��u0ˣ��s�������%B��#p�ot��)2��� c൹��������C��h�y�ev:�+(�Y�L���Fe��>O����Yp���ysS�<x�̮���°RNU�xza�kY��N.��?q~"t�8�;ˋj�6t�+ߌ��"�ܳ� c��C�pZ_&�4�(;K1��û�RS�7�@c$����q[BZ!���Ѧ8	0��[n&�9O�I%xlU��C���׋p��Z������G�B2Z�;z�!(ԳC1��]Y���8�]������&���ׅ*j4�Ж�=F��c�3`��&t�z�1/1u�}�~$��?�^Qc����I���ƞ �msW�����yղ��]� �=X����7�Vz�p >�j8o�����Ҹ���� $GE�BYF�o`�����W���(��/K�?�\PE<q�EX��Z���˨��Z��'��
�C�H7ժ	�\_JjƯ��JwV���G/|N��Gˎ�8N�@_�<���t�q:��#+���Ha�ݢB�ISN���ɨj����E7CdK�:7O�N��_�����2�-�U�L�K�. �R�i�o�:u�[��?�NP�U�{�A�Z�Ɓq���z����#6wCd��/r�|�z�"����նG���2�ݚ��~��qz�W�Y���Y�t$ ��r���&;���!G<�O�p����4�d��}A�C�G�o�����r�trѧU�n�R�J5�K��ڒ6�(�3��S����]��xw47�P�m���8�n����kot���*fʔO`I�'��i�=�g��9�zA�ygˌ����~t��f^��~ٷ!Se��.JA�n �'*�����xɘD��˴�b
д�6	����*��bEw��+�`	Z�kN�9�8�C����}��Wj8�U���:<�Y#i�s���G��A>�<��bbGQ��9^3�cDIp{�7��V�U�z���<���t'W���KՇ����P��0�[� �F��aԯ�|��U7Pm�[ށ��jf����9{���ٶ���h�^�B�g��W|�^!�p�#��#)��Y�qΚ�p؁:ۇ�b�X�r��l��k��6��wk�~��D9bzF�J�}���d����].%��Z)�󦟴 D0z3HW ��i� iAH�V�B�,����1o�\T�E����m dVq$�"P5W%~*#�;�o��1|^l���{S�k�i*DȜ��ӻXWV����(豬��C���6�p�t��F-����e��P�|��#��7�����������maU[4�h�p!g�*Gꠜ�T��c5�*G���nվ���U2PtK��� ����jS���M��o7�۸;�)lB�䜪I,e��dUwYa�`�y�c� 09V��R�(
a�d��t)<�:��S����aI��3�X��Ԍ��f���m̆i��gI�歉[]N�H�_��=�f�Ti�;����٨.�ĉr��-?��q2���O�`*y}�
�_�8�\L�R/����������yF�N����5i=F$ �T� ��W���UB>�y`*��d5�8�RZ��J�`�l�C��.�J9[����apV��r���Q�_$�s'-<����AP�)U���i||.�.p�a�LOj"����s���R��5�����%��Oĕ�#��"<G\����R�\�Rl�BWQ�,�6�dca|��ݒ�z��L\q.td���aw� �+�Ma��c��ȓ�hq�<�l�W>��i4˺9f�"~h�o�>N\���|�z�uR�K>��^��P(5u��Y/�bB� � �D�cg-p:�v�B@bY[On��PQd8��&�)�ᵙ^�)��I�;
��(b����$��ֳe��Gh������Q�f�!7E�+�&����N\��6����$�;��Z��u�N4���v�^�U�L��G����w���cz@���/+킢6N���=tc�BW�4��\i��3��wAm�Z [�Qc�#�VbY� �|�i`�}��(ǃz�9�)�U(F�9�D�(.���XZ>H%�ԭB�|e\0V�O�%6��>�zL�^�'�6n� ۚi�'
�����*y9�VH�j:����s�&(�#�!�[��|5{���7�>�V��
�r����#���Πʚ-<�_��A���AA={�5��B�v��1촮?S3UL_69�{>����,]c@��U��vG��$o�м<L� J���P��y�i���iA���)�د��̪��0��ī|.
��rǳ6���Ig�+rg�2����z��S�I�gbĜ�*��h�4Ps�[V�������TB�w\�]����,#�������<�r�Dv�H�U��M4Щ�ھ�&=3�gBͭ��7�Sc����ĕĕ P -��|��3�P|�xs����8Pn����cG�e�	;��3�4#J�DD(�����,��'�9m��Kcp=�x3��V�X�>�c�v6�iǊ���iڈM�Ձ�]L��2�5b���G�d�V��o+��5x�ky�\�.o� d�[��O{VN[��V��:1k��W��G�����DD��K��/j~��:p���w^�*�*����	�A���܅-쥝�]���BÐ��_0S�6���K��$�d�wLƨA�0�ߧ>O�lg�	;-c�b^D�gV0��4:U
PT�Z�L=`���e�rF�w�Ɛ��Uz�?k>6<���;'S��\�to��p�����k?� VOhPI5#.��2� |�xu_-�\�0a���ݟ4�&���?s�$YT��.��p��8�ƓA�nSAQ�(~�u��?/���sw? 5:�5e������5��)�m*��#V�ڈ5ݞ��``���Qܨ;-�\�k�2�>*w$l��	��+.-#΂­��\N�Ep�6R��=�/r:�n�h,�u�|���U4WV}�2�P{�)�]$���au/��Q��+<�Z&��*��Q��P!C¹���ޫ�3Gݢ���΂�9b!	{�n֩Z��4.�9:_ÜS�s�{��F�Zj��|%�+Y�Q���T�&9I�H�q;�{Z��P6ϸ��I�Fa|I�	#����I�G ���(<$�{��L�_���߇�E|;��N6��E�ۄ�������sB�`���pH��Ơ��ы�E�B^���V�a`�Ɍ�x���˱S��������R��ν����[	i	/��T$Ô�=1D�b�Vh!�E���g1@e�	:�ޚK��Z(���c�T8���R��J�P����y��
6ր@�x�|@��7D�ֈ���Uq�GW���V�I>�ޏ>2e��j�|D5�AciJ�dwC�W`��^�&�P�O��/g~s6p�A� �6;�ZB���z�������6��2D)�3Ȯ�z�\�'´R����z��o�j:5Q5L�*����%,�^��uz0�5�]BDwk��m�~+V�
�~5q�� 3����$Y����N2��������UBS�q�~#��	�i�p��dk��>o=l�;���l}TE���y�j; ح�m�AUL4.͊�չS���F�Ϣ6t�Aﱝ����Ȟ����꺥�W��T�!�;ǋqE�`%t*�!n��h��F��1��|`�3�]�Cs�j��u`ki��u��E=i:Ʉύ��_�;����e���lv���q�xi��ƥ��GBtzn�6 S��_�69l�p���[�m8����Y+q��C��t��f ��O9T�M�+�uR���+���0NDӾ�AO`�g8���l���9R�J��z+߹�Ic1��N�b�(R���8�Sd��v�\��3�S���T��$FOu�Ť���4�~���p��0)��Ը��<�"��G��;�E��a�(��r�ٌ�\(R۵&n3�z%�Nq1{8�9����!��_��T\P�*wAً\�Q	���u�5�[R�Cd�.Sĸ��P����XX�^��^21\᷒7y�VẨ/C�A��aI��b�=�:a����HO�x�H�/	����įD7b����q�o&l�Ԯ��ޢӄ���n�oc2�c�t?}i#/���-���w�߼��\�HA��T"ӎ��bϱ��>d��I��m%�i��m�;p!���KUOٯ�*�:y��b0Vx ��n!�Mt뇔d�]���Wyz��^�49�ah���a��~��\�i�[��%C�p�Bk&;��$H\�a��Iau�'�������
�t5���� �_�J�߆�̊��'Nu,�ŷ��zJ��-)g�R�wO,	\�r K���J�}{�`��YS�S�א��F���)@��W�>cb5�l��5���.5A��B�)��f������]�O����:�1�'0s\��B�!VG�y��*�GP�2:&ڵ�c9��$�u�ss�O(�kڼ�_�҉q�w�q 椱'D.�w4V�i<�\RaJ��i�
�ۓ��5'�l%<8�c�w)�� ] ���>S�f��w5��c�g̭P��DV�4�|���^�����	�F)��]A�(Fԋ?`�?�4D]��<�����(L�D�cD���0D$�'w!����%��\�y�$ց&�U3F�ؙ"�0���\��>��V�:�������KP���$�N 8
eG@hP7Ss�`%�c���`����Fh�]ɵ
2&/�ѕ��0�^q'v�Ȗ7��:��f����P�N�����2d	q�uM�S�X�-��� �xv[5�:�#FC�׿ñ�]Tb&Г	f0��%��8QG]R��9ě�Oz��6H�_9+{�3}#���,Pc�:�c(�A��5jpМ���_��=���iG���!֛��$oG����59�mTm{�vD�'��c���$|T�t��l�=Ԝh�	�ʿ�|���F���a�H�;�mST#�ӫ�
R1�2a_���x�y�62��2(�-�[_S%^�w�41�)0Lx�b� 3�|��Zڜ�tϑ�N�[y
�(���NF@^�����Yޫ@��+9.[�慅�۰�T�QF��Vg)����^#�?�	K?pj��`~��o=	MA�i&�v�io�Zo���{��)f�w�5q�Ӽw=!��є��k��˷��t������fg/sOl�OS��2h�Oc�D����L�?���T�Y�YGN���Ӣ(��B�8Z^^��l�MF�%�7c�Q�޼�s�!%��Q��Rs�U��9�w;ҟ�8��z�:��Y	:�>u���S�<�A.ԝVFZ{��:��y7A��! �a��o�(a�{�/H�����x��{�g��P7�'ׄ��e�6]�%�P�q���hN�K~�ԧTPC;���Zֻr�F�j���a�3`�l?9�X� r���{��S��3�_hU��ˠ���Q%/�wv'�e��d��E�x���i([c����l����|�{>M�[h��������r��G�'�z�Pƈ"JR�<nC\�U�ڍ���x�ax�$΀M.
:��/kۖ�C�耗�?��f�w�0�k���c�'*u��=-�Ì�L���^d�� @-�2� �Ua��|���g�!=b�=X�)̤��
=^N�u���=�2rj�(LV�o���_����3��:�M(����?�4(�E۵z,������71����E����)n��WnYo��ve*R��}�.I�	b\G��y����"A�<�>�F��(b�ku���̸|�S#��DV�~t�_����Z�@<�޿�~r�t!Nӣ
1�m2  BNa�����������L%�g�y�����X/�J�x��?����w<����=1�v�d�Є��>ψGRikc�\1[��|�?�w=��rXa�}����L���ب�!d�V��N�UZ�g���;��n��,/$`s3�Ex��:��`��8g�>H��l�օ�˖Y�:�e����ŵ��.�5�{D�EDR�w�Y..3Z ��D�ߒ�T�>+f�2���e�}�*b����.D�M���q��\Z�dQf�����(L��/ܸt��bW9"2���ǫ���7K�q���3"*u1�����X��6Ò��zl*$�r啷��ݑ�K*���k�Z�~��7m�/��v��3�h�kVclhG�G^7e.l� ���:��UF*��Qd�F�o���/�{AՌ�Wz3�W=�n�^.���r�C*�IKM'{���4�+�V�:]�p�f3b�P�^�7�B�=�>�n�x�x��J��wɋH"a�GT�����L>��X$���W���ܫq�<�ȷ���CS�o�r	�F��:Ѓ%c\��*�N�e�)D�5�M�U�m^���~�I�!�B.��9K[���������{���G渵}��:���o?�Dn���
�3��UA�!E�bF�y�v�G��@A>u�i����Wj��~<�V%����dh�p��5��,<~@Sf�^+���[Yy���OE��m��h���śܛ�pz�8^:���}� A�s�@��d��-[m��]Tߡ�sg�� 1�Xٚ�f�w�KO���N_��*�GI$AB�����K^pG� �\Wp�le��Eυ+x�$6i `H��]�����&u:�c�A�#�Z�h�E��^�| i ��텀��3j�0~�L�h�v� �ِ������a�݇��#��
%E�,!
�iȄ�Y�M�p`=�&����&ςS�_�B �vdU9Y��Y�M��Yx��KN���2AZ�h'�\,Q�U`9���)@�+{���w[�gȴ8���|��~9�o`|CYV��Z%�9{�s�S|(A�@V��<Y���OtL�����iR�8�>6��C�� �xQe5�ہ��En������GO�U����6�J��)�4��*���a��.)��/��	�#�|Լezd�=��DI#��[��쳢x����Km2����B����X��6������R�<�U��2�b2�;1�y��?��b�~d�RIq��e�|	<�;@�&���:�:fL�U�P�0QD���J���y�a��*�U�d�[:2+T�Kgf�^�NtE:K.�5��T������u>��N=��%��c<WD�Y�	b�rg��`���)�8!a ΅����ߦ�]�6 ��[�D!�q�S	@=	W/���%��iC����m�ȍx?:fk֔�@�����͛��X/�ǎ�m�b9e�8\wF.)��%�H�LB��o���i��i_T�������0�$`I��x����k�W�}u���#�\�
B��M�w��
��*�����t���g�����n��?S;�g���O�Ȭ��o[H^O������ً�
��AJ��n���M����5�5�&A��&�g�����q�!�'����	�uN�kZ�0���ykE�p����ۜaI��A(0�������t��r��tI��p�۵� A�pg�q������*B�͉:i��3���+�v����M�����l4[:�&!
8��=����Ĳ�~�;���X*�~[���ڊ�N�x���)|򔈷�<H�K
�z ��Χz8��ݱ0ҿ;skt�����5�M.(@,z�G������@��R��B��� 0���Ō�Č�֌VʋP�KA~pG���Φ��u�_�l����]w0�����4���s>��D��Q�1��?����z3����/m�8qC���3|y�6�ٝ�!1�f�1S&�r�dF�l��;�Y��߁���i�iXOr���`2��76��^+��B g+,��G���}��`�/�X�6�V�+Uq�qi������ц�%�U��ϝ3q-r��+v6YL�vL:Z����rX�����Q�n��g@���W���)gZ�[45�'F�2��vP���N�w��b����5��(n���k�
�j��v���������|�y�ӻ�F�8�I�4V��<�;�>jA�(C�U_`x��LhR܊�I<!瓴� ��8�h|O�$46T�3_�){h����B�^�d/[(����7h��N<	o&k��S�G�L�9x�J�_���9<U�07�[=%$�JC����G�9����W�)�Ե=�K���<"�	�j{KT���Q$
�C�?擓�^k-;$1������2d��. d�!���*6��9����_�˨i��H�%҆,��d�;͵H���ߦ������F(_tcs��ū���[@ͻh���2�"�(���A]l`�4��! �����t������
�˴��9c���3KCC�����e+�1DZK�ʶN��UW�����[�QB�����}+8]�2�\���L��j��ܻ��P���C�D-
�<���@9;H�s���^B�ƩcN1RA���,5�1�K��Lr����K�e�,c�6OI�k�b鴱t�N/��ȼ��/[}xS�<9����^xj-]��o�ڦn���ޔO2��J�'z �e��a{X"p����;��ߨq� }��I��੾���)�FZ�|a'�8(�7:��i�M��Ů���ƿ�BL}��]�i���Yƌ?i>��^fx�=�����=�G�MH6����C7��:1�0�3@����k[��?H�6SA��K��ޤXR��4�܅^.�Zw��D����Y�x۸܈�# �ǂD��:a��:�1���y�8��k��i��&��(J�5Z(в�:[�kA������7�Z���I�UQ�������[n�_.�q�������Pm>�p5G���%}�ɄhK���h6�zwq�[Slz�$��ʔ��y��g�4� ���C|Ӻ޾����(n�q����n��*�A\������);A�_�t{��M���a(F®�G�a�O��fqx٢�Nd��?1=�M���_-��Y���Nh�rk���H����G��Ӯ�Pg�w��1�,J`�Ee���������e�O�ݫ'��]�h��R�����ys�eY�$��;[]l?��"�Kn/JV��iVk�o<ar*��B���tX�ҡ:<f�	9>W$�e������v+
4�(��c��O(N��4����=����7KeG�����'$eQ�X{��|(1����8c�?�y����G��Ye�	���X����X��!�&w����͹�`���QI}.�]���Ŝy��f�%���&,�$xڰ�뫪G�jƢ���.��ԝ���jR�GzՋ�M�u��g�_�Ƕ�a����$(B�Dd��P��33�*(6�,�0��9?9o�z4^�S�����y�7>����y��*"ֱ<h#����%R����~�-�Z�!��U	"��{N�#n�������Y
�����i�V*o�'ԑD�W�K����p1:~f��]K�o:l"�մ,H�5��7�%�{�i_�8���!x�*qEп	dQ��EٮYɌ���;<;�]�P]X�7+eLT	������Wկ�n���w���Z8���^��M2�n�v���R���[�Z���GX'S�5�^�L�e�-LD�ژ��ڶ:�f$+)v���V��E�׉mU�V�CtT���/�}���ѷ�(�Y�n/�VL�Th�:�Y�H0�>�� �c;:�ݏ����%v�V 7Ԥھo	s�{F_=�Z�f�hw�3������p
ZT`����0��J�t��m�B���ླ�Ï.r�0���"�vp���H=���}���]�[�}��rXӣ�|G���lDA�W������	���q��՚������d�i�BU��`���o�\S��	�a4�$��>g�N��K��{#�]�Z��Y�����t�U���W�����M&X�]��v�?�[m�)��~�p��t���:Ա.����!����npۺ?'A����'�m2��骷r�i)�i	����U�PD�f%U�[�O�:��D��m�;x��y�\� ���߇fa<�P�yC�%��o�JFX���j0�L�iI���&mNPe��&F�D��Wp��[`��� L����oLz�v����b_\/S�A�ZD+��T�L�׾}Jp9YfFC:�$����V��S��ć��Z�я#tn������
G���0++�k*͝���[`]?I�T{(ݾ�A`����B+3J��y�-��,�:�]�F���]bS���e�C3�?�R�A"�Xz� L��<�;�X�Pk�a��'�6���'<�s���1V(ݾS�l�J"�5�4���i<�>�����W�9�݊��6@H�["�*Fd��(��;�=���N�2�N�n�Db;@9��n-v����d5��yUw�%;2{���#]+.2n-r 3�>�m�J�����x"�b�����f]�;�5e�暁�A�CU+JGò���\+"s2l��'�Q��J&����aJ�h׋iTZ��s�
���6����^�h��Q��T���^(�
���OD��'@n\�gps�z�>�Ea�s��%}"���j*ϡ6�ܛ�[��R5��� f��G��<�@A�f�N�CkN�0GH=xb��,�m�JKi���$��d<
��2fC��-��(�J�"-K��6���'\.#a{��������9y�s�@�?�1�v#�
�9�^�be.�6Yi��:|8�N{䄄�G, ���!�g�{��=��fw[���������O��t������W�o��y:Xʥ�g��;��%��/|"
K<v�I�h�*�;W��F��v.ű5d�堊ao�%΍��"L�=jK�_�T̗A��'�n��)�oQq��W`p�ܑU��4 ����K���6zS��i�rKō�'w���3��8���#��S�Bg��oP�ʽ�B�7�y�{���oU�*���\�pf�r�?��?7z�i�'�h�� 0T�7�r�gB_̃A�M���$�%������i�@��v%�	���"�I퉏&Fti�\G�ұ֝�@pa4O�hT��?$��N|\��9���^��4z9X�h�P��9(��	�� ��|�?k��'�J�dj>��]S�뷣re�ߩմ�(jax]���3Eoܻ �Ul�j�S�����Vbm��tv�V��չښ\�X��-��,��U�H-���1��@Kc'�
��hn7iz��J�Ge��f��x-nl�;a�˄�CѠ��ja[k�S�^h*�m�Z�>~@ d���|��
�'&����)s��������H�ӫ��c��%�i������hM��vg�Ro:��mN���4���!��S����f��?	p9g
���(+�l����4:Fy��E��r^��=ɶt��e�';�(@ܷ���r�����z+ұ�M��y�jU��C�9�4i�ƥK'��֕C�� ��=�fϹ8�J����D��f��GpJ���U������{�O*b $]r�����Ҷ���F��Y�4¾j7����>�[�P&T���<����DH`#Ӷ�+�g��Ɇ��H�R�`�S�~�2����㖽U%b=;Ҧ�.M���NGp��X�cs�V 4ϩ���c�s���LRTnH\�tS/�ap2H���0IkS	�"�8�ɼ�I����s�_�ז~���`~֒�N�u�V��v��G���B<�O&�w}M��;.F�Y�%Z�3�#�������L��)���آ[��0٩��I�ӑM��v�(�`5�l������k�^O9:�esɻ�
? /�>,�>�=��+.�s�r���~St��^)����L��N�ar�z����"�y
Sߢ7���3���� Sxl|� 8��j���r��:E?a�����bhbTyy޵�\>B�@^��\l#L���}������%I�<G����!��q�xK���8y��b^;��s��K,m�d�ض
Јt�H]�� ��g�y)����E��nP=_�P�|�(+쥥���p�щ����5�*��)�\݈�r���oEϜ�Y�C�/�kuC��(�[��UNW��^8c
g�����W�@���T\"����vv�
�y�o&^��`��,WK�cH�xokO3I��z�ߎt��X��� �� ���o�l���9����g��nPW�ut��
*��!{P�5��F��So�?m?/��"f�Ux�֥alɂ�-h���W#�n8�C�a��mf���:J*]։S^�o�\���44>B:H�Rt����5AYr���2l^�n@_�w�&.ӭ�*:-��ԯ�S�2K�t�dW��lU]��\���02V��ۣ��[?x�,��-�
� :��&Ϣ�^���V��.h?^o/R�r0Y5"�ǹ�D��޽�t�"pÌ�^���W���m�'���
�k���+����hS-	k��BT`�??�2��a/����`���aT5=F:�%�����꡷�f���(#"�����2��0Z�tUWo�ZJ���e{�ج��\�9@qgy��.A6B�y����ج��s��Blsjԏ��F�-�ўa_z�Qt-�bX�dyz7q_�	���1�ö>���&�j��!=�������[ߪ^�o��S�>#�8ڞ��O���op'�'@,�dٚ@R��rm�&�Z�#=nM�������ooCN�2��X
s&�Qo3��Ŝ�3:�>Vz��*�mx͕�Ɋl��+rJ��o��yC��4�}�y珆�#�W��f�cMڪ,
�=���˹�P��ؒ�y��Gp�=fgh�kY�t�+��e�r�� +�O-���rf(+o0r��h~^v5�f�H�B��7��V�������ώKa7R�[���}���*�G����#��:��[+�ȉ,No�n����~b�n�ҷ%��.��x��4��UE��Yf���. �H!E�y�}Q�Z!|������2��Ch�RzCH���b�������s2 8J&�Ɏ�@<�o U���%B�x�3[v�K�����$�Ǿ��i ��k����ۚ���4�'g�緢x�f<�<�.V����,V�F�S# 鹽Ii��~�u@�[s+��.�؆^� ���º]OV�����RW��%m�*��`����m��-2-`,O�*
@A8���;/�c>�"
	�A9 =��LmOl�T2ij0�$�ӭ,���Zz��$���,��E�\f&�P5�>����NMb�bi!ţ?���<D�9t���b��˩K�sIU�t}����(񂙇T�˖�z�U񓔦ϰ=l��=�J8�P�p�&>��K��؆�	���7�jnԑ�$b4����l�5D����w�hc{7��9��v�<���m������0�Ha�o�%g�,��� }��y�k!�V)1��zcPT0�4	0�c��Tg��s}ڭ��Ϟf��}F6�^մl*١����N�δ�MҀ*<��JVa^��D3R�g�ߎhB�s��2]*�=3�v�Ou0!_p6��5k� ���CC�o��Va\7)ڠ�5VI�d1�C(�>~H����0��v��KO3������Y ��B�׏��@a\�&������J�|���bΨ2rdfS0��i!8���ͻ�XfW�η���֟V{;;�Y�M�f��*Y�<�w��e�(�Ἓ�v�8W;���ӏ�l�-M�����H�I:@�&��5�	� �E���� ������Y�#wJ7,������Z 4�Lm���n���źSal*���Jm���:X}����� 2�f�И��$�� �ŭk0����\�@��V�Ug����D�M���v��	�������˒�˄�W�-\T	��H�yT�y��j��S�F��D��~t����o�A*�:�ܭ�~��J�@��g%�"̦�x3�L��uo��i��*��4|N�;҉��9g�� +>7�]�s9���Jy��!G7ѽ��I��$���o��(��-�\IBl7C�m42�K�Z��1��Fy٨,<��C3a�w��R����bw� �j~����I���f��=�@ᘪ���;�&�F�׳�����-�5)�6-�J���\�NW����ƻՁ���t{c�^�h�P>�٘�+Z���`t
���-ef�4jH��w~F̔G�s�k8>Y���'8����j��$)�/����6
�Z�ԁ��� T�����.�c�~k%���� ����D����FN�+u������<B�!J�F�{�	*�E�u���-�v?o�3������A]3,	���G	1��z�m���ItI��<�,��%�ݯ��Izr����hZSU�3�>���w���l��o�e�z��������s&���-W��\����=�w]l�Ξ�����|Ib�s��j��&EZY���|�0cq���!?�! �+���X����;f����.h�ޒPz׏���*�*[f�:���z��X�$<?A��p���3�!��i$�<���x�'>�2~h.�¼��yB1���!!�Ku%�%v��q6�0�m��'�|�u1�,���~m�Ꮢ��"��G yn� k���=`@G��$ ar�VM�	 1�Ʉ��.�B�UTw���rd0rk�Ztd,��Ğc����I� 
g�-���u��|$��c�B��*l3��i�2Y��ǊR@K�G����lΣx�E28�B���Z��|�>�(>Ҩz��^6L�f���l2���B��r��^��dK���#�-���*�nM��!�
����`�\��D
Đ)~�U�@� �^T�pri?D�%e�J݈%�1�v�PdO�#XW�q�) F���Ǵ	�+_���y��K�0��	ߏ=�	u�:3��d��0�� �R3����$60�]�B?O@���z��������3��0�S��J��)m�J������)�K��ܳ0V�Dl~�7�U���m'��'_^�ì�C��|#�_�Q���䴆��X�Q�#�.$P��4�_��I�\+Y�5�����D�$��P���IX"�P�y����j������x������Z���������g��X�b>��JesY�����a <r�9�n�vU�^�D�\����p�������Pl$`��FXA���o�QM�f� |���<� @��w����(����z�؃얟k���C�c\s����_{��c`�R��-<�?u�X�_y�>���=�9P�ZԤj
�R�~'3���;��{{���j����]&pt����'��F'�r}�a�����F�6D���3+7�Ղ�4���z��Y�Ⱦ%����Y�@�H��:�T�	?��v��XcY�RwK��g��ɳS-Ǐ$ڑc����<�۷3�Ȳ|cg`G���%\�]G��;{9V��<*�����N�߽7�RU���i��Ҋ�K\�+�ˬ���d�P�)$��̖G;���W�x;!��91�5·�������2�	烖�!H� d�,���h�������TY��R����M�T��OGC>ag�e��}�k�N��sdA��D���?��,�� �����D�6�l��nh�چa"@�{�v06��P_�9���VC���o@��!�I���J8�G���}�6n�� R0��#s5{@�3]\��^����+ ĕ�Cxh�F��Xt`t���x|:)o�AY��Q�BkM���p�Ͳ��O�>S��<�g4�Ux�fBgz/�ݠ�2IPm0�3�A<dan��!rc���%�n�P���7P(�+��
,�����P�i&��ޅ��������ʫG�9��$��!8HL2��f^���%"/˿2�ӈ�Y��~���)��{-��e�Kg���2�N嘇[��ɁP�@��k���u���C"��-T,�8v��,Ԧ{��^��f��f�eu5�Α-�1<Ũ��JB�qe�ͻFr��7au%e#���v�dޑu4ve�s����.�����T8a��Ly�|G*��n�uO���� ��f�^���l�2���x9~�[l��%Q!�mXol<��\e�K8Zj���>��pT�R����������+~\d������������bP^�i�vc7��x�`���ī+�0�?Tj�uJ��<��*�i�P�����C"ɭ��C�
I���^��|{�SO@;Oa1i~.�<?�-�*#'�P�������V#��z��#�l#��m�~�![Hh���XuO�K�n���v���A#�0z�>�k�Ԅ*0d�����/:+c��8{��)���_� ���D��J1ʵ�=�*�[16=V<�K�6���ubH�^��ҹ�G�k��� ��{�Dl�ʂc��;���=��P�w	 J���Y�S������et�6�7�]�1�ԛ�b�7 ���S�ӄ��+8�b>/ܰ��`���Ui3o�=�h1�eO4T�>�&'sC�-A/�XȬȸ��?B�Q�$\�&F���Y�_ZI�Z�Ww���X�XR@��ه���΀;^����J�c(T��'_j1�f&(i۟%|}��)� �s�� Y l����:�T?���g�1��4��U)TY�� �d�[AM����(�x�!�Yxd���	Q��R�u�J�ʫ��nW�ތ*3��1� H�dJj߃��ԟ9RBBr~�9�8�1W���y�P�@��qRg7S��8*b�ofnТ%�C�fAI�P�bxL0�]OW�ȈlE�h�ŉ��s�}Ɛ�"��)�O�x'��g:��$Bi�zi!�"�i� Z���i���7�wJ��uvںO���&��ȧtu�7�'���F�S&���:rF̭)��'F�j"�Av�Q���s��;�-���@�yh�+g�d�c���^�hi��_=�?�oG$U��y~��!�IKѱ������uE9w$/0lOO�yC����V���$��\.ԛ��C$O��=3���$יme��L֘���%��N���ɹ�0��M4�q:P}ƴ�&`��aV� 1��}Q�\�k9�7e��J_�H��A��wj��1�Ѽ��|��2j�4N��R���W��s'��C��<����-f�U8<����|����`K>�{
���f��ԋJd3���;|[:d2	1�5�%\G�"�|�0��>�T�쩅�q3�����!Jq�V�#~��3��B[k�)~bn���|���*${���VN�_����ܓ�Q�y��v �����LPF�ư�1f�����BAD�Z�W$�԰՗'�{/.�;ܢ]PoѷdRrwQIS���(�����w�Ht�g�Sޯ0�`pU�.�Ӗ§���Ǐ��DZ���,8�䩔6T�x�-(\��N��e���^&yO'�b���SU˅z � ���ȼ�BO�b�q~M�S�M-��l=�MhtT2/aI���K�44��O@�>-K������lG�u@��#ا�׸	����B-9v3Ȟ��Pb��!,��$Ob*d3D�PÑ�ረ�VW��"��[�� �9����GF�v�:"˛h-�H�5dH�Zga��}�W�i��ˇ��^~mFC��Qx�nV�!_�N�S��Z����Y|l�G�rLb[?��1Z��Y�J4�g���퇂5�f���Q� 5���ਙ&�X����e�f��C�<��1�H�ڥ�:���m
,#��S��:;��s?�h`8�xJly0K�u	�Z�9h[�Lh%��pX
t�S	V>А����=��]]!�o`�z����ߝ�>�$�_�?D��J�A�3�����hK�P�C7�B�cx��&p���Ft���a���P�vc~����]x'U\]S\�.`�B�1��Z�~�aN�5�>��dz���e�E�H�0cJ3r���2��"d���I��[GNLx�pZ��Z��shYK+��NK��Q�=Ș���e����:�ۏ��gJ�r����(����u�J�ߛ�:0�j��I#��+��F���I�K%F�Wbk?�� ���9�O�O�a?��|�q�Y.��V�k���z8���J�e���=>��?����4�(ḋ"��o�ٹf���z_XD�)��MH!��t|�F��__؍��&�ɄF���C>&,s�J?�$�p��c;�����pT��sn��
XX�W=#h�z̐�&�7����#�P+��MZG��*�9j�����Z��yX�i7ѕF]�p�N��6�_=��7!��\��g����,J��&��������������{,�Z�V�^o��Z�&
��:��}�f��vkϙ;	l����<�H+ P������eh�݁t��6["�#�'5�j���}8��H'�.���S׋�5T_
1M���)�Q��:\�U6nߌ>	3��7������/�-vYա���$&���q���!���;*oK;V0��T~�4�A���u��-��bMJh��kIb��z�qt^��m�u%s\�YV��0�p��� t涧��g���2F���MfR6�)�f�ޗ�G��r�*��FF0]�paV��lZ7��r�+M|�� ʭD�BT+��i+��y�����{�|FuE��"WÑ=�fXA@ľ�	�R�tC`I��y�Wx�K'u�b�Z�T;��]�hb�Ll��yS%dF��z�vk��.,���]9��t(�{����k'Ǡ����y�H�\�����������oEtL2 �i]�P���4�[�2)�3�*��\Z���_IuS���pi�����J����g���@(��H��I�e%K��"�
b�hX燕�7ϪީT:Cʶ�#i�nd�p�w���Tܪ.�AYⒿ�<�k�6�_���Vu%���i���L�GxY�MZ�=���I=����դY7t���bzɏ�D�$E�x���L��'��x�j�gYX��2�\$LD�_���4��s"��vM�ͦB�C}=�^�ĞфI��^��	s4�24t�W�hS�M��h�<ͪ��0o�9o&�^٢ �#<k=���4 �7�\崍U�`7��,�['V|n�T�RO���A
�mj?w^v�6 k��H�zL��_�ε�Ĥ�N�P�����t���|�Ń!��Ț����e�>D�]+�]��%��;����uW�wѫҶ������?H<�ż�AH�����,v�~�� �H���hw��ݸ=��Ӛ��c���)��xN�d{��g��<��I0�g&���-�0]�[�*;G=,��}覾�T�� Ad���o(��P���@ԕv�Z� �r�\E�vu��<2�`��}g��f�%)�@n�6���Ȉ(w�p[o��+X:+�4�$v����R�[9�0�j]��ѯ�J��<� J�yR
Ek�`�+��J�����kYƟ�UH�L�����	����$4��	'x��0}hO���`0�������2kL)��!�sC"���m*��u������85�!h�.XE{-!��O�;I>��\�r��ݐ.}r����h�po<��b�uN�+9��	�Ln}^��=�%D_V����<;�Βh��V�z�3�DN���mq����o1�!�4�å��׼���g"+�����w�/�t��-&l$[�v�oi��F�ۏ�NH��5���jg������X��>�U�J'6�E�b��(E�!b�ڝ|N&��oh�e�c�n� ����;��fK4�}�v��Ԣ\��.G�T3jS����S֚�LUߓ���~��)T���>��a����Ym"���l��r��c�'�r�z�d���@�S$ۂzS��RTz�.�8ǖl�{ʳ� I8D�(2l�-��޷��kRw�3���$	��_�ؾ�bk�}��hkT?�%�6�� sI��k�d;^p���xt���ӟ����ޢ��km:2�^j�L@�F\��<C�g������d�>e+6h�+�
��Ь������?	������\/G�9#9�U�&^�tɥki�Tv��	��k)n:lg��9z�T\'�i���\��`�]�3j��Xӣ+!��R�Q0K'� lO���6��Ѻ�*n�,�,�Ǔ�I��	8�˧_7� �Ԇ�ʇೂ�&��h.	Mi���h���$�&��!")�=gE\���K��gauy�*������N<�sle�k��x�aF��%u��F��:lY��MjD�w�v�dJ�:���B	�N�{�aor�\6���£���}� L�ٽ"�]�¡I���]�ݸ9Y6��Ŧ�9f���L�vr�ċ�����D(Δ��ZN}�?��G&�u���a�r���x$�of�����4%��!�M�0�����$��E"
웈�Ef�S?��h#D��/?����i3��R�<w�\��_n��f��90������>�3ou4���t�끑�%S�?�U�2a����B�a%�^�9K�������p�ѓ�т��H�/�w��i�;��d��a�z�jYʚ��v�[q�+�)8��D�RJҎ�h(XS��;���
~+�[#?���k)�,ʇ��A��GaX�aDx�c�L,�U�n�Ĳ�}�Eis����m�L���@����X��j�耿�
M�l	��
t̟�k_uQL��D~��˥7E��7�[6{a #�<�ȶ�P���r�������)�@П�w�ȷ�A�攎(�Q�<n2�e�k���*�$)�P���608�ˬ?��c�G��<B���Z����[�/5ʚ^=6�sb���jBU���-%s���K `����M4i�;ŏ�I�g���bhϼM8w�O����f5�:4ٔd ��Fv����ġnB?�/�0���a��?����.S��IzQ�����_G��� ܧ*%@���Sn�э��J�9S^YӜ�'/n��, s�����&��zn�F�iG!^_��ǹ��H�}}��-�G%���.��z�~0`+T���w�ǔ�����ۮ�%���.o�?�g"�r=C�PAk�"�E���&�5Ax�R��\/��ҫ��)��,��m�0U�\�i��Z�L,�V �,���x5���������"<�|��>"�+�&
d�=�:������$Dm�д��$��YL��±�8s�J>�B~Ry�Rq�7n�����[�?�GU/�^`��#iEc�V�����S����B�$�k����{�h4�i�X��Z�����T�6^ø\�щ�龙ͻ���ׅ��0|�Ә��+-4Y�!�}IqV�����e�l�9�� ��D@��X�y4����8I����]��M83���Y8	����k$��"��9w�CP��J��TIP�ݔ#p2r�x(a�"��%��0�+eW����t�rH/BN�l�	 d|�B}C��S