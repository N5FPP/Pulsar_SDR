��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��e�ik3�������w$����g|��J^]ؽ�V��S�j��������)vIV��N/��~�@ʖ��-�����=C��(r��劧G�n������r�7iD��a�)�O�~�A�� G�Jk��Y�j���`�py".�}��**�̤��=���%�M�2]�K0A-?FY�M�Wjۘ_�7_7�1�Mp��O���:�KH'gAG4nD��_>��7�aڧB��&�}��A��b@��]��̡`Z�Ʈ�$GL���4��ϵB���̩�@�"��m���=�q[h&�N^n������u.�(q?��mC���0����$����|�Z�V�>��|7|�*�[���}���C�g��^�B(v���Rȧ�LCE�-(������I�`���9F��V���Po���%�3~ƾɞED�_1��G)��;�!�7�<����jS6��lܞ�ʄ�#',+$�<6'q�5��� {���m���#��^�DJ7q����/}2�*_a-�E������㺗,���3�٣�k��¶����H�Nn�nrI����P�G�º�4�Fg:0�IRz.ʒN
5�o�L<z�.��^����벬�P��漫�fz����T������(X��]��r�Xdm[0Bz��+QҶ�+Sj�>���3����t�����r�&`1|���u9�5�b���"1q�*���޽����5�!�����1��j�QL�k�#���٤w�ZB�!-U\r�&?'�'�\)�ɖ{�q����%��Z�'��1LwzSic�d��[I��>�n�W�������As��E��Ak�PB���YT+�v��u��d>�,���$�D�L���xςq�pJ��G��;���"#~�����&m�qj�i@���	��`o�p4n7L��U����W���{B�Q��o���!�5	؎ڤfʳA�~T�#�t���E�jF�Q0��R��Ĳ����l�G	uW�ܰqW:��ށ��s�Iwߺ�3gУ��CԴh��*V���>�*⠨!Y���y�LV���:����e`C��3׿L�N�,�u�����c΀����lrK锢����<f�����t�!9�����I5�"��37f�_��ז<?�55k�o�?���sF�s�S�~C�Y��w��h�FҠ�5��*�1%��
���pO�s�������q+~��m��tX��s��ػوt6��9����I�%���j
�)�$C��O��.>�Ph�W]o�}����:�X� ۓ[K�
D"bXP1-����L�y)�Ǵ'f�bO^'�R]�LG����am� in����G�cv���$��O�+̵ziOI����IWy�U����D*��[��8�V?����.4�+3�[�49�Qz�1鲸mt~��t�.��Y�N^tB�q' D�@Y|�NXփ9�16�>���Sa�-�͋a�s�����u��J��!Ψ��Z�U�D�}�a[\k�:7�	j�+V�R��=�jj3��+Ѓq���35w7��	ەK�PD�$��e~�h�e[�U7�1v�bn�7>�c
�2�F�"�#ws�o�eW�@��[ �gS�Np*6t����n�B�>��|��q�=� An�9w�N��zc\y�6���#�ƪ$ma�R�⚬a���V쐸���!�?���p���%p��p�v`Ud�ڷ�+s��NϜ�+'Oq�|V#��  ��?ӏEu�x"QJ3�UL�-���g�K�vN���Z�����Cͭ��g�왅���P�f8���)�����H��/��L�12'�e�:�澋��=�v۱&��c�$3�I��y%_�(uu��ǳ�N���^Jj�Ty�a��W4�BS� ��kC+S[\G���u�N3�\- qou-�t�`��������l=<	���x�s{��i���lJP��p������ەd"'ʠ�/�WY����^�qD�|���s.,�x���Y�Q��6os׺�ZқJ��K%(���`��BVA-A5m���d�)�ٛ,R�X�������bh��~_�К	H�����uײ����F��{��;rLq0��l�,R���]��	��|�޼��B�ܩu��=��b���d.M��=�%��׈���o!��֝�σ������ˣ�3�t2En{�G^�l 4�obb{�
hd�!e�;�"5�^M��^��W�����M��l�����Mβq�ڿ��r�o���CQ�_"���ԩ�#UAt5Vc����;��Z㠇�-��N��Lq��w�˱X0K
i�|lΦ_pB��@���o`N��Fy��ݎR���[�ꖻ|�N�'�\�Ɩer���p�����}�c�oK0&(�+H������Fn8A���Z���6����6��?�&�e��/�d��7q������4+�7�WF�=�6�KP�K�/�>�.?\�{��)HP��4m�)�R���٦����.��k���b�^:q��6�6�\`3��6�f`%J�r-�o;gPO9�b���fd\v��k҄��� ���fN�;�u1�]�vZ+��wyt0��mkH����u��f��M��mH*|�,#i�.p�*�����^?N�S*��>R��W��ӝε�(X"�{}�}['���5�ygQ�'�_K$�B+\B|�,$?_rS�����͈+�����D%oD��n���!��dQ�g�gUn�
������g��A*��	0�;-����h��m���]�7���ҧV��j��MOӍ�Io��`?�ӊ�6�^3�YM�YU�>_�a��5d1��Y��>x��<�ՙ�[���4�f�\�e����kD�mW��xLy�f����AaR���GĐʁ�����7-Ȥy�0���r���Z���X��?��}�S�KN����OX_먼�|܄�E��7����-�E��3KT9/ȼ�E�
Qa�D��:�FHۅ�5D�<_�4"�Ą�f4��P�QV��CSEž�0���Jk:�z�_��.R�
o{�H�_�~{ki�7�Hܐ�`�.MN�,٤��e� �=���?�H�