��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY����B|����c���!令Bh�	 ��H���TR%uom�ʮ�Y�*���{�QHw��Jw�}��N� p�������Iv���ʪ�"�^q���[�:�M��ݘ<̞0������5[G�	���p�S�Q��,U�H�uci�h�\�#k�\��8*��8�΁�	�
$M����ۃZ�;�?|�ŗ�@Ja��h�K,]1k�"r�%�K���[�>ֽȪ�����]�}�ل$7����6���o�G�VJT��a=J�,bc\�!dvLc��R]pc}�@���s��lmb�XE�g��Qڗ264�=к���l�uIԕ���x ���3�Jd��x@�C0(�{���O�W���}�R?ϓ��5z���3\�I�������W$�Ű7���4�K�EqNi��D�xܠf:���R#��}!V+��=�9a9|2Cx�8�Qe9�zG��e`���n�㝑���<�療��lX�ˁk�s�=�
1>�.��Dj��~���SJ>!-�爌�_������f�D�$�����\����h��+�E�����#��� �8�v��	e��]�S�'9F�Εl�ɖ�Yo����MJ�p�G�La.G>Z���X�TI��s���y�����ÿ�	U�KL&@�,�9�����3��P�&� x��d{+�z=���d�>q&�B���7�E	�_��m�W�ߝ�`3��W:��	)wҞ��wEⓡ�c���Qk�..�H7�Rܻ�����^\���y��C����K	����s&#Kv'�=�=#7�ܻ�9�	𑃿�Z�c)RY��6�{6����t���B�EL� �;�Q�c�u��S����̺�$���J��X�ֿ��$�D۴���ߔ3�v����\Okw���aR��B[���+ō����qè^qp#,��8P��&V��X#���Y<k�-� TCѷ'�O�e~R�S�xoME���~��`f�M:����M����l�I�.R�vW�Ӆ�J��LH?:b�ԘY�Fcl�P�6�CҜ��c;�˓��L��'�!��d�|C���l{�������~>����¦�/�5�l�ݘ^��'l�w�s���#3�z��gk�K�i0:������p�p}��c����DR�L�Lf��s��ۢ���o�	"�g7J������1ӱ���"�i�dD]�������W<��s�:��\Q��4� &qR����1D��J�V�	�Ɏt�T������H�~�)�!��±2�{#�3��t���d% F7���X|<��$l><��F�]�R�|r��#�r��7n�'�B��ƌ�_�!�A�h���I;�/y��K9�/�;=�7mC��ؗ��j,���/��>t������\�mế��g˷�o����&x �)ߺg�)��>���A��ir �ײ&<q!��@{��3 8�^%P��T.��������섙F[��?}:c?�S�\��EOe-�xŻ�>�C�d�;�����6�}�����Je�^(�hf>p���}��w0�XLK<dE6�N�@�Y ��ߦ����1���L�O�Jc�:hx�ც++�|R�k�b�ޓY�NE_�n��O(7ъڥ�"Gr�ȇ����T�!M)y��X-��ؚ�v�9���, ��DB��	�������J3X�g��^��׬�@*���\���g�+^�"��\,��HyQ�1�F-�����s�B#JܭĘ���H��v�:rX E)Iѕ�\�_i���j���	��_1"��a	�O�䩗��.Q�������z���9o��mF\�p��.ь7ڪ�nT�:�F ;OSe1�j��Ga��o�"�{b�wj����V�+Ee�D�)���ײ��>�{{�G�*d\�g0����y�=S�Q_|M&���O)����8���/�oG¶�[����*���*'aG+7~�,E���	��7|^�=�Ѥ�=��#�5�]�M���jg�1��i�C�DY�0�����&�C�uaI��
�	faQ��ʧ�
7��n�@E�6�Ly:o���A�#X���6�^���q����}��d���h�+��p�������$DŚ"��U���Jg
�m�е��&pI���	�-g��KS���8)��S*4ƫT�l$
d�y��9Ѫf���Wقm6�%-`$������(��]��u��b!f't����*�Пl��)�t\V�l��	�[�T��u�>_Թޤ�p���:�^�N׽�'���Y���p�Yk}UI�����fְ��7��ɭ?�d��B�h2L�J�]oP|�X�����\l�1ʬB�A}x���}^�rNi�ZH���,��P�yNC8ws�qF"�\�r�й�B^B{1���ǒ��tL$:��#��_�@V?�j��
�ږD�"�h;���6.����r\�pT�3b�դ�u��n����-�.|�+��� �m}�P�2Bӂ"x����>Gx<cО�#�:r)?>���~���;7oR�2���-�9��n�5�p��~�_��<a?�$X���!��\�B��*i���C�Eķ��f	 ��OoT�tV���)�L�(b�eٸk_-[o9����5L< 6�?�Ӹ;�����!	��>鈯�v�T�qL�Y��'d*0Ae��YC�G�.j�+�ҀK��ډFw�.M3���;�'�E���ծ��oVa~"8�U7����Osa����$th��R�R���q"�����H�4b� ����&guD���42&1�@�r�]H�`���U���#�%�ӜF��	�iu���S�Sla��2[Ɠ�� ��+�� ^�6�I��N�?.�h ^e�_��0tdO�4	gB뒈�{f�K��g\"H/hp�K-H����fx
��,K(�T�*�NH�wN�]��g5/�i6�B�=�x�AZ&� �Qı�|R��e�ԮK����G�HǼ�RX��4[7���X�lV��F
����y���ŸJ3���n��Ꞹ��n��ez�i���" ��˳�̻�ˉ*7������	"M
@:;�D���lVb��:=B��gI�e�+(�3���Lъ��	E����L�d(�C6�療�$3wO
�(TR��L����F�ŖT�u)����z�&��� {����S�բ+y�( ���P��>�e$ �����Ϛ1w������c��e �P[����ϾT�sF �K�^�)��Y%P�.Q|���		 �A�(���Z"%����c��&��5dsq��������#;W��z+��1��s�w_1a����oL���פn�V�;�X����R���$ڔ�k�E��2/������"�ȻLB	iǔ>LB��`2�S��L�̚�%� ��S▼%�^�I��E�<M�G�X�����0�����$����qs5�J��L8��E��0~�oY9��:��T�A����@�,�{C����&Q$�b�T���˜V��j=j��X�׵�?)� ����[����(Ig�QޮX����~�� lC�	��i��c�������0������8���vU��Μ�����K��eV	1�0�B�e�5Ɠa��tY�Dߦ#��C����Qs�23#yR���e�-���xG�0_u (U* �|''���X�8;r��e[`���SA�6�J!��\����NlI�ZA�g����b:EGl`�YO���J���ߚ}Pbd��<�׵�Nz��7FpA��<��B�i����ƪ!�Mi�I�~���r��݇rv�:/Ȩ�*�ƍ�4?ëx�$Xy�^a;}>ٖC�k%���%�o���;z̥ʿ(ڏ_m�H���Ȫ]�oY�mDԽh�	mFsx�B��6�|9z_C��\z�F*[,��	�yO�� ����i�?��B���{�G5ٿ��k#��X_�qy?e3C\3���o��^���^����cgf�JP]"$�:3� ����4.$G`A��zLOY���?�u����6R����K��/Oj�z�G¬�`�ت#��u,�is)6���C̾�"t�f�k�f~渟��A�w���X`l�nRL����і�VH��I6�g���1ꡳWa�.p�4_z7���ْ�)C��.?�b9cK!�Έ�H�����+����$�Y�9�{�y'Pz�Wd]�L���'���}�}��Ò��	�����"U�!9~G��ؚ~��8��Q-PD�4��!+\|�V�Q�K�tqv�Q`�45ޣ��W�Ƣ,�<�@>������x���\����͇�d��u�D�YL��r���*��f�d�̏�Z<Y=�*|�!��-��a�aĔ����c"�9]O��{�YP�j�i��AZb�B8_7�R|\H��-���FU� �b��%�a�e}�G��@��7��.4���;IYK5;]4�1V�(F]�[)��ғ[�X��]���=.j9S��<;XS�$(��#يXp\y;1Lj1zcZ��mm& ��^�P$�?p
��a�g����uPPJnI�-!C�p�O	-B��GѴ�͗�M�B��Ѯ_��m�A���J�[�kn�T�õ�Ni�"����=�
)����ۺ$��.���49�G�<���~Q�!Fr�l�z����[�z�Z�˳]��+w�Y;�X�����nG;&w�0��,U�7�ynRᜏ���/�����ï�O����bB���X���G���F�����]jY��̡�{�P��|���j��㈚ �݆�S�b�d_u�k�)��R���U�6<R�~h� �	��z�n����P;�� :�wBi��A�� �%���b�I���R�!�DP��W>�^ؗ��2 ��� �I54��z���p��ܮߡ
�D��Mow@+�"��q� ��D���Պ���,�����.��u�S�p^����1����8��3�����NʹX�I�24ZI<�kN�#$X�q��3$H���nՍ;K#u�?W�3������
`DH�\oGW��K��#1�ml��>Lg������6�"k=�!�`:�:[#'�".�aTΐ(z'��o��a�)t�31�E�E�"�̌��mK�Ǘ����<��;���X��.�_� q�0��љ�)�'?�0R0C�]I�yj��J�� =_V6{8O��,@i��~��ۻ�0B���0����:J�M�mw��<�����n$�6%���	����)^��f�1��eɺ� �{����z������K�)�:�0�sr�_D�*�;�&�����CV�w��"M��/O>ۍ{+�+vQy�v\����N�%��stc��	h���)�9D��-�d|. %'�LG����`�q����� ﶴI#��c֐�o�?��7�g�n�0����F8eFKl �FV�����]�G�l�>*2�Dh�z��P=2����R����6�{�H-����K���'-�>�A�t��,F��;J�s������׭d�!�/����$r�i��&�m��2��}�h�� ��* U���^W���<�s�ݽ����ʂ�U�yV����fo\>��jƛ�y^fb`�.kX{m�M�� ��$e��ҁD���1VT�י�-zU��"+�Q����W���e����h>&�6a2 'A6��0��R�o�~�J>S<a�%f�c��>l��YE��3Aß�`�Y��̙�G&�$�9քhm0�c���D�
-�h�čn@��/�̓��)�/�u-�c=��8:'�P�nj{�?d	��R����=�9��q�����p� ނ78Xo�T1���q�	���J�K,߃ j�j�O��頄���U^>�_B.WxԷ;���l�:��4h�"oyӌV���`�Ťy�9�� �N
�K��^4�ĜJ4�t�,��7�*g���qZA����;�8�����
__��>qnT�/�`�+� %�!��U�8�N+ʸ�6̮�?�#��~��~���������P����f"9����@}e�}"��R���I�X��` ����JԼ@̥P+]a��T��w���sԙ���K'��3�-�h߯������6�]9hdc`R�����o��b,Y�#��䠺s��f��b�4:�F��I>�h4�T�<���^FJ�s���3/�	��F�k�}�X�%��܏�T��D��;{|��#W}��ж�-� ®nI�V��2��W�bkX�c<�B\ꜳ1��S��;pS_Ɋ��l�Nr+��RE��/���s�����X�2���������+6�����n����� �gi|z�dČk[�Xmp��sF�4
l����ì�dv������~�������C��']8}�Ǖ~��P^V��UH>��]SPJ����K#fA:Wv_!uV�%��'�q�-V���g����W]�����h��W�!�A�"��vǸ���[+wn`z�v��q�J���GD�s�H�7 >���.TZx���_�Aû�
T�!�D�:�/�?4����}+����:�&�g*8�2�7
r�KH���miܒZ7�˰���E9I�����}	(�M��B ���6(\���R�B�4]�=�P1��r/M��2a�kcD��p�Ӈ�&�zי��gI,�]�����d�\-P�� rjw8�1�+}@ L�k���d��&���	Aዸ&���~��Sք�1	���L|a�i�u�brW�i�&s`�:]���w�xF�R(�,��2�����wK4�.��g���e��g�^�rw�̖$6�7�]��4�}iI�㚳R�&��7xQ�W��Aِ�ˤ�.a^��z�O��ƒ�ߌ��W�Ͻ��;E��?Zx�:��@��=��&����s�
�]�Bb�Ԝ������.a�Ju���d����$�'8���V���������9�
k��:�Қ�&W�������Q��6	G8_+�Z�-��E�H�"�I�J�J��?��ǅ����JZ]��	��/�:���N���/�m�b�+�|0�͒���c��?��� 4;�z���k�n����>���)	�0��lI=p�cR���)_�1��e]���.\ˤ�[
�@��\$�_�}ށ&�I�"+ݬ�Ij�7UZ�������\�����g6ut�Ϳ@�oW��������1%�h7�;��7��h"��?Ё"�!�a��$ٶ۵jg�S`R1��P(�6ve�����KLo;�`K>70nx���AcN�2��M��"��tS�cm�h�\.��@�Lcށ�ϼs�+¡�hˡĀP�<�f/�Y�<� %d�d��|�Df��ms��>�9�?	�l|�G����`ut�.;&������m��	��s4�T����!���B�˕�p5������y�Ah�H=��?NR��*�$}�=�3�44����EN��B�l�cɄ���o-kLY�3�y�F
/��}A�9��8Tm��77 D�D~�a�ȯxv1�8��>�0g'��n��v��.�V0�T6����>E�̭����}��/;�4k���収!��(����Z�:eLXUw=AF7�B�)IE�H��C��N�F��0�8������(f�'|��m�k���a�jϧȶ��v������(��xDؼ�[��kK�����2ކ=?;U8=W�	<'g,�/l�������"��"�+����B�����ߛo+�
+=7�3�m��s��@�u����2�b-�m��(�%kܺ���-��]n=��|	��g%\��G�pz/�^q�,d|@=V;�R�
\˔U	��d��5�Ir��H]l��!$�1�<���Jڿ�Jmi�ؐ���	u��#�j�p�qWy��������c�W��$�+��P	���&��},��9�^�䤩/��}���9�����ý4Z����;��ޛ� {��=���M�q3^�)Je2��[N���E��Lv
E�h�]���A�V�<9�_F*j|\*{�
��Q=��g9��@���q�́�x�R'~n>��J�o=)���@_�z�����ص���&g.y�p�_�{�� "��f.�����K�L$��dv~&E}!�E�`�U���A�4/O��`��!2��>�����h�#�(&�p`ӧ��/����vXI�0�8��j��<X�N#�F�j���Md>x���[ �V�����*�����|��(rP�қ�E灆o�D
�-+�߲��@߾Tݬ����d�K��
K�Te!N?"�#+�>��m�J��}�|ܻ��S��:;f{��M�K��]�U$�|���))V�� �@�R�`4�U���z��J�����pIv��ޟl��\&�:g�nS�"��I���2��
<��%��V�Of�0���2揟(�a/���}Pà����������y�J�ʭ����@�9{t70PM�Ҧ�4ԧ��-�G4��>y�n�{�c*q��ÅjO T�u��[̟��3�
'��kD���e�����	a�D8U-��~�`�WA<���C���~��c(��.8_�C�����>;J$4�����h*����Y�u(0>[�6��27r�X޲���9�$?��5�8���O;s�]
pXn˅1���rX�\��3��x���WQ��;�~��$���_�֕�Q�/�V���r|)d� W�8tD��>v}$�_��Cc�f����ٜ=�h�٨<���t�(��E�����/N�rEƦqv�^W�ަ/�*�����t��ӗ��]|rOM	�V-�/���|�!".�T32e��Vo�Q�y^��9��#�NZ�.饤����^G�x���jh����� ��:<���p�(��`|�?�qe~��`���s��'��gmvi���y��:�x)V{��y}S���G[�J��4����HaZƣ�~�=\��ǐ�	FFỄPԅ|�b�T8�M��e2,���ŖM�e,����I:�,O�t��hI�R��e�F��'$��Ij��lz��P\O�"�\>��e��Itj�h2BR�<ȃ��*�S�(d1h����o�ёp-��Z^���(Z������fg�w�����\/�(4ݾ2���^��bj�i�=�I}*��H:��vi���L�w��!��:N��vu"�(���)��[ƣ=)��u�7yyߣ����VO�'��$�A8��w(�>�:�4�4�%v�)J�08������Ł�i��(�7�)g
�+>9�
�ϭ���Z	.�))�za�ӈW7#E��wC���%��b��2��]��=�Li����8|���Z�B�>��N���,�jw����Oت���/ĦS]�9/uDI�M.������q�>����A�u�ʟ���,sW<�/��2Z�8֢73�m.�bc��y�c�J.��u�A���f\�DZ7%��צ�Ao���Ui�(*�m�QN/��en�7�s~`9s$��2�Wa��w�AGe����7~N���/1�bG9�:�R�w��G ~#���Y�*� ���j'�XQ��&�}Q?CRCm���.,�/Ui�=C�2�������VχOU��m�����t@�/�И�R*-Kÿ,\g��=)��ԝ�t�Y>��WۙJ��;j����%#פ�.�çj�2��<#���4L��'�oJ��UuK?1�X0RCفo�w��/G�CI1!e�`�֭�:����=Qę��5���H��)t;�6K��	�C;P�t���nR@k�/�y�8x��Ra�=�ʯ�GP\���S�,oC�P�̇aø�Q�H���0e�e��O.���%�\XF0[AthDN��gN�H+�����_��q���&�H-3�V�ؚ�0Z�=$BX	^uh�v�sԑK�
�9�QFZl����;�T+��ʀ��'�e;5֋�o'��K�rB5 ~�*����2�ͫ�����V�	a��X�A���J�����b�/��u��;qL���EF���`k���(/5R�P�q�*��
N ����4�T����s��)?��)�O?�`�ˋ�la1�3U��t����V�Х��9��	�^]lVvz:ֻ�B.!d�2ߞ/
��\�ǵ;�	������>Q���'
l���g���k_�<�a�)^�Ot��=m?y��Z��B�O1P�P��F$\]}$�H�q�h^Ĥ�Y\0�X�\�F6 ��Y�	
�GsX�<:�+�	!G���F|���