��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY&�O9�fǶj���{I?7H�?o�6i��nE�UƇ�ќښy�g�\�pĚ����P�h��/�n;47[NmHZ�������Ȥq�g�.E�k��o���Pe{�5��aY�ɢv���U��A�O�qx���Q�Ľ��~R�6�N
ϗw���	�׮lNA��I7o/F����Pѽ�ױ՗�?\�17]I훗h�b��$N��J,��y��������F��"^�*�T36�^TX�!��'����vBC_�Y`���Ls
�Ђ+|F{������F��L�� �	��z��[�n��W�i������C/���+����zXV��M�v'��l��+"��8��R�G$���u?5UY�$C?� �۽0��S^��9�]��`[�9�:.@#�D-�a\>�Kл�gL���@Ou�?�3];Z�]����]Q�?	f�i�Ƃ�`2�V+��|�&g��<��*Q���k��ćf�R�Ji���/x^B˥)���$H�!L���8���'0� {���;|E�X��T����;���t)��>~�
HL�Vֹ����DY~M�ieSa�%t����&;��-�.q%H��.V����UΔ���I�O�F�~wygUO/V��<����F���(1�9���
�z�4(	>������Lo7d���P#2R��!�]����7@ݠN�Ew�L�}_��M �Y3�U�A[�m�Z�S�bx����c�
�l��=G�ګ�#�pd��鲝E̦}?L?޴4A}�`������*��r��ʑ�;@R���$w�&:�{�A��ׅ�Z<�c<}�!)��P�"����Z=���[����9{?&�C�L���א Oj�L<iL$X�����:�|Q���0&�&���@��=R�b�i��#��ˍXȞ2��rH�-�$��_�N�p�����4��f������ږkҮ�e4r��H�
2���	�Ԣ��W3�t���	��Ի3�`� ���Q��&�x�)�p��k`�TOܼ]-���z|ŭ�s�ZR��%iC2��\���@����������ҍ�� ���'Zo]��QVS4�!��k�SLR��4�i�+�w���Y��d��q z|9ʸ�^����%8Ԩ� ࠤ:h©�x�t��K�+�J�p�>4�'VB�q +�|6���ص��s����`ȗʨ��	@��#\o(�݊��XW������Ҥ���<�]LD?��"��y���_������3����NLE��{�8�u����P#�O:F	o�z�.���*�|��"���$���-�#?`���d'䯹+4��;[<�p�+���ͽ��A$i!(�b>�˲���t�6����\��,;ȸ<FG��|ܱ��B�Ȭ뻉�������ߊ��p���1����P���1v��<�Yq_��9�r�?��B-�i�U��~����:����j�(��h�.�_4���'3m!	�.ra{�f{*e�S�=w��/����ㅜ.,���؀H�Q�Uz�=�8/}�Y����6k��{%��:���, m�	�0�>��*�P�J�m�$�:]����u�\cџ's݊Bg��V�To+m"E�XǑ�k<�s�r/�:��DeY!����.N�a��������(4�P��B*V=4s�mV�2*+?W>�$���MjY���6$#���M�7�WJ����OR��m�μ֩et�� 6D��$'٨�� ���=�Ժ��8����ֹ������ce�[ӌ��C6�S���%�^:rC�ь$5��D2�^�(' r6%�G��:��<،�����
I����'Jp����@��o=�N�.�����xĮ=�S����q�[�1i�!�@��mc[r��Ay�v`�sǲ�M�$b���\&r$z�,s���U��R�{�����E�N���!*4SD��v��u�i�l*���7]ξ�� ���Nͦ��Z��b �{����`���Mvr�Vs����tN��ں�QtD�Y��g�x�y2��H�_���%�Dq�Y��-�:�20	��n��}RC�/c-0Pz���s�I�D��3���tC�
��k����ڹ]}^�^�`	ݱ�����Q�
������ڎDU�91*�m4���EWF�Gr���尐�2�쿁�\��
G�&�o"�u'b�3g�OB�������$�w8��ڀ�[��!y<���a��rŨ�%G�`�L���k��s������ښؼ�<U1�Kw��� �.U�:��\�	���1��Tm�P���α�RJ!d'l�0���˦��A�nFc�>|ZܨB˵B,Vt�����~1�y�p/=�#�X�O���0���ds��Bq�PXri�<"o��@4`*^N	�|U�l�b�f�k@Ob���]�(h���~a��G��@a�gѯX�	Ubnڕ���I]@O�?�:\��.��sHӓHڵ�~=�}���a�X1A@^���Bim�?.}a�k-����(��yP��/�j��Z�6�|H�NCS�tzEk�1�?���-�"�k1@&Z�?��G;}1
�hl�ĎSn�g�E��N(BKH���3�!v^5 AE��'o���->5����܈��9�]�ޞ_5X(ǒ̋o���i��DaL���]�pl�{���~��X<�E,F��r�ãu�(>�$&�����y*-��t���/K���M��1��op�,����J��$#�¥yk�wv�u���\��k���QwH	}��l"@��RI�s	�7O-5�Nl"Q�5�C��.y��I䩰I�X��Ϡ��)BP�Ƞg��|���"�T�
��6bX-g�a�h;R���IQDd��=o'D�C�k&}������_���b���؁�vǸ��ǝ�6��ċ=Li �/�ܰ�Y��{��Z�b�Y���o��.�)T�!�bI�sN��ⵠb�[ߋ���X��٫J��� �.�b�IkF��T^�خ��:�_��(�R��Qq?����o�jC�S�{e��ɰ~��EڸE�2+�B��/%��'2xLɑ��C��8�π�b���FeE����F��jP�����׎T���廃��h�瑹������J��j[Y�?��S�3�	հ���#��O�(i���P{pHj�O>j�4���;��,�b��O�^W\���~d�h��'n4���Y���n���39@7�m�?9Ex����x�S����W�pp�h V������JGv{��	'�]Ԕ�/�����U�mN7��}�8yW��:m�--��&;ޚ��8���-lD�?��ᙸ������Gr� \�����b?�D�N(�Iq�`)���
���Bh�B9�w����	#g��* ����#_��!;7,~��7���������ZmHM<���6*����5?%��U ��r��TTex���G�)q8!�,�!���	]�4�7ݑ�c�����>���&��9HK��
���((Gf��z�����妐��'�U��K��Ȃ�����D������@���W�i��:b��ȧ��{l�Ԑ/ZGh�b=_"gȬ-VO�m;q$�ך��-m��!��ߛ�M��@�{A��)>aH�5Y�6Z�Le��h����Z���7qс���!9G�vx)t�	�>��{L�mAf�yb���6ֶ,$F�ܬ���w�9�f�M�?P�� ������=s�v�
��n���ރ?�w��c���%�j�$�&�ݧ`�
0�HO�y�]Q?�c
 �ls�@?�v]��qL�mzsP�����#��f����cv�u�z=�� p��B��\$�~�jT� cV�Lw*j��KM�PA�wx����jM��m^7
�l*H���V-�xXt�j̓�R	_DԌ{yR!�Da-
��@�v ��t'��� B�$o�񂃑x.��hzL�L�#)�e�})u�Z���>R���nI�08�zM>q��	��tXi��2�����@?��X�n4�+�+�K�1�1vE�Q:jm�`�c�C_vC�Y��]"����f(� ��
t;���)�_(�DDj� �Lכ9O��'�����@�m���&��B���K��e����j7�16��R�33���pu�0Z�������d��U�-��l�j���Pz������z#�f�L:��ҳ6ea���an�gc�.p C����Bm�<��0^7m��ؙF�믾\�<+̶��zh5~�ʽofJ�[�U��b&":��Q������ �eh����'ۛf��\�����Iˮ��!�J�t�9 }�/���^34��P��3>��
e������.��)J#J٥�jK|��B6�i
{��";���~�S`73f7˃O{��(�/�8�}�X���Yj#�� C����hh��������(��qDe����g7����΢�#��?���A�h�7Z_f�5����� �>d� �z�{���	�`���,�D�n�5a~#�I������Q�]�n��&���Zӭ-䀹`�&#���BJ���ֈ�YG�ʚ�K�/$��&�ʗ9|�8�j?y�yLL������㟐�`IK�|�U�G1s�~gn����?Ae(�5���Ϯ+��I#'|�W��,���K,��q��٬RK��]{�<*, Nĭ�E�wW�^��C��:���;)�/�A�9�~_Q���pP����_�~R���]h�(tߘ���Z*���:�O�xy:!���ߍ�l�(,�~ǋ(�]����)�&sH�F����:�R� F�0Ψa��ܰ"`��w�H�(CO�yȓ3��V��+�Rm�N�r޻��}L�t�.�챂����d���/ߣH1Z!�7���o�A����Uzv��D�z�If��7w�#n�7�����5�Ն��>Ó+��elrMm$R��rw�&#[�lj��{C�t(A1,	%�{��,���IUd�ڔ�i��p�ޫ]QÛ�B�Ep���ʉ/̹����,�B��r5@F�K4K��K��<���MF�E�'G�'1bf:��@�u�`e��j*��#A8<�h.]��i������	�O�����EF:Q4�9!��N�����C���+��o����Eؓȏ��ˠ���C�6�ɩ�}�bhN��V]4��A��9c	�8�t�ۼ�W=7Y��w���^YF��RH\����M���w��P8�}�P<�7��2����1|�_���O�����q��jq�2�^�1i@�b�U�����٫�nr��?���6���*#�B�c��7נMA��%�"�_�t�£Q7V�}nJ��B�Ey�ֆ�pQ�e���rw����G�$6qTٶ<������^�ŀ��Y��-��}!���X�y�?hN���f��hӨ*���ڜ`����R�y�*3�#�V����!����%)D!�v�TiSC���)����$L����[,�y���9��\GXZ0!��0��א'�&�2�eZ1�$m���� #��:����xd�0Ax�k�U|��ب$���N�7����jR�7c��rw�R����Ѻ
�b;�]˗T��'�=ߺ�e�Îh�z!Od�Fj�z�FZ!k����ӛ��W�R����u���Z�tM4�_¢�Y	.f��e}�MhnH)]<��D���*������?O�ٜ�@}y@�YsAH��ɂQE��W��Q�{Z�J��;���+�+�V���_�1���Ҩ���4�Y��Ii����S��35���d��������|����veT#�ce�.��9\��ѡ���_cd�`��?��;qL1Z���EhBν�j'�K�j���e�V�U�AA)��!�B*����@{�vX���Q`�(�M��.�����TMg�h�딲'_�"8�q�W���̵�7��[?@����w[���g9�;��⒄�	2��i���Rڋ����V����<@�;��R�S�O+30֩�|efF����*9�r���	�@���>D�Q�G��<��,{�򳝚$�<�Z/f��|P&� 8�fPt�dd��$� �f~��{'�)�WR��H�q CV����V;p���Z}R�H$���`��Ou�)=d,�@������OL9���l�p28��o|��l{2md������0 >�wJ�*���[��j�9c�^|E�Vo2u-j���� am��NnάY�/B8&e%�w�vp�P�TF��)z8�{����q۾9�������@����3�f6ˊKE���qZL�i9�M�ߏ��l2�B��Ԩ��o�	�q�� $8���(��lW�8����=�p9�vRjτP8�֘�.�"�o
������B�^h}i}W�՛Z4AAD��Q�r�����S	���Ŧu�6����Zz	\���f55��Y��m�?���{ 4u�Tqn�c���q�
.��Ui������P�-�����+pL�S`K Ba�nrZA��Œ|_w3)�K����(���'�ME6�v�u�%#}���q���b�KF1�N(�GS�?���&��/y�_HɃ�!Z}���t�7F~�����Iֽ6�.����H��F3P�vI��ٜg���9�e��p�2�91�0k2�i�G�0ز�-���\w�ߥc�t�XT���1����?��e������fc5��;�ͱ���#>�Y�`���C��f������'�8/�� �Y^�[�Tx�U�y>:U_Ùu:�9��V�4�&�>n�*"�fn�4W\vF�X8��_��!��)�����"!�}���DB'(��l�۵?�JQ��/�[n��#'P
�A g��
�D��u �H4�d�E���7ҙ�2��W��\�EF��D縜�$�B w����T˅H�=��HQ��x�W�hTU��i����]Z����Iw�]5�S�x>=�6��W��]�LDF'�rf�bֿf����d�0�\eR(���n�x�sg6����P#,Jy����%����y��j�,��I��X�7*�E'��S0L�O�����KpI�� ł_�h�����e�+��"!g�e�o�������<}�ج���[���2�¨� ��Y�ōK��2�����|�<N��y�(bjf�����xmm�_s��ӓ�3�rڝ��(�5̽2b:G�A[\d�ϵ՘�����*�+S�5�wD4}�(�&�)�`�Թ	#�a�3��hηf���i���á�B�֑�yߦ��`/�60��'�/�̗��:��_w&u˞S a��n�k�9 h2�PS�9t��V��H�1�܅���"��y�ɂ�{�`��Yֆ[d݄�wR��S D�AH�HL}1z0D�i����p&�FN�SZwT��3�����4���J��`�g���q�W���j�j�-+�D&^���B�#��p����L�e���xi���Y'�N���,��8�ba	��=Bf��� 	]���KOnG��CC�衡�Nٱ�C���s�$~G+��5�cTVIƿ$�.I���j�����
��ِrs�f�r(v��	�
:oD����o�=:{����k+�z�t�r`<���|eĞ
2�d���-�!,�+�E� �ڰ�Q̆2m�ѓ<6�&��m�G�/x��6E���ӄ�U�Lw8 �^X��H?���~4��e�.ڱL,����^��������4ZPaP���� iӨ���߈��|����"�l�oH1~�=�/Io��*�O)����o��+�6�[,�i��a��z�xj�3WHI"���P�~347��������ɻ�z�܏'�$�F�1ɟW��Ԏ��~��k�mE�����t�~q�YKn�.�5�x��il�iEM��{Y��ދeS�\�`.�Z�����XVRT���Ժ��������l��~>}Ԟ�L�J���� �S��U#^I�P?(Q���%X� ���n��B{.�</�lF��"�ܱ2w��|���΃�I|/x���1�=\���{���T �U���m,�TIx�#��Ϧ�$��s���|��j���[�&	�����e��c���A�z-����Ik��ͯRP@r��y���C�gy�c_u�͞�]�zM_W��{��Jq7T�Cl��Ge�|��!Ng�����Pv:s���1�sˇ��m~ (z���q|�j'�	Q��� V��#�&��hH�v �k* к��g%m��X;_6��wV<x��nB
>��q�ʟ�'l�OcXE���LM�(�0�(_�!���0�w�1:H0�Q9? Z��>����U�e�yã����g�?m�k��;��I�EZ�)���,[�|i�N�5&;�M�&�g�>���=4O�V�hrY�G�۷��?\C���E+�%ు��˥���U��(SE8-����X�4�y��r�		L�޿���)���_��u���n�/�?Zk�@�tcs�s�`�ԓ爧~l����0��t�-���������e (�5dv%[��LA+�+�-���y���p���HpXM˲x�T
)��#a�M�1�6��-�������$}@�("��$θb�jp���/M���#��ؼ��5�$�7�:�G'����4��sxџ��8�91���֭��31�$:���d;6֭�/����͒UK��=�4�i�p�W�[x5��BSw� ͩč!�n�8�t�+,�������Z%*p�k�:�<F6���Ru6:g�:���/���)��z>a/o).~,8~%���}�lP�R��f��i�V� ��X��I2Ox�\Al@m@�a�+�7{l��(Y����gs
.�34cW0�0>ƉtD!S@�t �Gj,���{��s?W5&}��W�X�r�Y�����Yk���֩Q0�u�(~�Q,@>p�R:J%����h:��_տ��d�/S�"T̿�,�����d�J�i��8�l��`�0Jm!��k��,�X�Ү[��M���ܕ�����uc�"���v��5b9;�6������R�9��Ͱ��K��m���*�VAJ�o!��[�Z/}��*�3�B|��^B`�@0z����"b��i�E��5��g��`�XL2c�J9W�cز}c�8�q�ܧ�9?LΗ%�8f#I$�kb�$�$�D��6/��α���A:m������Is�vFh�oxP��y�=6�'�]���<�-i���n���1Mª�.�uv:�����E\�RQ����0xx/ĻH`��������gZ�Ј=!��X��{_�w-dh��C�1��q�������$p)g�XO��dY���W���X �u�����[���6�ƊӬU���I���sf��P�*2��C�\i��O���a�lT/��sA��_����;ܱ�T{N	kv����;�&��g��SY�/SM�����c C1�v��!�����z%�f"2ĿT�/��x�`����'ۆɴ,��D��f��ҡ�~���h����aғ9ƒ��\Y�MW�LZez��`��d���q^�1p��Uȫ3���{��#-T�CU ��I��R�=�ӕ�Q��;Z�?���a�-���q9�ڱs��w97����hY��<�$��j�7�������S�n;�yD姥k΅T���ɱ>�qJu%����b`��P�	�����2$��Ddg�ѧG`d�3,%�|^F	�$�z����s�jS~z�ύ.��|����@�ݑ��8��5`Uj�����M-�HQa<��� #/$&�5}�$��q9����Z���@*˂C�J)u����Oť�Iu���>u���	�	��>q��������9����@,t���� 'v�r�di���"G����=�N�0�S�;�%Ĭ$�E�C�o���q��m��D��l�� ~���+'F�	�a
R�����H<!�Q�,P��uQA��7(�8ө7�Z�ͫV�x�PI���ΧR3�r���Rp��L�?h�J����a�s�,nW}R�p����b��#��^�/E0WY�ɽ�%u�=������n�!v꼒���-ߔIqq;���hc�!��s�'@���7P��#�oM�M�E=���������I��t�� � $'ڬV	(��b�8����9ѩT�褞�$���q6E�n�����7��5��^���`�G�C��#x��˷R��b��>S��Uݭ"�-�4(����[W\+��ˊi[J�ns<��q��m >������^��5&	��V0��O��c�A��J�*�r��H���'Tx���`58G��z�=:��ҿ}�S�b;)��@5�Wܖ䵧(���Ԉ����F_��x]��+��������!�s���дn�x�N2��9��)�`�F�ć�""�=t�'C#�X���2:��˟�Q���
���cLY��>4����&�c��mG�o�'����a[L�u�����'72�:p����0K��&5�F�ߪkq�Ӳ�G��>ba8/����=&m����x��� �� Uk���4{
Y�}���~����o�����-��̼�X1��j�N���1�9"��+�{�l��Ȱ֨X�-�?_��PX��c��#�v�ﺂ�|�W�W�� �\h�֮�"Hkրg<�:�,6:7Ku0?�٫���8/�������7)�+���H�}0*R��A<�#f���T1�8�G��%�}�tzI}@P��� �5j9<r��� �{��߹m37��Ӵ>�I��wUk|,ኆ���NU�aNP.�Y4�l@%15Xj qV�o�%v�V�7�7E��UP��2�]�G��[
%�Ѥ�ǧ��G��,�����=c�^�^��YT1�x*�N� �_�7F�ls�����ԑ2n�3gjs�-	�'Ѽ�{��`���9�,�W�u�:��Q���5���
�M�p^dm��,�LF{�1����%��c����4F���A����CX&h��w��2���ּM�\��R�}WtkA�2�6�~a!�H[�Cvį��;nZU)'��\2�l@��CB{�e�C�*������}����?���4o$s`٤q�3��X�9����5�,�ꆪ�)����C�\7ui�S2a�M��P�x�8�&Co+َ��\p��o�Î�U-,�����&+2:�߆��5T���<*�r�j��'O�-sؗ���F�N��,�X�~ӓ��y�0���f�#W����p�i��:S�B�]*JR�����ʀ���U�?1`/��:�=I���t�C�d��+�=9ϘJ����,��v��=<熰z����M�nk��wH ��?��������⏫K��2!ԼJ�N�g�F�(�9U�[V'�rB���"U���n^���,��yT��:����(�S��
e�.��T��̓^�_� �a¬-2CU�0$��﹖�=rY̹#L-�� �w�g�d��-b;&s�|Uē5I5�OA���BY݄��A������T���9RьUnX[-�|
r�U�����F`�g�La�х��zZ���闡�ǝ�օ���}��^��r��]���$����ݚ*� %���	�N�	'�[���	��^�l1�?/�p/�ec��s�#'}sx�}V�s!�A�y�9����@��|{��b!�	�¾;N���/��Wv���.m#3����L�V#�#=ҫ�����x�I�<t�ZT=|CɨT�n��;0��p��	\}��0M��v�9����&�<N9{rid�r4E�L����1֩��:��^�����#�6K4��c*���F�oL�w��L���[�m����^�N��k��j�X��-[@����8��;�Y��{	:cD�ay�oS��|E"Yb;���v�Xz��f?5���;��t��Z�C¹�򒨝��,e��HP��!��mb�ג>ó������A+��Lz썎'ŷː�3���/ ����a�0(��.Ř�{�����$!PxSy+t�mǖ�B^�'3�d�������̤�g(�cMV���-Ҹ8g��7��׾���b���Y��}a�wC���G��48� ]��hqQ)EC�&B��{ ��{j��u�8����j�.�#91#���)�I�i�Fcw�?g�$�Ʈ��z��`����4~�9���X��{儳y�P_����+w�.I򽪙�jr�4ɮ�'�;��:�!DS���[� Sl��!I3Wt���'@.5���B��66P��O�cP�	�y��o ܁s�D�����6�p��ύ�`B��_!����e�`jՆv�U�Y�:�^0��rҖAI	�iM�CF6�$��=��*����cp�\��>�F����{��7fi)��+.�9n��>��t�l�9��i�,�g^G�F�\A�	�YB�7���+�g.�F_0T}o\�4^�Rv�O�*:�:�8 ��nZKg�� مJ+#�-�??�)�`�!����僵��-�DO��3�}��Z�bVi˕��j*th-�Պǧ��\@IOK�q(���?�l�B��@Ť����WҦyW�׎r��Í'fw$�Yp~4�y��|	)e���/��(`c��~hf�f��w�XfV���]b�%~��Q�x� e�2
\Y��H~�� �1�d�O���%"@�2Z:��ga��IY�_��~���w�s��6�~$(�k��];G�S�w�&��J���%K��%��Z�|�� �����e�����-�ǫ�tl�D� {*�X��b�jnJ��O��A�� "�����Ճ��U|���Ү���>��u> \�;ý��ݠ�R�i�]*�Y�(�=����A�a2x��	�m��,�W�/z��mѥ`	_B�p�s;�N�z��I��\�k�U��-�l��3�w~�sq�N6�,:rٯ>�L|��#�6dxCD���2_��_�D�������7m�9�]X$R�����!�l���K�i�h&�b�*��Ӊ����Ɨ��[�X�;e�
>S�L�\��z�W�u���Y�_�q~J'�Z0�5�P ���u�{�K���s���\V��ٓ��m(��r�U�)��w��9�Vtb�@�p��D�9��R�C�����&�PF�F%Tev߹Ro:��^��<�����u��!@�R^!s��]��rڵ�,�q��+�1�qk��£��$s n6�"�O�"�k�1����?cB�c���,��t�if�����iݠ��n��f
?���4�k��5ĳ�V��CRL:�e7UDO�y�}�qgb��E������3���tS~��Mv���ʽi\(���!�o�OyTΝ��*�/�H����P�foPQ����h玭�T����A���H�����}ľ�����6�ޯd��Bl�η���g���Z�x�ְ�f��m��T6�[�IA�|�lk�W���v���u�㾫��T{1tהI�jӌr�\r��zC��85���A�g�Ab�]I|=V�OJ���c�O�\�1� &rTT5��I�$l�h<����ڙ	-R��d�̻NiW��l�-�����s,A��Q�Bsˋ6{u�ר�����iHh��D� :���\
�*|�)�f��>Q�c'e5��S�v3��}�\]�Y�t�Y�O@�����[���t[����ҹ�o�a!%����%w��V��n�KO���ӯ4�ڔN��'�>�K�t�p{\l���ɉ�� >�&(̱@Aa�����6�%���NQ�F��)t'�6;ҫS��;���e�j�S8U�P�l��b�s��M�02!kf�]�TF��̀�z���#6�޶Sf�-gx���[WT%�<K��i�X4fۚv��7^�秓V?eZ�6�@���T�I!%���\�Q
�v��uŨ=�=%
QsQ��.�
nX�����z�p\�Z�S����G�vCY�}�+��Zoǫ,������3�C-���p��u�x�bO��A��ǥa����J�fd�HȃO�]���ˣ��+�J,���[����f��� �O+�����No79��2]_w#�k���;3>�C\��m)#�S��X�Ꮘ%غ�-��p��C�l5������yf/*��kU] L����5��\߅�K1=��<?��S�^��5I��?s��0��"��_��\��)c�jU&R�T�L	�?4{�^-J��SDY���-]��ٱE��J�W֫<�Y�Ë�y{���G���9�����Nc��q@eۍ�tЂ���Mzh�{z�7��Gâ���e����ңfϭEUa�d��)6�D�23����7��3H��b
��e�]��,�\�� �%�?��vxmz�K�?nM��䚇��8���7* ��_�w�T�PF��j��W�MSC���^�%e�|�xt�@>��f!�s?R�ճ^So���PBoN�,`A#)%�����זh�������-N�Ժ�M�B�/��{Jlq��g���=�.����=4�u	ے�b�g��r��L�����z 8�i�˔�a$�/
� �T��r� ���;o{�X��� ��/�d�0*��'��|�i�,ˍ=)�η���5��Z���2��E�4��������+�ɜ+O��P��q�!g�=�t�(n���%t��ߕ5��[+�=�5v��v��Tx�]S�!mD�R%��y��
��e�`�æ�0�H͟�t�����H/�f��CJ�MM{N��}�)�|{��TD�}��`Fw�%x�1�xx�f(n;���[
�(��W_z��Y��g��xn���ar{��S�M���ي��X�������.�aeQء��!hl�	���lt��\%�ۡ���CC1�̃"V�9;�}�q�SD��u�.�� &|�V��n��׸�K�DB�0��\��J��QS=ѻ�"4��ّ�'\�[H�n���@Y��?x��,��δ�g>ɂ��2���qڊ�?���ݕ��b�w�W&��w����zʌ�w-���  o$
b=�����5Ffa �7Lm�'߬���쎂��Q����2f��efh����L�5�
"�tM>�~ŉO}��&�YЊ����,ȟ2�t�Ri�[�ĕv��8��)�f�؏H_�� 8 ��n1�gE�3UƼ�R��)�ei'����Q�:����E9Q�ԋ�G��3�s�(�Dɏ��-Aek��%-SB�y�썻弽�_�X��u2K;�X�W�h�-�A�����`�	��a�fFpQ+w��l�\�p6��ʠ�[y�K9;w]�����<�R��T�b�S�Xe F����0l��Sr��ͅI�T���c7g�8��Wƚ�å8����Mʃ�G�{�{Ǳ��|J]׺~<�]b?�bxQ�2yF��^+EIM����d� �S�m�w�12�,�����h��&q�M"ԅ�tH7�fϥ��H�\6���+����N�*�py
��&��j)	��~"�.� c���(�SbN���a�b<�J�D��Z���6I�
0�Ú7�k��zM��=�2�#�F�N��Ǟa&"g�xr�N�zm�9���<7̱`]�/׺�y�;^�*��;�Ab���Jb&WR�UQ怓��&�,�&���Ҧ���ι�,Ze�
��w+W��Q��ql�R���LPV�<�L�I�-ʅ��'�$�'��QC�'�f�g�2���ic����؝�
{BTS&7�O��4�/Dl���1�+���w�&ڀ�R�i�(-0���y�B� ,#�.<οs�q���(��X�-#X��Cį�ߪ︤��!��L�?P�M���@1��0��UZ��{�J�<����M���O�LQh�$�����b�e����~BR����R\u+�s�?�Y3pxYo �oc�QE��(5?
`k�����1?�,riD\ĳe���ox%�8�H>༳�$�GB�����\��S�T�D͜(��"sK��t���P�����O�4��bb;��v�L,	�ڑ
���[�(��"�����tk�0Y�^^²mc���f�ya���E��bZ	c�f��?�(:������G�������} ��1q����}���r�-Uѓϑ�� �a���E"3Z�Mu͒�Xb9�y�s4����+сF:ҥ�,��d{|���8a�uv)��K6��eODp]�_f�C�uQeŕԐ���C��0,�>ؿb
/�IqG�=R�V�c�9s�v��L~z�u=Y"9��:c����.�OP4_�lt����|��M"�G�� 	��f�1���$l��.*矓�+(�F�Sٝq�?�_�JGK9�,6^ϸ��?��Qi��颚��d+�w���Z�C.誺��ҏ�(b#�ƀ�`�w��������֪O�y�82�36/��"��P�;�����u�t��g�FΙ�@4��0�.��Z>5O!l.'��*�޲}u�ɍ��rͷCZ���d�楯6X��k��省WM���li�����V��ۄ.��83�C��>ғf��	W{$�.]Za��l�2�i/����?�8GƖ��X��pPȂ�ٕ�d�x�κ�Ř�,���l!�����+�؉��Uj4��(��@��'�JԱ9�����Q����p`I�B��j�`�xi3��-c���_�Y�� ޳�q�Y9��;�(����>��mY�DT���h��b̘0��שּ���<L����"{���<j�a�-_,�C��
�Val�o�)��+�m���-Q��Ӎ���`ͅm`�!"�U4e������CV㝩��d���#n�@�P�yԬ��;x�B̥�Z�4ޡ�W��5"^�,|�ϳ�n�z"M�>Kw=��M3d0"�5��"��j	AH�XJ�!&h�7��o��T�� �sw�:4�_#��K���٩�ෘ͖%CIZq+ż|9�����9�}?�C��]��V7�v-��R�مq�0��������<����I�҂����E�C�yKP����ި�oU�DyĶԏ"�Ԕq��J�Fb�il*���?�2��x��"A=EF�o�.zgH���ҳ��~�`2X���O�W���rS�����}����"�ʄ��i9>9��ֵ�6~>�e��#8 �9h9�?X�{��z��p�Y�������Bӆ(H?��>�����k-h�ܧ�Ens�Wˢ"m��Mu��T�<�r۱�J�>$���Hoe+���t;i:R��S��Q(j����=��L�

/Q̴5T	R�a�"��~�#i]��u,i����خ�[B��̄�;Xw/�xMޖ��r����aW�ZGw�hY���4���b����56(������weh�r��Q��3ֿ��6�m���lmmx�z�݈�z����~�	�{�s׊�ru�����l��Hġ���|Sα��^[�_M��u�������Ĉ��\,E'l�6
�R��kt�X�d�-�1=�U�������\o�����^���!imw'̒^@ÌN�`1�/���=��E&E㧳��P�觉��~{����G҂�,|�	E�B�3�7�Ұ��1<b2`jzrn/�9�3��^���.�26ύ�5�:��O�c���{��n޳���$S]3��ATX�7x�ѭ�J6Kf�Kp4�74S%���#���}�dmQ�S!���|/�"X˛9U���m�uk�����@�/��Q/����97OI���ju����SJP�KC��X�?^��cqo�`�&G=/�S�FzL�]hb	�0 �ְg�|A1|��ӽ�����Bӆ�)�U�����%0ĥ{GgC ���ì;<X1�k1�2x�6�yݡ�?8�k�5�%�K�~�)#lo�f�c�Z%X\���So��0����������7R5�r�r�g��SZ-���b�W�t���!b�W$�����!ٯ�ej0��5�6�8�q
\3b�ȇg�cD�F�F�J&6�)���B�Ȼ���q��VO3�aL�K:�2�:����Vs���i��_|~ͯ���0�p���kU�NB����=r�z���!R��Xw��=��_����馝,ΰ��M�l]�1��U����~�ې�2��eGuq8]32q0,��!N�lk�3~s��Џ}�P�`{ujů$�f�h���@���#`h���i���Z�谳�-J/׫M�X�{�8@�2��{ʴm��lp�� ў�3z�C�n~�.⟈���~Sg}+<'�1��^!��Ƒ����$v��(c���0�>pH���Y�<	��ښ�$ƇU�"M��lHlkzT��}��Y�R���%�{XX{ �X�I�]�u����b*��e�`&(�����qV�Nń�q��v܉��)1���x�P�7cCA��0�.�8�˥A��E�(�� 	��m(p��)�ŕ��B|�#G%�O$��&�̇���4<9�-2�g��������ނ��6��l��2�E<����%X�{R�\x�2lZ�N���P�<�̠7}�����M�^HB���l�_ˍR��57]̪���T(���T����̸l=X�D�;;P���Bف���S��J��?�m�5�PL ;yb6���B����ȍ�S� lb1�>��f�{6�yi�Q�&V��Ck"�G�WEh�՟w�@X��(��~�J%�!^{�����U�����N)&�~H��-a2���QՔc�k� .|��.��'���D��{�d*�O��C<ǋ\)�V~Gѷ��B�T�SC\�'-y����$�ct��&��ҥ� �;�v�|3��+�Nu��J�U#�f��D���[��:.Ă&��W���MƇ�f~R�⊴�Db�(yx`;�K%��U���ofn�g��	���X�.% �ī����,7��~V٬sVU���D@O��Ѽ�F�T��ؿ�i��?OW~�����Ԋb��bY�9N���[�Ǎ,�����wh���{��@�ST=�<�rL��wwu$��Mkd���@E� �D��	�-�Nͅ�����]Y�c?��~��*��_H@�m��>@1M���)B�T-�o�|NصO=�k߁&�����H�?w��A�m�Ϣ�C� W̨f1-��s�O6�i|��i���H��8�(.=C=����	�G�#o��r�����(����ZrʶpȸH2��RZN@'���`�Y���`�))a�fTq'�Xg��O�	�0 �۾��{���#-y�����`�����/�����U
�W��T>�V
֩W.ņ��b���J�
'Ϻ$EB�a��a�v.��z��$�����IܿW�J�7U�1�_�LL�Z��.�Ք�I��>&����!�=9I�N�� �}�sL<�bM��n"�{n2V�~{����U����1ߖ׽
=w˦P0�@hh���M�Lazx��>����;t��h�~�sf�`��6��*�F��x�7|��O�wYeM�O�1�7�vzs�ȍL��o��(ՙT8�^RM��*B�g)P:��V��4��)����Gd=�_��S�rF�e����6E	;M4d���h�Å�K�1`���+�e����·H�J�]}�زx�q�P:	X+����<��6K�:��ACp��b>'�ٙ]Zz���[����{1�F4�jͺ�_�L�hL[�g��k����@'��o&��;(h|�DY�����4h� ��o�D�3�d��7���R4�� ��>ץ�NEv���w�L��SH^09S����J�b/%�֔��:t�c|��M�"0���l�6�uP��x�i�N;)���΄�u:���6�C1(�+39`4'�ް�:�8��/Eoqp�8s����t%�c5���)�m��R
y��=�*o��𕟤���o�����|݁1��TS�R��dwq���k|��,6b5�ehB�DN�K�l�2J��g G�1l��`n�K�/�>6hK�37�M^-���9!m�l��U_�P?�2��%Qhp'D��_�63����گ�;�q�x!�kH��ǐT��o�c ���d}�M��CUA��>�I�^u͖��yV��o�}/�3�*����-]W*�.�N5�I�`��(Ϗ�
KȷF���X�C�ٸ��x���B %D�'�{Η�c9���g�w�+�(�ѽ�-Lt� ��H�L�͘~#�Uʮ�p��Y:
��ޮ'�F��Vj3R��>%�����4����+�b�s�}�� �3|���4s+�?��ᩬ�fi_���ⅅ4>1!)����Q<m��8L�t��KBo��A��K&�B�`yZ�I�zXdћ��|�I̴�z�Nx�;��w�������,���+^'����&�24N�A}{�1�C�9gGU������ef���\h��Eg���3m��v1fZr���K������,R)�<�ϒ�J�yA����6X33����2K�b���h4���,#7*ڮ2���Y�5R{�0o4 gp}�d��M�Ko�iNM��?5|:y#�6w�8`�^��H��.0��O�N��Dx�G��r��{����(R�I�ay�;���i-����_1sP���{�/AR�TH�%�4ڷ$v������s��C��c��	ͩJt����p`?��a~(n���$�jN����4�ϨP3�q}\��
���6� .]���u�ބu���Ԫ�D�����m\%M$���1�dU����كn0Z���ڙ�e{�O+�#Ω�ӈJV���SLi|��&�n>����:�P���eX�V�%������h���,z�7�����R�W�?�-E�}~1r�[ �h�h��j"�1ͷ�|(7�3�U��6��a�ˋ�|����~�o�i�(��G�������Rn/�+���Rٮ��]�}Y�3�i��P���;cݠ�pZ�舄7���ʿ^扈������}[���R�ϙr�j� ��O.�d��h>�MR�B�m#�y�#��-8e6�_�PV�A,X���U�8�˷���a��m�5,0)�@�$/Ϭ�2`ţϱ ��R�bE��B���,gg������k�Zo!�</�Ɣ�/G��9]VI��ߏN�K� ��$s�k�[���&�F�ȱ+>�9K�N��Q'����(�E��n`��S��?I�ǿE1U���f5߇� �4�#7?�gM��U�\�egKW�v���|5�h��Q��7	,`����\��$Z�6R W0�Pܳi���q���Y먐��T�%��������蜸m��~��`5jSTk���lk{������@�On�Ì���싪�d�<T(!'�.�AȒ�H�3oh���q։�M��XADnU֛�ݱ��pS�>�U�Nt{�l�T;'�<%�%v�J�f�g��f��h��߿�;������A/�L�K���r,�v*���[ �[h���}(���D����N��}������>m!��zפ����Q�S8�Ʀ6��;O�{���n���Ȇ����������3S����Naq2��fuu&)�<�Jp*ͩE�����u��~?�H8�l����g�<���J�<i�yz8G��%�A�3\Ã�z�s�,���nc"�AqSO&і��Ʌ��	ؑ	�A/����B�3�Go��2YD.��^b�;��9ؔ�!�x�>aJ�"�� �`(N�9�t{?ҠaQ�Us���XR�t5L��<SJ��L��L��X �q�����I�)!b7���]%�ۂ����N�7n�{��⚏W��Ə7�p���s֝ghyݾ�t�R��3DJ���;J�^������:A������k��
�Ɏ͚@�T��usN��� ��N�&(:����è�4+�
�U����������M�$¾䵹��fd���kvc�(�.�C��X9R�J��k��w؝A��M{�rUn�^��8���wAJ�"�Y=���zx����/���f��/)T03��	q-���:�H��ۈ�BZ�B�$	@�9We�&��d��߉0��vB3eQ�1ߦ��p�� Go��nGrV��4}��f�Ӓ؝��k&�5���bVݦ�kZ�,	�����>}��)�Ë��*=y?M/���C��1z��f��)�p@����"�/��\�v��bӎ�ީ����++z���zw�����6&C���	�b)f�����A��68��;�� �M�N�A��ݟ������o�U�[J��ϱ�z���Z��j��:v.�S�K��&|J>�W�l5�[��m4��T�+�ۊ��I}�_�bj�x�T����H��L�� d��)[q����}7���M_�Px��С��V	���2g�S�6��왵33y����4�^_��ݙ�i�cO���l���=�Cy�Ǧ��afW�W�1�g�τ�/�f]B+g�!b���?��iZ}^]�6��K��5���:��~��.G��F�[�
}�pbf�#-�H^�ʸ�l��
9y�&^8�H��͸ �a鵝�ݠ;�r��_��Jh7�� �`�����-��y��|�p��U������{7F}a5̫g�MD����'>�����Z��B���*0�>��!���z��z����Z��u]ǅ�`Ry��F�#$����s��m���������"	��a���5i����=6�"P������iq<�]����i�M���J;b�`*��\S�@�(�_|()Ȥ�㎯�dd�Fks��^KS���!�L����������O���E~��O3�nPZ��m� ~���YVzlm�r��¤>
�5�v&J�4�S0{c�#ogA�������F��0����%�&C��C������>�2�ѿ6>* '��Y�H�JO�����w�dYR�R�=X�7�JxH�S�/L�#7�B�ɵl��AA^��>�=��z�彅��ݛ�y��9�Q���:�YN:����6��=!�'h�K�b��{2i/T�eG��n����oqv�Z|Q�Ԭͳ��쉬}\>}| ���t�_N٧u��������&^4"�{<�=X�7os�#��"{<<�X��k��F7��m��&<P�0'�5[rm�ʍ�D}��jԖAa���O�ʢ �7`R3���g�v��5�^& ��YN��� =�S��V
��e���y-�s��������D�C�e1�����L���d�?&��	T*V�1�x�J��osUh�)���ץ��aϑa�愧
BJE2;�A�H�@vR�x�?p[��'UnDq����p]G״Hq$�9�����i/�ДI���_p7���vI��ҤXf��`T4O�3/#Q.ͬt���ųݿ�z��L7���B6L-p�9�)]%�/-��-|*lՓmRvn�S>,�p�<���J;��۬]��V�z���y�8��b�lN�"\���q����eҀRs�k�c��ld�rgna�6��o|FxƅgU,�\r�{�R*� ��A �Uם�X)����S�dfT0Nm��Z�\�*���Lѝ��\��7P��yĘqm$'o/u�����8��f�;z�L>G����(��2��[�d��Y�����K9}�"k�h8y$�1�FҼH:vM��������7�Ֆ�s���j����g�K�S�0�:C^��b��b2��1�6�K���옯���,6��VYQ����x��o�+�0�ӈ�����fX1��;A��Hh�r���Y�3�D� U�$�X|��I$+sMg�w��j'��ʳ�K�����&2>�jO��l�;$�|T�☃���S�~J�Mx����v���Qq+�R��GF��-��>�`Y�&��я�k��˚ם��Q����q�{��Xw�R�
ȋ��j���Z��[�F't�1X[%A�����?��bee��\��N��i�����e�b���Nk �b�����{N�r��}
cpq/7�1������}W� jQ��ج0iU'��Zg�!U��ϐ#��<�����e���������=�vU���<R\�ºȔ:�sJ��:��-���݀�^��j�a8R7������ş�nɝ7F����v���B���ݾyq���d���U�`�j��*&P)90�P�����/������Xd�Bn,��x�����u]1 üm�����Y�|no��!����yZѐC`M�͖�lm��_~���Vf��G���<�zou�<Ȏ~�R_i�%�T%�����N=���:?TRGix�y0U���Kc�0H~�f��&r�2�����'Il�9��<�|��e:�Xk6@��s���\6�K�"�y��#Y�?�˖��zA�,A�'����~F�����]���(��ԯ���z��R�
ԭW��w�����Iy>R��P����rx�0�LdIC�z��M1hJ�3��+@-c��9��QMNK֖H��6g&���}�$���S���J�+Z
�Y(׆�+>Y���|98\f-��]����ao�@G���L��� \g�0`��[��m+�ag^��W)��ߕ�b&��&�N�c)<�������,����?��+�L
�ʧ��n�˂��D���v��I���>�A��E�v@nx����+,�c?��
,�O6{f6��9�_|�l���O�
#��.�V��f�ưf�n��[�;�����@��Tr
��6��L���+D׌f��ÀE����n��]x')}J�H �p"�CmP�ܑf�j4��..ݧ'o1��(z��Z��xe��=e_�@-غ,q���z7��J�l����ȴ�n�yﾞ��B��ؑX��܋�/�."�YxLM�����x��v��=��%ے]�s��ՠG6����)3��:&�Y����N���{�ٱ4�ù��o$$�聵n�Gזs4�gf��=;�C�C{l_���f-{*6q�236�y�w��@������3	���H��Y�W���OxXL5�̗��m��5|*��t/D�hsHm���|����#��aL�����6e�M�usR�ĵ�b��>�[[N"��A'!�����<�?IO��$1��&��g�����=�Z4����R�Tv!|��L+�� ��8�`zݱi���Yg=T*_�Q�����:�~w�'-�I��u]�7fc��Ǭ��$�c
)��F�|f<Y!�:��g,�y�N=��� �&�Ը�g��:���J� ���>��[1�D1;{��	_��xP�j�����UB�gt�k2���mU\$����.a�"o��&ā[O�$��6�����?G��c��{{�gc���"���9�=6'm 䁡�q�-�2��^b!�V��P��O���(�-�[Z�G|���]�ֱՓ�_G{�{q�,�V+ýX�6�ˤX_��(�>)5�sA����ʾ�w�I�<?�1V���Ru�ڊ���W���8Կo��Z��՗9(w�a�#�{�m %�O'J�ީ�����*��+M�q�@��꼎,���?6�Z�W��T0
�;���?���'yA{e���J0�^5���^ȫ�_�7�ש��&�7�\Q~�+�Z^�v,�ۭ�����-ko�Gܠ>0�_����ۈ�D
����g��>���;[CS��aE���Oz\�j	 �{����B����K�Aɒ�7̦�Qg������IΧ��띇��j'E�B��.����3������f8[�	� me��n�L�+R����Ϛ<�!���vR38�Ơj�F�-��ٲ�99�Ξ�<�@ת:>���e&�����Ͳ�L�����s"q`\CX�'�Vj����Q�A�r�򹯈�������H%�5b�Є�U���E���\`9����D��	�;�X�F�嗹8�%2.?���k�>>W����;\"�[c����å�2�i¿��f-Vٷ�'[?��_�a�.��0r��`�yS+Ȟz��[���67�	�h��M-p��ɨ'�e�!%�L��)	=4.%��,B_3�H�Z)e��Մ>Q��Ϝ����K�&g�������+��e��ä�"\���P'�Β�:ȅK��n!��Mj�B���C����b��0��1�����ߋ8�����(�R�]�G���r	KI�3o��O��M��Ř�쮁mI�k�Z��ͅ�-�:�i<�y`K\�/q&�e-j"%DW���S����a�#9�~^�����k�W"̕�"�A�.D�ի�ޏ�F�0�?WQ�phb�̔��f}�c]Ra��MA�*��-��EڐJ�/�|�Dj�(��������u��iT�"��imdҥJXއ%}� עf^S؝7�kg����l�""c���R@XNp8�j�{��[$�Gh�'�k���G߈V��������X�ۋ�&��^!"��@u�v!�t�'�������F�DԼ��p>s�D[������_.����f(f0�
�����a��n��^'��um_�e߉�ۍ����%��/;mZ+˥=����(U���G5�� !�ڙ�R�|�{�i�����A+�ry��\l�������q�7������\�T��J\w�@����w�,,�'�z!��
p����w2�m���y7"/��=�/�=���?��.�Ez�WN}����~B�8��OI?|9H��x�s{Ho�:=( ��C��N��
w�o�;�вF7.���@��5�#Or��2 ���ݰ�t��4�>Kٕ.sX58�Ʊ�8�wFfБ��͋s����X��;�7C����t�Tg��n])͝�PNa���j���O�.�r$=�@����F��#��W���m��w~-��8���9Yɐ�F��(/9��o�CU Sc5�Α��F!� �X�JyѠt��K�����>`_����#�ي����up��s��V,3�>�/�ɜJ%�R�<v�*�M��}��[������������&o׿�.{[�Őf��~`���_B>S�i��]�m@��A �������d2�vA�,iS{� �1y������l��?��V:��S��UDs��]��6?�F'�á7[8
�w�A�[4��XE�}��ʺ�[����=3*��a�ҵm��z�	y3"sV����u��/N����!7H�3�eu���y��~�Ct��Ns{ zcP�cn=�����o��t��b�e�:��y�-�2�,Rqs������M�1���� ����(�q��3q~����i�8��u���|�q6H��B��lp�� ��$��@�S)Wd"7�T����7��U� 6"k3�o�6����V�a�?32\Vy;�FY�YNBއ�O��э�Y�5�QQh��c�B����?Pf����L�P�G������$?��&��$VM���N[�2��>�邈ҡ����u"9���=s}�]�DgD��_�)s�Dq	���	�fX(?x��,sOR��so$$^��Y?��T�E��4]U̓��� ���e.l�cc�+5��]s����B�P���"lS;v� Ɂ�`7F��5��֫w��[@r�ȸJR��� ���e����]�)����H�6��X$���ƝQp�7��e�5��u�+z̓��e�K�n�` ]�
.m|�ρ+o��Ҽ�2}��}֌̓Єe
���3˜�l���,#q��
� �B�uKC����_X�1��f���S�y��9��Pd1?}�H���5޼^'�Q�����z@ā7ߍ� ���]�oXgi9%�г��G���.�6��2��->N�:�q5�V\��^r�<�M
�z��6�l����^kՈ�}M3� ����G�z�C�t��;Z��N#��P����1w�I�z%vz=yu^�Ax�E\	�|����c�;-�zl&J�\���c�n��n�g�}�P�(��q�X�;w�S2���·��E� j�z��W*����ΗoJ�;ߟ����n��W��|S޾F����d����!����}�d+9p֢iӍ���<4��L��@�ߑ*iԤO�!>8�#�ELʡ����J7Y��$�b9�!z�)8�p��J`�U��B�s�W�V�`q
��}I��	��Y��s��RQ*��F�SkS|V{��#�ǨB�M&��@�	���FV.>\劋0�l2@b<ɯ���mjT��d/bf�����[1�4_N�d�'|����Т��gW������>#y�֒�n
�xv�{|*R�g��*��A�P����ۧ�{a�/���x��4���֐������T�z��/vM����f4��+���s�u��O���k0�nҷ���з�;�	������Dϳ_����Ƹ�����Nw�Bt��X7��\��{k{�{���
N[��`�6�/*��{Rd9�Cd3���+�ǽ�̗۝�1�+ۣ�������]N�[1��#�8�3k˯� E)9�ԇw���dw�nG_E|ʏ6F5�����N@켈�xz�c-��n�),6���s8v�e�b'�KS�Հ�ݑ���������5R��7��O����H�׿��_��O��Kq�֭Y��y��l�}٥5/�5���t�&!l� V�xacT�����e��3��{)4W���|bӤ�P���s��]L��9�2]iy���:�(�6�_F�n��޺n=-~m��H��ͼ�,���9���ZYt����������;k2�[I>�.�1��?����`�7~�	Wz���'��|~���j�g̯y�X��O�ء	�o��Y��u�m�^w��l�<�j���� ���4a�@��8[����>� �x�-� � ����&��N&T�%���Iu\A)��$�����a���Fٟ��C� o��ҙޡ�2��X��_%��������'�k|f/ȶrZM�O��Zǃ��b����f�tH��#B�Q�3z��~��m�J���j^��ӫ�����k~�@B���#Ҁ<������r�2hE��u�ͨ�~��ܯK���_�IT���̷� �������)������:"#����HuC{�|��^��3o�u!7	IӜ��V��N�����е	���gn�9o��!A���3�ݺK���	�m�~B�7���8����x��[JL|O�H�;l ��\�ܚj8D������w��$�Z����ʲ !��F3��Ys	�y��m�ݲ܎1�@
�VA�o�w�~M��?"]��_���N�����X���?d�'�0��G	���g��g��6��.������kV7N ܭ�e�8��xLbߝ!14�Uzļ�Pw���r� �{��-�Ə�6��Hy��a��:l���1��p�UO\�E���^/D���U��R���R�E�d���a_3������i�R�ߌ�I����%\�pJ쨉���Q�PN<ވp�%h��e�z��E�Ρ���HM���cF5yo�L$������+2�Le���;�]NCkg�c^�n�ͧ�̟ۚ��AM�3o��_�����������
[��Ő���2�M���8�z�n�Hzn[�4%^`mG<xV�u��ŝ�+ҙ	Ísd��7�z�\ݼ�甚d @��G�� ���'t���O��с�V]���Bϵ}Ma���gڴbҳ��D��,ݹmfA��	�����gN��0*f=�w�y��!������ENHS��~�j�4��}(���35A/UZ�B��t}��񠬺DdvNgr��Y�N��q��4+hNYE�5�� �«4`���!q(�{gH��&�񹯐��'��,���o��wjmo�s�|����9�U�$1ڤk��Z���ї�>m��+��Pq6�\����
2/�"�>��^lO]�}՗�զ��,V|����{�A.Bvᴅ��S���B�:�>���74�Hżl����Z������HH��@l�L�Cb�8�9Jb�&�Z�q/(xz���R%�b�U^��W�����풚����b� f�!���v�KӤ�,���ab库�M����)�� @���v��&5es�rn]N9S�dl�f��c��J$�	�|=	t\�/Yq~���ې���3`����x�_��+ܶ�İ�pӋx$��wV��'�4��=ρ�귇,�˓�g�M�I>	5u��@yc�p��2l��=�_1�M��!��	��,��bhA
�C��v�C�E�\|����e�L ��þ�D?��@KNZl��X
��'~\kH[d���NM3�Tꗴ��%� Ҽ���|z�*Iu{bl�# )g�++�ԃ�3���jWbHt���m�Y�'A:� ���Y2���F?�8�e�<)��v*b��B���f��=m���"mp+��k�EGkU�T��&���t��b�{a��󭼰��伡�T}D��*o����U�TA|��g�&,s<�)���!�\�ˇ?A����4�~�8i�IE���>�K��t����m�e���nk�Z�DWP�@&1K�Dc���� ��v�5��O��̖a+}��GNx!�W�>�8(�<;����dw�5|._��:���I�9A�	�G7)�,��	J-p�1��������Hzq�����X��(^-�O�vm�� ��d�l�N@o������ ��`*���H����pov������o������du�J��Ôq���A��g�Y��WOObfSOdf�a(gz(��јr*���A�m�%����=��sy��6k�X' N�Xu�a����+Lʜ��ڧsA�]!l����y���bS'��ɋ�¦K��e�F���Q��GC��T��Z�O_�a��뜚N�yi�e�s��kxh�x�Q/ׄ _,K��v\��Y�䮝�;7�d�F�S
�ۇ�(�~��V-��O���cd�Wt���;�+g�(���L-��f���2���9�� 	$������W&�Z��w��*�d?��JyS�����h��ZH���9*xrX5:�++bQ��:�e�8	[
Q�.�v]��I��0�[Vǐ/`,����!GI�$f���ҧыX�XRaa�ffV>�C��T\�l���+�!���q�0;�	i�bȃ����qM�*V�Q]� �]� @�_�:V`�T_���;(<��Pi|Q�o�k��ڀ�&$@�K�x
�0��S�F�F��S��*�����ƌG�3���ӹ�Y��jE��S1R����T?���]�l��>lUw�ҕ�EGFlۻY�C��Y�3u+^(�j�����D��h�&��r��
C6|��Ee6�^D5�~�s[����
�n,�*(>�����+�6��2
�'楔,���=�Y�K��ʈ_��.�JS���AM���J�0"��ʔ�R���ƠOR���'`�n�T������?%@k�6B]���~ЁX�#�x������xF<����]ӹgEs�/�2���&�������CV�� ����$BT,'��ީ��3�:odJ�R�!ޤ��#z݈2�n��ܷ�4$�ôa�� >;9MB�1~��ݢ�/�!Ə���
B��4��?�vP�;�K���A���zFN��s0[�ޓ/ �b.�:���T��m��=��xˏؘ6�������5�ϖ�.�Ej;=��/P�g���!�m4�^:gN���v:N�����ڞ�����帜F�<�E�`XFޗ�4��؆�9j����e��\n_�SaOcn��Q[7]�|�93ܤ~p#��+~9�du�,�v�_c(�-�8^�a�t
2�I���r6
������V8�6�~H(��Tꕌ=m$�S_�Ş(��Xpє}�!�� *�+�zc��d�1�Ǵ�l�J�ho�D%�=�бW�II4�0WQ�� �����օ������s�-�]���Lڤ��B��RW������{�M�4`q!Mi�V�ݳ�-�H�gģ�T<��}R᥈y����e�BI��Tb�|{Z�>�c���z�����E�'���{@��p@�Ƒ� o�9�d�X�WH=q4�'��m�V����@`Q)"�kG�^�F�<�_���᪥��µf�K�6)uXP��Cȍ�!3���;�3��w���?M-C�'<�����;11�	}]�wH�
C�<� Q���˻��r�E�v�p�d�u��L�<�������^�֕v}��\�'e��G�(d��%���,|�e���MG�o6��" �F�pEF"8;'ḉI<�L��O��q�ཊ<����]$*����/uy�ܧs4Z�!�3M]\�i����XH�z�q�o�g���F	�้ S{~���O-ӼW�����8H���0��_��EF���m�%��v6-���LҊ�E���/�)XE�m��N������Wo�Ю��w��,��h�_������Kv �(#��yrT`5�zh!* �a�:�yݙ�Y	s�H�/X��#ݣkG��4���ʦ4a߯.��H�:�J��:Kr2��į�� �������٬k̹���se)�dl'����'?���~����0���f���n� �_��x�bO�L�?H
�t���C�_Ƶ��4ù�a�1����shFf���_Q��&y(�+Dl�Mu�zm����윋�t��E�S{�eѴ�˙l��{�M�T��.4��� �Z��N�I�S%��0i���e����r�n��3Bf脞�
3Ou��	���dk2�*��#/�b0�hn�ZR�����o�¤��@-�=��C����z��i0�v`܀Q�y���r'�Cz��/<��= C0�|U��|<���5k�꫏B��?�8 �[R2�m�*|#�}N)]�?�8T�n3̦·�aqoB��l�i3��] ��vĳdz��;����+~DiFj��j>��(�sK��")� R��M%��1'�Uj�+���U���5K��#6y~T/�cv^t�����]h�V,W$�P1�D��5O8��� )OK"�`=��a�����R���H�j��Y@h ط��"d�V�B։��K�z1�܅�ޮ����Pj���T�1�@I7R���j����NM-<��������r��5-}�w�><Z~`�J�Μ���	^Q)I6*��C�Az����#�N2�H�����>�Ĉ 虾}�)�g몧���
���q Ks�3yJq�����V�R������2 ��Z������ۙ~	6��D��R���f����<)��  �7�#G[�z�%���Y�/	���~폙jDD�=٤	�s6��<,��yG�t'���7���*����{�W�SpA�
���P��!Cn�xvK�xˡ*g�$$�Ά�����0���E$����p(0��ǢT���cx�V���)VS9��U(��!�[Nu��]p��C��	�9�Zu�K"N��G9���s�d�D�9��M�z7^�bb�� �hB��zwPk�f�}�ܸN9�Fe��{6�0��)B�_4$��7��paN�ւ��]������s#��J��{�0�nn�Z(W���M�e�)��+�g���W�j�#4ve�	���߆��Y¼��\���@b�y�+;��Q���{��z�iY�b,��E3�z.`Z��9������,��W6{�d:LnN�B՘Gt!�GL)��6�ܺM;�p�6�.���)�m ;�;S4AE��U�
wՇu��ˉTei���|��c��拋j�$�L�q�>�\$p��b�V����$욈���T�k/�_��^F}!��꺸��SVC,[(�#X�m}B�G/LAT��h\u�r��d��x��z��m���p�3�:O!�1ƛ��_	���a}����-	wϏN�pIf(�C�?Rh�}�wW��������~9��� �U�X�@j����d��#T��ی��E.��%�As��:��m/��v�2k�{P��t��=��2������-����'�R����G�j��bl0W�9�T�Ow�@���v�19���{�0�J���;Hq��Rӥ~��dm�/�; �]��5��X��������$p����~>w�K� l���򤕐��2m�Qxny/~!2� �6Hq�#�9t��}�~s5P\4���q_K�|�{��A���VP,@��&���3[�2��3b V�g�▔��وPlԬ��~[Y�~�����^�e���雸HYX�n���/fm��cB{��'�u�q`ǷP�����\�u%U"O�Α���#7�6�)�q�~�{B|� ���H�v9�-�J*q�u�� �$�/k�?��r�x�#����u'��=	��h՗�y�F;!�V����`u��'��ڸG�+��*#?����/iC}�g�T	���v��zwR����Df�����J�un[�Y�"�b2��
�/OSq��wN�@"��qY�{%�<�u�P�@��7�!���r�GLpz:���f�R<Sx���Ɇ�����MmJ����Iװ7ٯ�Oo}�O��I>�[����f��H&٤KX.���	<[�K$Ҝ����[H��.
�x���������&�tt��m�S3H��*��g��@���TT����wV¬O�t�'���yX���jtQ��PS[�(X�Px�kY_&pX�r=��&So�#w{�:R��~��R�-D�K�ɁK�$�'��-@�g^T��vh��s����bNp����@��
Ж��'�]���ݖ��s /I�Ƃu���㍖xQ�}�b���d�l����L2�T3�z,��cP��|�j�������ޔ�&q>��!7�R����k��%�
�cд�b�ź�}�x�{����`�Ҿ#��' ��t=���9K�O�1,�������*�kVB;!F�'E��Wt��~�����I�6F��BRQ�B�x�1v�$�q�C�I͹�UM����w^�>�S�k���PC)�R4~@O��C�k� ���!��J7L4��L�j��^��-JO�)ό6�_�9�S�t�R ��3g6D&y:w�Q1�0|�~Q# ��T>�RQ����2%�����6,i�N����x�¹ \��T���������\���+��N���Fy-��FX��M�{u2�Vӓ���<	R�j г�/1�?�����<�~ȹ�HmfRlEi�f����?h6'�A�o����M�MYt�o��]%�j/���ƚ��L냒�0���k�x���D㶰���C���8�&�!���?w���:�1�Ґ(Q
MT�d�� V�<��t\��K���x���tWa[<��Ed�!���>����K���I���;u�ޥ7}9XU���%}���8N@������v(5����B%���l��n�VF���81�=�lQ �m6���s�@��o������?��L���vS�SN:7�9C�X�@�Lt	��B� � (�u�+����.ɰT��|ײ$�%PX	����)8CGttx٥�Y���V�TI�9��G�p������<�@7>�Q�%6��	�Yl��@��daħJ��^-8�0U�d_d?�Tw�)����,G=�O���A�h����_]� �����Xh��8�����n$n��>+7hqW5���%4���\
�g�QP�8� ���Е�ȖHt�!��]���}���S44��i���rR���A+�Hf3�j�2����zd=Z�"Ϻɴ�����Z��ڞ$R�v0��9;Ҙ�X<1��7����L�?mz��AC듦t2-o���HDfa�3�����;Cg���_�&-4�X3�I�}5�Hxx��I��+W���uޛc�¨;����J��E���&� �* DG���ɇ��ף���0����:�6
Ӵ����1*�� �uV��j��%�g��&����ޗ��_�p�+�a�^�$`o'd�	c�Ǥ:��J!�W,�1�)��d�����Q� �C\
�a�H��DW9K[��ӧ�"��u�v
�5�ˍ8_s$��3���/�	�������;����QT�5F�:ȯ�5���=;}hd�?�E����Jn�
�P�K�<)�������q�� =$��}ɱ��l���9%���`��E�L��\bHL$�L���ڟSu�Y�����dAn{�w�� ��!
���^lmuB��5�T���#����Բ.�����e���:���/�(%�rv�E��i)y��
P�/��p��4=�񇦪N����j��Y���ʭ75�����Fz�Z���pv��&{xxm��%�	k|�qi��2F���lw�S�c�#+�����h�H���$wiZ*�"���+pF��Eu�n�v̒���q=��~�sZY�{�V_��Oe�������Oe&b�?\�ƉK����0����Dv=��\t0e���r�+�t!�g��7`�Z��Oj$O3�A2�Rw�U�q�0��{:\T3z����Y� ��i����UY�]��1ҬVΑ�
�Qحv�]����B��׀�%$luW���岲ڦ ����H�t]{.�n��J`̛0�_z��������:�7�V������k'��WdZ
M��d�*��(�Z�U��`�Y�z���`%�"�����=S�P�pt�GvpL7�eC_*�B�'+5�p�pE�/a�+G�#	��<���-E,i��;���ڒ�)�2=Joɤ-����?P�kU~`cwM�r����>��b���%��nZd>�Jyn>��Zn)B\��&���5����:�$ǖ�ir^�"�^c���H�]��n�����[�"�=�qT�׈���t�*����s�pF@pX-�7�F$~i4)O����Ti�����H���n��w1n�[�`��T���m��gb��>w�Q�`F� �ͧO�����K�"��'NVJx;t�[�P��=�V��<_��iý��@h�-�s�! �����a~JJI�I�\y���T�@lF�
'�.)q���%4�݌�@ ��qF�n�Hg��B��b�6�)�"x�fX�\�/�`G�$Kz��x5�����28���@�UI�(�?�)�h�l��-���/��"N��Q�8G���ey@
�֧"��(WrO�?^@&o�Y.��P�+��hG�0'jR_��o '�3iѩ��H�&h�N�Gɏ�
#N��F-3��m�d�rRl>Ivv���#��������C�%���tZ֧�J2��ez�-�
�bC�%��t@��10��7H�]8�bi��$$_�a\j)��-O?j�k��5�����S0��,����M;ET�+e��G:��n��7 ��n��,ܴ��.� {8-E�����d$h��9�jm��,4:聠k-�  �̍�d�%VL�u��j�e���y�T���{N%�v@���K�P��|�pS #���	잆ߕ��3<\uHC8?�&l={�������
�}�".������\��Go��Չ	�$��5pȜ)��;�j��A�\D���A.�M���SO:5n&t�>�.�0;����$a㛰�D��W�)�b"����X\HQ�ͤU�k��h^g�����_,�Q8g���]R*hw
4t�:d�c>:�+I�L�,KK�PԲ��?/�NW%�3?��_�[N~� (�Ƽ�[3�^T��h+�®�![���,�:Coh,*�>a��a5�7,���)������6~r ^ދ�(�"��|��__j�F��6��ϹV8�
t�>8�]Bǳ=� ��/�&�C��:��i��n�dWől2E8�$��}�������_nyŶ���1�g)
t�C�ٶ�"�#:6i�5q�	��βi�c.����(�V�5�����YUg5?���9/�x'��-s�H.J�]�D"����ާ�l;K�twp�q���^���$�?'+$�3t�Y�$(��؞y}x#+���BH6��w����\,��[��F9��La83n�Gg��������v,>���b���'�Iڀ�	���dY]��|��@�Rt�>��;#��	ev�a���dJB��ܛq=A�>?V8Ρ �s�&�ݪ�v�!x�44u�`�3��t���1{ި�|��*'�0������`�|�.�<���&K*�����@u����G�&��҂�V�+k̀��R�;�Q�|e���ǣ�g�7�Q�@-ЏS��z�Z7+>�e2¢x�`L^��YaC���)
��r�h���3���b�B���=I�IE󬽇p<�}�?9�=��zA� p?P�0�*��tr�{ٰ�F���㜩,E�7d�B��U��k]j���Q�&�?h���G�����[�^E\]a� _C���=9��M!�i�4��N��Cf-H��q$�5ic���o�-�1�~D���݂�c�����я�:p5.��C��ݑ�z�Q�}�<��R����ܲ��"|(���.� �>���M�Z���d�53���i�j��A~:�����{�n)f�j��0t��#���*_�d����CBd�8�lk��޷(�Ɇ���RhW��^��EZJ�O�/J·�ne�j�H6P�2��T��?�6Z��5F�G�f�$ >$��/���P�A��*�>�6��T��J
�@	tP �zS����g�A�W1�NQ ~<F!��������p��T����T-�Pg3 PwƜ��NX�Ĳ7�9R�h~����q�vJ��|��H�o��:���뒂${�S��j��>v�CG�xk���It]t���U�q�˹��(�T"m<DT%��i���:��xˣ���͆��x�Il;͌2�~2yc#v������ ��N}Ve\Bޘ����}GJׅ0���'Qv��D%iX��|�͍8�zW�5�2Hч}���p������,�����P��^��MQ�)��+ R�^�a�%w`�B�jǜu)�ح%&�b��_�	��z����
�ˎ��p��J#0�;�B��\��]V���W�Bf����;xq�lj��Br(H��;�4���&��OD��򵓀"`:ޯܐϰL#��b����s��D�_���-�;��]�׋�
�4T'b��K��/GӞ`c��[��II�q�2��4Kc����}1�c�^_�V�(lh�ѨCU|׳�Bl^�ݦǴZ[ȃ��z��M����B�Ę��8S�I���k�}d;���tS6eϬ�CA��;`������f1Y*�l���վ�_�6oy��|��W��؏�
b�1v9K_x�%!��}�MM���z��t�9졶�G���l7{�r�Uˣ�9/#�,�z�,C��#���룄��"e�"s�U�F����F�}{�'�n��եg���<G3>&+�Y[�L�@ÓKB��Z� D���T4=��=�4\!g��	��{��ڽ�^�'�gqJ	$�1�g$>�����_mf�{X����C��Y+�Vy�b$��#F8F�����2'��סڈ*�o}�[y�vҸCU!���2�z�E �=�M"�:�]��f����,\Uv�������霊Һ·� �w0�2�r����@���";���W}�����R�é�u��<E~k�);�/A,M�L�I��6F��5/��H�t�ؤӕ�;��|��/7_l�X�7-��=�CZF�:�:�����Y��3�沮+'%��W�ew�La�M�'�����Ǭ�����FZ�}p�s"|�ކ1�]�1��Xm{��JS�}J_���z���*�Q�@�j�����p�T��bQ1������b� �nqH��Y�`dA�,a��W����@</�)���-��$#�p@d���́�)尤V�{��+��@�� �uc:���0�Z#��1N{��e������X���+�)|]`�7��!���,���m�)��нgY�H!���6 l���%voi��
�	�U��%��U�<��zm�	^���;N������cu�q~�ol>�����/'9�%�̦�<9��Z9�m� �3|hH�[^E���ǀ����*�F��U��qo)lñ�*�f��ɲǑ]s�%2�N�u�s�� ���I�(�:2�,�T�j
�y��0�%{��,��.ٷ��=�΃Hc�A 8I)��fYa�0����:����Qx�dM��@��lI���8� ��<��>l\��X����tt���uer0��%�����gHOu����b�m]���>J��
���������D²B��T��dJ7�vF�)+�'�3��I��P��K�O�d؂K�4�bz����o�Z�����#Oa^R5�O����[ne�{K�2��Ϝ����vVI�7�������	>�T�Ā�|A���� �9��P�u�~�;���%($O/ie�$�b0͏?9 ט�e�?h9��ٖ�5U��l%<[YFaL�������"&H�6be������X ZdT�+v�6z��*A\���	ŧZ#�sK�"�Dm$S!�U�����EV�%�����8>�
o?��cD�]G�}/.c0����xě2QZ1~{�\[��)�,����!*��)7�g�∎ɲ�����7%��nG�!�.�ݡE����v,� �WodĊ�h��{������un��4�qLC℠�R�a���hԥ}�p��d�f4	U�����\�	ʿ�|�@U�j}1v��"C�e��N�!�O�(Wc?�'Ү�I�F3��}��z��[��.�↬����K�؅�'[��N��P.�ѣ����k�ޙ/_W�=�q�(=�P�rR�� ��t���6%�pA�dؒ�ɸ�Cg��ʳ�s�EZ})r��<���-���@:^��FVcY�I��w������;WBa���R _��u�:~��k�K�5x��?�4;C��Mj�Ns�iA.�����K`����	s%���W�¸+lV/�KZ-G�c�0��z��u����ڊ1����E�0���>gd�sTW`��سk\''�
�L�9��/�~'P,�dm�9ԅ���O����ݞ��0�'Z����!-!�/��z���t�9���ç+�͙{��e6�2�<���I17�M+f� @</yd��WV%ǌ?����<�ET�#| ,Ⱥq.S��[�E-�0���a�|��pY�ģf�̙R�A!b��U��D{Z��fZ߲�
F�v^��p�������1�(v.���ͷ�B�4�Lpw4$X��)ߜ�na���<!�)"����ܦ*�b=����=�@مB��5��I�괦�?B��S����s�º���#Ӻ�9UZ�?{#ZC�iU�?6~�#0]^��y��Z��|*<A8�c���e���N���"#y��q�������py�W �,ϲ�X�����	�\ss��d�j,�&hxW��Sa��ewVq\C�em-�1��u���{���H�-8���#�A�<�>3*�x���ꪚjӦ�}WM �^��>��Lc�,�����?��c�;��b%�uSU�qly ��(N��� �3����� Ox��K�2�[$6�X���T��SZT�Al\��z��DOU���f����ĉ�e͠d�T+�d�������(y���Bg��AZ��\X�qΓMf��y&��hy��D����5~��b�ŕ�9���o��!-F	/2 ?��,���R_�m4 ��Z�y�̈P������T`���ߏ�`?�b;vB��֢)�k5pj|Uaǐ���Zj����Mj8� 1
�R�mUd������n?w��S��ơ/��eYO�b����L)�=JRϦ�@�p�S��
�9XQ�˫f,���e��-�YZ�y��,���L�o���w@[]�{x1��[j+�d.zy=r�R����T�9q�3k�k xXZ߇��)�^�;�cmE4�%��YLaҵ�7\O`3�+"��~|�]V���x�9Uf$H�m$Oj�\�FDE���ʰ�� +�O�7����#�vA��?Y��Z�vpvW�g�5��f4Г�*kn��8q��G�]���M�T>���L��'#-2�&�d�J4~�	߹(�&���:C��~ۖ-��:�rY���}?��ѐ����?�ƿ n�s.����Ӆ%0�2�sTq�^��5�g#��*�����UT�7x
3n����A��l�SnY�v��&_f��G*3=�y���ߗ�Iz%�W��*ك�X(���E�ל�5mL���0��(��|�e��ʜMܱ�'��1.�l�J|Ԛ!9�	��x�!�	�C�`����|�۫�U$2�F�/�)���d՜u��O�H�*��?�U_m�+�
<YO�_������K��	FU'���*�}��+~�S�b3�D���^�ݟD��� ���>��=d��~V�.�6��	�(��r4E�\McZ���_>�v&;^bNa��a���rn�ϖ��tr���VsF�o�M���[�qz���ը[�����Jષ<��Lʜk���xɹ�(�.	�=��)�����UK�i��a�S>@�)r��b7v
s�r=������;���H�p-��pj ��%BݨO����.2z��	yq�dsE�v&��hUF��N�$b��y����}�W��(�b0F����X���+�l�3Pv�F	)V������?IIM~�9��F{\��N�w�hm�I�Y�k1Nҽ�Hى�z?�c ��2�c,&�uu%�j��Xk}��~�mѣ%�MEA�H/\QcM����
WG�Ȟ��~r��#Qo�4,s���Y�㗦�Y '�65=�0a�o1��qQq���'�h���e�-?���7��������{9�[��/��5u�A k�(H`{�><�Eb�M������4�������un��̥у=��^�ۦ�L�}�{�Z$ӈC��k"�i�㝃q������yu7{������p0��i�����e!�~��T�B�S�9��Py��:!��L��d�.,�Eq]nH��E'��P����/���5�t�2Q�>��vR	a�N�P���l�G�O*@�n�3��;U'4���令�ǘ��tM�KČ�¼���Y� �A_�/u>"&L����\-���p�\?x��j:�Fd��R��=b�x;(,ÉԪ����C!O5֖�6o�O-Ӌ:��BKܑ������@��JJ0��^�����X�)�$�@+��J"C�f4?��'���ω���qށ�`���A��?���Hs��śt��ϸ;�x��W���g9]r��y���<��Oj�J'(㭉|PS(rj�3�>�����S�hoc0]P��x<)bh���Ы�\�x$�Z��{���8��?R��v��HWET�Ƨ"���l���y��|��~�;:�he|��1���7cy�@3X��@�͋���l.���4�H��L&y1�k��:��!��7�il��"�"T�>�!�K��<���tʶ���&��n�$��-O[�`���%����+����Wؙ� ��+��Jb	�2�`/�-�o��S�Һ����{�,�5�^D���n��hnl�fH�)ɟ�$^h#S_Ո՟��"��ՙ^x�����a�@�������9��%Z��Ȭ��q��dMT��d�OG�� ��*T�t���+L��S�d���_̨��_���B]'�XNG�(`��*����
y�������8�!Z��c�f��\�Nx��W�蟓��^V:\Sќ�{j%D��v:�p&c3�)�g�g6���Q��2�bJh��n�t3�Q�%h��&n�����<˕����s�_;�i�� ��Oh�6S3 Ff�����^��hNT��`Ul�Srn���h�C�^�td|�UQh�g[��*\�����G�p�-�t��d�M����V6<-�/��B �p9��E[)ef�K�$��>�����[.�d�q���4�p�q��e��	0�A4>�5[���}��1�q/�nso�=��j{Q&�Msԍ�}�*�5�s)D��m�q�KƉ�j�,��\p�T>8�\z%M� ��2�4�/"/����{��XӦ1��HCg��M��l�3���1 ���A��t���Цo��Y}��a��_U՞'N6��=n]r��� ��:f��E�\�!f�h�բ�(�N	{�0O��H�����Ȁ����� �Q���q�M\m*��*��l_��J21�'�Sa�@�.�p���yE9��=� ����j�@֪#�� ����`A�M<�b����­����D(�6�R����OĠ�ɗl\}�P_a1*Ki�$o�.H	�]T�'��Y�`�U�K2�Kf���PU�N�`&�Ϝ@eM>C��{�����E�zVzs��?s��L�I,�3Ɣ��j�a,�A}]��;-�&l��Pu!o�Xy�䇜a��nЅU��3�?�����|��F�X�O�u�E�Wޤ��ú&�N�1�[�S.G$�2J;�أ��o�4�1"" ��YR�_��νl���ّTέ�yVs�t��<��,�4d�W!�s#}�!�&�v�
�ސ0��C[�E�s�Ku��d8MCi����%�)� G����Or��]�xi�*퓐�^�x��-�i@�ړ����e��"wV}qv{�/������i�A���w���@u_�v��4�}Yz���_'�L?w�����,���Ǒ��g�$h��M}�2Z�.E)~�B:jS_�X�.�e2�
����W�$<]�����a&[7��ǡmkyA�� �̋7^���r-�� �Q��,5�Z�;��	�{2���/}�$��d�ʆ��2b�qb��,��	�,�|K�d&wG{�9�+߀~�FP^�ƅ@���
�Ь��mx�Pڹx0�'���^��bN���}2۾­h>==�{�B~���G}	���[��� b����'�%C�d��tKN���2�("�F���j$��ڙ�*Ϧ��������p�1z����#z�:�@�x��,�}�T�t�BF�T���:�'�{G#��:a��5n�;��y�hX1(��:$u�R�m�5�p��0g�Vqw=ܠf�HrX���19�H ���،R%�ʦ3��=���S�3�'�,����E��YҾ�턺Ma_��Ty��s�BxHi-��$�ض����aG��峺���QW�"�P��+��t}���/�R�T��u�Sb���re@�/���?�l�~�)��|��)^;6;-˛�(Iy��2Z�z����J^�z<Hz�忳���]I�g�:ǯx�cX%U��{�N_k�}w� ���	m�����6���֑��o�b���үg'�!�{��9�> )Pp�6�;�J�y3R���4�Q����S�����8��JN��l�[�(�j&���}IN.v
��!��w����^<3޺��2^�˦D(�TKq�S#/l;��l-�e��$X4�qTh��r`�1�Ƥ�V��	q1A�S��Z��:�$o��4O���j�<����X*)��0�?2o����3��߽V��ѻ���:�s�9i@[E��Çy^p��v[���g�/����S� ���m1���o)8��i��I��0���ʢg��͚�>g�s���7Q��%L�k��c�����d\�>�`����ݚޛ���R��ʚ?��RB"e1n�v���n�GG���ci��R���c�޺ٓ�:�>��P(aZ,WZ��&���æ:i���R,��X>��,Sq�R.{-z-C�Q��/j�f�m,��t'�_M,@$�d��ǌ��x(�Њ�����fw}��+Q�����	�����`F�7��_G�e���s�$���-�wP�'�nC��ݎ�X)�y����p܇c\JB��3h�{:����co����V	i�/|�$I�� �_��|�mN)N`�N- Ih��Iv�dX��sI,�������BD���ݣ�2��$�z���	S�p��a��m>G� �Fm�5�}u�z��@�����h5���xA�k�9}z�#�:�;KF��,��2+�|5m7����Ж�n�Q.�^w��;)����:�'}�z�L�s8�~��U^ɺ[Iu�O�Ǎ
�0�����5o�GC��!�69���ﮩW���
q#��/��g�CJmY,P�Q4���T�oA!�!ǫu���X�O)���L�`�$m$'��ϵ�u�3��<Z%���z��"�g�Ko�
Π� i�d�}�;a*h�Dk��D伫 �1o9�y��Ju��
P��E��I*r�����7?^�=����/����xqۛR��	���Rٖ�l�4�M�f�,���h��WE�b2%�A;����]Җ���K�[?�f3��( �N@��e���:_��~Jv�w�,�/�=mϱ�S�����V�1D�����R�>�B����?2�����8DF�;RG���,�B�� ���/�<O��>M���"ձ�izK���&���#ER~���D�`HK|6�.�v� Q�?c�hE�wi�6�Cg�&���W���s� j'�߳]!��:�����D~0��d��*<��>z��B���9�Z��f,���ի3�Ml�YǭHf��އJ����]Ŵed��FTV�l�<��%��r��,�߂w��,��E����h�Y�TXs� D�y���:ĳU7�t?�����H�yg���`z��͔0��C�D6ge��Xp5��x�|��F#�Z,����f���UNO���'�{<�hO��G���4�Z��?[6�ĵ����2V�ϙ+o��$m5n~�&A��W���>|u��"z$��6�@�5��Dr����-�t�[t0ń�L��9=E���e��V��nx������M+��L'#�g�L��ѢnS�!���zѫ�9z���(�2_��k 7��˚t��(uc庫P���F(���LcG�5,	Ψ?�@��(��J�Ur��A��ħO�����nD�8�RL�a}�T�V?�� ���5w�B6+K^E��/�vN��(f��!~oI��Q	�;��k7K9�bfJ���(!�C��S�+b��琎�d�$��+ ޚS4�_`�����qI]&�3[J�����VC��!=�<���6��49�W,�*���0��k~iQa�Cȫ�t��Klk�U�hg.���-⍼��M��������pUR�6����SD|0���L���a�
9y�+a��b���!��O��%�(�{L9/�}�I��v�s���B���E^�he�e0~	_o]�%���cЬ�U�Ҽ4��L���ݖ���+���2����Yz6�@��W}�S��"�3 �.�_���)���ӫ�y*��W��r�C$+=:փ0�BV�ԤƜ�:R���[��:.4mL���^6���(�$I Am��׾P�\Ӓ�v��`��V�� lW�߂��2�!˜;�V&=Ϥ�dZ�S)�u�66��>-ti�=��#����"x��C��$�:m�V�}M[����,h��Y���t^�>54]�����*������ @Ő9��%���v	���C��nTi�\_l�-�h�*��To�!�z���ơ?�R�E7���N�)? ��7�Q���ѓ��\NT�&��YyM����G�{zk
m����
�f��m*&���]�#V���S�\�{�\��h��UؚD����92X1�S`�-���ǼD�����j�+Hĉ%�or�\Ա��2̘�u�}�z`�B��#U:�)їS���BvR�ā�����q�w��:R���M~ߍ���Nv�r`G'mv�1]Ν�'^39�{0p˖6� R%��!1��ݑ{5�������ly�
� ��=��%�I���ә��?�7���`4:Cľ����j �{*]��?����w�I���\���G�Ês�h(�*J����Z�WՈ�a3Ot g�5򁨬��}Hɑ���fVzs_Q��r�"7�*�N�q�����K%؁:r�ư/�y8�-H�	��Q�Y�O<.�F!���&�z-�Q�.kxa�7�����d��~�Zp
������I�3ػXPvnNO[�Z�l��7�l��>ߡn���.�z`u�C�&w�е+�U�`3�g��#��G�K����)E�:�����W�e�jM�l����T��hu'_PT9UhVm�/�9����37׳nlz]Y��Z]���X�g,_��R��� �V��E�`WC�ܿ�3�����+Ĭ΢6������\$�4�_$?�,��J`�����^T�����T,X�2��-����ڻCdZ3���Եփi� !���fP�o����k��4�N�#	Ą����݃��*/g��I-�E�1�է�)ps�	�k ��л�!�Y�x��V���ʊ��/�k��y�������-JV�;�>��r_̆e*��+1�9נ�+�����пc�&�+�P�X��V��<���E�M	*��K��T#y�_Ս��#��E>D���4$�� �\'����B?����#� ;_��5�iQ��&I�U}&��Iv��Cf:�.מ���3���n�S^0MmpӇl���1t�r�_�����A�r2)�\n�8.R��acn�e-�ǭ{N����m/��Q�-�}#�z���:�&<�����cA�S ��: p�s�#��2�)n�������-&s'�q@���	-�&�Α��e'D`�*���VY�98a�0�<z����e�����[�>�k*��v]�DT�������I��q���bF�9�F_5�`x�&J�ui�_��\.s���}�g�?E/��ߟ���_R*�0�1d�J��c&�&d�x˼�L "���u���]*�,�?0(�YsQ&,_G��z���i�Ѱ�k���^�؅�V���2E'N௟A���kL��[,����#����y4ѫ�i:\j	
�ٮ�3|���ǠҤ����#�I!���E��Dߑe�������݄�BD���-�S����P�keѿ��|KX7���� �F�8����怗�7�82�b�i��x���9 6�.��c.,�Jj�r!H�x�k���+�ⅈ'0�����:-M���!�r����j�ͽ�����e��w�kR�򩠔�Yf�v�і��o�Y:X�b�&�K�Ͱ��"�̜t�<�U|=�/.v�Oy;�0S�7���� 6�9@�č�)X��O���F�R�X��+Ov����E�L}q��U�`���6�s�n'�${F�1�'��j�S-�f�V�пbw�y���-h���ƭ���Q4�-g�l�L4*�>�}�i���1�p��.C��'X��aX�-*&+�Os�pc��*�K��|1
�9���z;[*��Pc���|�`TsGz�An�s���@��D�[{�J:��u��ΑUƙ�^Ь�z�Ag���Qbǖϛk�g=6ܘ;b#^q�
�i��ô/ƥ��ߋo��j��.�rd	tc��$	�_z0*R��>�������I_���}��e�;���/=>s`5�[��h��������</V1����'A%�"i�/���;+�/����5�;8`�p�t����Y��ŐW��Y����K�H`�*�03���Q
�b]���sS
L8��B�� �l����?|ZU�u���8u�
�xO��2$]�m`�>�
�Μp���+�F�}�xf��b����NUO�n.�3�y H�IJ$�[y��e|��L7:�Ł������R�3b͜P%e��~퐚�ϸ�ة�Q��� ��K��Y�z4��4�����b�bb�Y�\(9�����k;�g��\.?6��a�4!����jE�]r�q�C��!�>�C�����	؊p�Ewx���Rݹ�oA�}u����m/X����D�EO&@:�t�.��d� ��Wu���l�����!_x��Q`]|��~:�m +�g�i=�!;�	7\R������2+��HzU�mr��迡O�H!��&�x�X�[��q*C ;�$Yai/�TX�m?�B"&[�Ӹ^Ǣ.x9�r.����կեCKY6�=:Լ�����p#��C=u��Y�)9�K�ϻ ����B�Y�)e e����-�_�=f����t�����"������H�jx�\�@yQ����u��;�������0�&�]3BV�ʉ|8d�-�ڢ���������" �G���}6#63�_,�5����x8��_s]x��mi`<O���� ��"f���m�=� @M��R���!m'\Td��~��ˉ�4���t!*m�y�>m@Z�����J���_�k;�x�]��)̄L�Lu%���ɯY ���M�,�J�˓��A ���Sy��'�,��eA@#f���K��&��ҙ�XwдG�3�q����r�� %id����_)�]6܆�qOfl�%�ʺ��yy�&O�0CBO����I�#39xF�P�^S=�"�������\ �ˍIh��ʇ�f�l,g�R�'8i޴����m��K�3?d&o��-����'�b�A�w��=���ɱ�[\v59z:����Ssn������f3:]��U�δ}�4��ƶ~�?�~�x�`���rJ��g��S�P%ɅA�^>H`������:�C���<~ֶuHk��gn��
`��m#�h�g��x�[��&���{���������������JJJ|�\����9�҆�\�����ҢZCV�R�a�r̳�/()<�҉4 1�)���q�3��q'V`���E����ؕ(.X����N���ӆlh�g���J�)��I�?N�̒yp���Αlv5���?�X�'��^�L�Y���	�r��G��)�-�m�����Z>�&Lۨ�9_<�����H?���~���B��.s
eݰ�.�,ۗ$�&�.,����p�bh�%����Qy��IM�9D�B�<���O(Y��н~�Y��1��x����i����r���3}#��sr�� ]�2*���RHK��#3��D�<٠��r0lߔ4x��9X�y3p��;57	f�G4`�7��>n���9��~��GQ��8�x� �y9ubek��xa�(�p;ʄ�]�����$�_�{/s�7^�ɱ�0�}��A����~aU�e	�Ӄ$��
 ��ik�� ]���
��j���#-��t�����i�r��Ry��.������{SѤ*lI�$���rJ��?AS� �@�x(�b�^ʝP[Z)^R�څ-��7[��L�qY�l$�Q߫{nz��)S�z�o�_����UJ�\�y)c����������h���]�"TWjv*JSz.Xj�Is�8a���Hdπ*��{�'U~��]ͦ�EH��u^���j/w��Wj��[?#�S��3џX1��l0'Żۙ��*g�j�@���.,Pq�a�Ψ7MB�}����<#m�VN�)��,�0��l�dX�4wꔖ���>cׅj�{��b��t%]��E�O7�u]ӆ�?��^�7]����:X��<WV'�~�f��R�9��_?���?>\��G�F&�=�Ԁ�˚�rʑ�_��L�5��Ԇ�]���@��Ț8�g%���@-�$v��[�M21@���f�p�*hLv+ţ�dfQ�r�9:w�_ڨךb�W�+��;��P�Y#e\�BF���km��eP��]B����5u��a;�hA7�Y���6m����¤���x;��(E&"�������s�<������kHАBF9&q�0�1���}ItJ]��f/�tZ)��nKl��d|$G�ۊٓt@���3�e�&�93��u�pG �������rRJ�K���Y�#D���� 3���C�CP�y�I�,(���kO��Q�-�>sS�����0�s���O,�]i��
�$�e��Rv��6�`aTu���ٍ�K�@�Gă!t汤ov�l=�d`��k�bfTq��L�|s��:����T��1�M�(U���'��[!� q ��yx��z�wU�2����$��#�xO|�3� ���G�|��m���F�X�SV(e7F�Áu��7��ez]�&&!#0s��<��e�F�a9�'�����7L�-���$���$�)�Q$i}E��D�<I���NB*�a.K���cQ�(��e�M��j���<]��K�& �o��^v/��iE�
�+Yd�0;���N������}CR�vB���ˋ�QT��۲w�`��G%>��[��md�����t��SE5x �����͋w���s����h���p�NV��fI��/TI�u!����
��)�����y�P�x"���]���e<�,f�u!z�@��B�m-�*�Zn�Nv� �e��	`�-?p`�_MP�"tD;�j{G	����,��ګi� ����0��??�I�^�Gr6eV2���ܸBy�V�_{��;���Y�S���qڅ��+(��K��sN�A���N	S��4ȍ�[ih�oL!��`���߱cnI�����S��[��ڜ�9(�:���)���N��2O�+�?��ߤ��c��1�п"ޫ
�_��li�4��3�E�*�:��a7؈���/�P���J{���P���IwQ�P��ysbf��(N����S�^�>WC ��d(@�UXv�J�;�R|�F
�&J��L{(S9�xS�T�����-2���F�+[[i�-Sis-��\�`z^"�2MZ������`"_)��D�h�~�C-;���uxD�t�B%^0��t��%�u(kh;a�P`U,hI�ќ��ގZk���1o�ͳ��O��d'�p�9=^m��0ˍׄ�A��P+#�������k���v(��*�^����R�y�~~��� (��-U2.�!�$�� ��.H�� C���� +�/k��+��b�$:����aӑ.;Ő��%�+^�5=�ݖ��ͳ���Gs�ڻ�vq���ϸ I����a@@��}�B�7L<5$rX�D�x-*|��4$����kGMa2�| ��s��upE���6?�ڔ|;\��T\�����Q�M�|la�%d�9�S5ظ�4����sJ���� �}P��|mm��H�#��D�B��bM��,=.�1�tQS�Sq{"��]��ٻ$P�98�9�{��z���