��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��We����kɄ�Dߒ����{����}w:/�$|�c|/^h�c�4A�|���<�r��}_�����SY���ʹUZK��;_��+��0�$0"�E�D%r6��2C+/S�o6�P�25�z+R���.��I<�%
W�,����\^��Ϟ�4�-t3l�+l}�م����,�[���<%��\i�3nL��:)i�:y�g�Z�eBl-SP�G���9∊"�H@⏊'n�n��l��}��֚ؕL�.?���'�Pl;at�k�ͧ�6�i�K�5�7� �T�ჷf���O�x��!h�:@���MǷإ�q�_by���u�J��`����CԾ�e��=�sϑ<}ci@��<D���I����wDo���R/�$$�|6������AsW���uR��Շ�By�F�KN������c$�����V����)��R�I�o˶w�f	���XBf�y�d��7��쀩;з�su6��WOH!��ܘ_���D�-�N�APⰸ�W�(x9Z]~WYq���ᣣV-ε�r!P���]�s���n�-՚q3f��)����Be��Y���%�Ƿ�Ը>���+?�.?}˟�Y�����Κz�k0,��"�}{���
�!�SČ�0��?(�#��L�N,&p�	P���8B퍑@�9.{������2�[��1r9S��1)[]���L��H�ey%�L`$�w�v"u2�T��%=�/�֓�.������&W��I���ش9�nYW�?�,+t�Z��`�6W�?Y>$Xp{�V�����(tWq��\�Q�}ū@��3�u�)�f�V�!�a{H4^�r+v*��:�!�^�T�zl� �o}����\�@JXx$��hGr��P
�RC-6[����Ь�Il�S�v�T�ik���2��zN�,��T��tJ�U���b�sP�`7��vp�\�~��?k�c[��'��Bs�e���u�>���蔤����Kנz$�i�cE曯=��2���O���"�	�.�"nɬ~�V�eE�rL��݂���U	��t0l��ƺ嫿�W�������G��#_��Ob9k��7^1����/�m�E�+
v>���k�*'�B��!�b�B�݇[n{{v���N>��BW�~���R�f��	V�H����x�	Z��+g�����"�(�O�b��UVĺ�!�;{�6�Hq�P鮭#�j\���:`:
�q�����u;'C�y���|.#���ڊq�jN�ƹ�x�k���hU�1�%oW;�I�R���,J�Ȗ��s���M�H�=G����I�o�7��9Ghz�b�^�Ӓ�nG��Ļخ�)4h�cW��_=�����x�l׸C�f�ӸT��h׬�n��.��2��awn�&2!)l���DU�uÈ�L�rL�&�FR�bW��x/����?א�(�xZVm��W�p��r�E�'��H�$n��њjGk5��)�m�C˝Z�� ��<T �#�;��d̉߶NZH�$�x�{��pқ����R]��_p|�!�t�p6��6��qZ�w�lk�?�Y�u�Á�~��<�-��^v#=��`6�9�Y�r�������}F�{�'O6��h⬭X���Yg�(��C����%!>�6�Ea_Ӥ��F���m��Fpx��n �uget�
��=����7�w�%��p�a_�� s�9����&�y��!f-n�L䵇i-R���Ah^�*��	���BoK��o
�Y��-R ��7[�$Ki$��da�����b'�0i�A��6e�+�O��#�4��t�4���+*N/WЈF?Tu���H=�ro��ظ�m���լ�@�J�tC�B*b�X
Lt�-�d3��J����jsW�$����������5*���T{Ej�����݋^X��Ƚ���5BFyI�)�Յ�Y�+Y��t�\ܥ��G~f��[H���yi����f(��A����_��b�u�����r�d���#�̐�%El6���Ƈq�/���$`F^S���ؘ[�I���� ���Կ�E��^�CC���|S��v���6]���{uR��$o��fY7�f�~/5/�&�j���
���K����B��N"�+�
 ��@�@.�ol�RH80?\4Q���߻�cFK�o��~9�r�?џ�7����Doq<����h�lE����
�B��K�Y�̏l a�mѿ��;��wiϹ�#7A�DȇE����Q���KxP�o~|�솣��q�,�<Q	{',n�5�s����67�p�����6\�<r��bkYA��+�!�ȯ<��v��@N=��̧b>�;�րc�}�z����/+��X��x���k,v��a�͗�_�z���C=o�� �I3�A�1���<.i[��簯H�D�f֍�ۨ ..�cn����� X��b��2�!����5�F�1�!b�Vv��>�/ϴy<o���9��J1s��av�8\�칌y7�c.|o�J�g��eg7���h�$�?S�Jp���9�*�nj� +c���a��H{�����0�(�-���.�!e-��	[!�韡�C�s�"�EO�1�^��r��Y��9���9�"
[�G�^~��D��'�4� K��w���4�AA��9�f)cbD/����U� �%+�&�~޷�����x��� zϵOS{V�V��&� � &�f	���.$�%���{�Tt%�l�J�Qjx_׵k�GH�$�絇�R�`��B��� " �K����	C��xy�l��$�M��=eI����%l5q��(�0�Lc� i�T�#�'�}���!�.V��L��#�o�1��B�����T�mh��ݭSW�Y%��5�#{GVb[
���J
�n-ۭ\���9 m�tE����b#&��F�&�%��n)�#sM	O	�dH�뢀�뙂.܂��k�-�nxN��ؾK>Z�i3� *��H�����+���ݢ
l�|���(Q���V�eTv��@�G�EM 6�Z�L��v�"& 9 �6]3�ą�c�M� �n��M�Є�k�y[���
o��b�o��ΞX6=���J��;�O!p������J��h�%!���§��/Je�~)�R�q�?�f6�����V�!!E���&�mԝMD���<�����"��Ա!����|��'ӛ9����&t3�a�hU�c�/V�b?)���t�v�����/.���w�����j��~����7�r=��1�w�O�'B�i���xW�&���q��΀�m�nm^��0#d7��9a��b�����@!�y)_�z:3}�s�E�@y���t�� !�t%�M���8�0z���JA�<MI.�� �LC�~�9U�'oq+�q��cjƪ�x$�N?��}�Q�M,�G_���(���#�����*�Y��w����@a>i^� 1���*����Lq�G����2B1b��R�B��9z;
wg�#,���͂Q2�`��wTJ����!���������r��i~�z���W���;D�80[�'!r�1� Ff�af'Òm��Hʝ�Y����Ђ�>F���fU�C��1���$�6fb8�l�D��<
y��a�K^���&���%�]e_�kҬ�*_{�A�"b{,./��}��ϕ�N:^���'�ys0��M���)|���b�1�5}u����
���.*">����A�^�����m�Ǻy�LJ�5V�jv0�]�4��
�j�����=ک�!X|��7Jpk�F�o��xL��斞y-��2�`�̨���F���jH���0\���}����BB���P��px���"�&Jb#qxF�����%��Ϥ:��
{0��^��@ʆ���g7Q-)Zł�V��s��w�hK��l���(��0�5��h���'bR�VT��v��������?�]7�ӆ`��)ա|7����A>�^-�"|g*0�AY� !e�X�]��}�V4e��-R$ܽ���G������_�����WM��7�b��+����#��6y�F�<	�B��`p�4��̰1º���۴�x(�"?�jP�	���i���$P8���Uױ��L�*]�\�Ci �jӣ��d_38J��&h�6bdc�y�4PFz��i˖�@*T��i
N� &��&`<�{x�mޫ��a{EU!��J��Z+���9S�p1	����XQ� q�����o�Ԩ�L�NKT31���|]�y����1� �*[���V2|_��`���;6d��
�$�U�����HD:4��8?��y�~��-���ԓ�_i�����dv5����^>�}�J������@�V0.�+/J�yL�m�l&���ϟy�B�aV�������m����F��8���n.�v�f�/b�r��*�p����	c�T�n��Q�F�����V��^�tG��K�ČMtl���n�.���z�7Usd��S����A��T��<�'�([���lT�V�Ė~��;D886+��V��u<�e[�xwT�[��Gw��X�v�>5
)s�O�\�+�5�7��5$��'�Ҙӡ��KŞ�!P{A_\?h%�ݺ ���B�}Q)L���C�0�t�g�x0�ұf���qMʣ^�����M�d�޲m	y0��?�ߐ�ܯQ=��T�;zK�L��D{kΆg��z��4p��26�
�^� r� �h�q�( Ad�s���Wr|%[�B�":-��e�7���颫Ek����F�θ�sI�V�� ��ͭ9C�.�<��t ?̑O��0}Yc;��$GD���-S�G�Fh���p�o����M.�ρr ��� �������U�"��"~Ũ����4ۙ��֭��D�6o�K�L�ύ�H�P��ۀ`Ӝ�I�K�:�*�Un�����*��U�w�g�{}�Zb���O������Q�?�r�ʾY+W�7.%�CT��.�����`m����	�_
NB�$���@��i����ɧݧI��<�d	��|x�H�N��>L�Czv�)�}5��/R덍(��M��Zm�OP���mt�'��e�X�%�1O?�
!{4�Y��ؤ��5-�����ܥ�ච�G7��^X҄�N�������&��y�*���u��L���:�bo��9a��`���x��	�" �.ܙk-?-�4,SR�}a���W�x����b%$�9ᙄ:�m�l�O���/˃`(�`r0Ao:���_$��ۄAa�3�#���K�,!4�+�JG �+��C��q�kL���6������aV��uݴ +f���-]�g�?�Y�'��I�?�b&��,
��L-�R���9�<Ќ�.!{^ع$���+�+ �%*x���I�Cv��AN&�}YUB��ߕGS��v!���z�$UH2�i���vT'�?���]%?y���I��a��ܹQu&���[K����&bFg��t�ͫ��1�NҠ�CI�=�7�}.hğO��W�yO�m#�(�%'�p��n�;5������$|L��:ք������+3�q��n��(�e.�O6m �B�U��(�y2�$
G��p��-'<�C�����j�]��KYq*����Q#2�L��J��?aH�'K�m�)�ˋ0
&��0��s�=��B޼�?�!�%���et+��9_NUJ�X��������{�44���w\ag9������Ȑ��bD'e���"��-o�0��Bl��{�;WzAo�p����3���3R�B��m]�x���m�MKP�ɥ���C�h��x1���́E�i���fh���*��MnU�<Fj�!^�`��|�g�x�N��͜��ͧ�/�Ԥ���#^�sI��'��>9�{!���E!3G}�Q�\ZC����ݎ�Jm13��y��e"w�-Ă�w�v�q���s)P!zf��������P��|�4�N�����gV����pS(��sɩ��-�=.�=��v�{�?sTk�E�W���M��懱�txp����>���S�jF�lx��t�4>Ԙ���/C�/2�kQ�$�"�����]���oTf���i��X�� ���/@Xج�$��v��M�J�5A��Jt��]<?P��>I�����d��#�Y�]^�5w߼�c]Co�������A���8�@�D�s�&�QT�R��m�J��!�������R�kg'5	ᷴ	ҥ�~7���CgQ{J��q���z;�ֈ�儩�ro���嬼��t�����x��NR�/�
f�&�x������sƆ|*�9�����Z�%��"et-͖F$�ĕ7�~�ѠZ_̥�	��Z�V��� H�9َ��e��Ψ�s� j޵�-�����h�Xiz[�\�`�]݂R�k ����(T�p\�%�TaRGOİ��i�~���>�1��[�wѤ��*�� ?٩��M�>x���v�F�q�� o�3��x����(��O��	o��_��%�-*��6s-�~S��+�T���#)���B�Ō�,N����3An�'��;4R�C%<��P��I�Xd�B+����ӹ��kN��S��;�<�^��n/���Z%Z ��`�ևl�Z���(���F!���[Hգ���#RjTh�OhN�A���Q����˥�s�䬪���t�$7
���F�Yǁ!7�ٯ.��YO�O�Č�js(�.I]>�7�'���1q5>��)��|3��ߋx0VN&�ר��<1r�:�>޷�R�Ǡ	ɼ�U�Oe7Z��.w��{Q��bHa�6j%NP���t�G˾\7F���F�I-D_ S�B�f�"ȓ)
�×x5��L�|3>~Y?�-*o.��{M����\f��`7�aR�dW�xs]`-��s@-V�A�!�(҅�(B"zg�S0�C���/�?h������h�M���b�No[� �ڄٚ� ���"�����M.CW"�܂K�±}����_\��ri�C��p"Dz���3��"�{��8|�d���$���������n�-��
��;2ݲ�s;�\
�����ۀ�qP�+u���`�����ٺ��Tn�h,-���v;�y�� ;.�q�P��2�>5�i����l�U����*��A��'�{���Pn��j�Q����N���r��R1nJm[M��	���̮`<Ba�� g!d�#���}SZ8�:�&]��ũ+��w�㱬�����u��fNM��U'��җ���#�gG����I�P�/th:7�j6C��-�(u2��bŵ�v�}M��l&1s�8U5�Ԗ/��2� <1��ȫ�^�a��{eW���V^�, �����2�$f�U���Kz�$2�����s�?˦u�A�Ěg�0G 6�-d�ϣ=���o�Z7�/,"��1˂�r��
��DHPܨ5����P��b�~��F�	���>K�y~�zh]K�k5�
A��Rj����#+V� ���ۊ�YOM��p�V�������D!�y����H ���ă�(a�;hY�^��H޴������Gp�ƛ�{
�k�;�d]nRv�wY�^M!*�F�B����P�&�B��eq��{�v�2�X��$ϵ��eA�@�y�����U
�ЌV*�O��Y�͎8F��|��d�B�G2Yq?����G_S�2�O@y!Q��jyJˎ��f�yuP��KB1�(W��#�`�E����q�Vj����||�=�9a�b������(ƚ_۹���`u�N2�	ط�E����ZՐV�k��D��-w�*S��ޙyQψ_6�+��L���d(�A��e���c��A����"���v%o�h�Oq���=/�9���ߊ�F=2n1���'��V�,T�@���	�����<\cb����R�PV�Nn���[+dXs��J�5��`�a9����N�X����X�'�B� ׉���-����gQ?�hM�|\&�	oXir��[���o �_�� �BB}����(�Y����#�%�Ρ��˷�o�V�[�#�������8|Ρ�uLy:if
�߾헨�A�!����8��q\�t�_2rdϯ)_¬�T�\�M�wd��i�l�\�M��C2tt�\���v7��H�{d��@�:��Y�X��+B�����@/zN��ޓ�MPm�kyJ�ޔ�i\V�)��` �p$k�ej��n��e�$VI�q&KgͰ�B:
�A����?�>���d�(�Éhמ� �M8���_?���"R+J,؊��|�Z���þs��cƸi(WGCPhb��јIh*;Ψ�y�U����ۂ��ڱ9/Y��~�9W�	���������͚5i�#�l�%+����vE��xyD2��p������&�����
)1�MeU�Y^[Ҟ�я�u)�wL@.�G��x�p�̀ի��B�x$ ����Y���a?T<�ب����w�=q�~�̠����L�;�Q���=ѠDE4�ÕE<Z�H�ؿ��̕�m$���%�11����㾿�0l�V��'���S��s�{���1>�m�E�C�F�#3�E@�>hhCܓeto*�]�|�x+�q4�P��e.l�{�L߉W�D�>4��w�������V�K�<�ARGq$.e]X�w�X�����mR#�s��\��*�o�zI}�Pm=��7�ה����n)�K�96��ي�BI�R�������U���L�5�o��sSN�꯶��Co�-ߚ��9e�WW���9 %t�)��ΰc����L�{2=bE�ql��U^����4=u�[����K�����s�*��&�
m��=|bv�4n��iD��`�x3���&O�8)`��d+v,���� �����Ad|A %%��U�&]d��[�f��Ϸ�`�ގӃ\z�ˡ�������[�;�(��$���,�1�zm*_��]�R�ޒs��~/ܹ��$��ѿ�p�J�
�!��������W��i�9���E}?�`�o`�����݌��LQ�_�_�K�.�Z��v�-�Oi�V�Ĵ��kGTCsl����Es�����.B�$���A�����ȏ_C��>��"���$F^�D���J� |��`��C��બ/�S��1��L+�.���V�voJ-ެ�|�E��[��@L���n�݇6;��ҵ���z�!�_Ձz��� ���ku�xmIW���t��^��o��j� 8��ح�=jCL� �u�c@�i�,wO�it#�����2ЪEj��Ό˶|D�⌛�r0s�\A��L2�{EHθ�-���5�[6�e�2t�}ķA�@&�jf��7���T��9 ���9���/U��7��ZC���c�x4O7 �����#�y�KW`3�Ӓ�Z/�B���f*�}�9���s�� �f�mtk1b�	mI_�G���_�M눰zdݞ�`�] �߻��|��Xa�Ju�72k5���=���� y�'%�m���S��+��y��3(d��N������2P��#��v�6�O�?���"���b���?�(VHӶD�~�m,aO�� 3�pt�Y���*U��`��h��j�X�A�o�k�ɳ�r�EE璴%qdݨף��ʓ�b,��(�x8t��W*�̕��MI�8rH'�u������9߷�.8�~�ʡ\	p|�e's��Jg^�"[o�p�M|���O�5�%ň���ܙA�Y�F��׌K�Il�+�%svcY�8����dt忆P�L��H��D8P����3��]��7[��H��-�Z� df�ݑ�{�v~]�]$  ,��h���3�bA���h�|P7Ҙ��#����F)�cӜl���^!�y�����\3WO�+��\�g����Tف�����@�<��^�[�C��=��tU� ��	��S�Gn�����7ւ�=ouX���*m�U&l�D���v�ʺ�6,�7s31��)w���7�B`	�ŃU�A�iQ�C5�X�=P��V�����$���:"ǌ���~�a��	nK+����UB��#0��F�} �h�,X^Л�}�D�� ���&p 㟄&+s���h����ܠփ�2�s���iQ+�$u��2~4�EŐ	p���x�:<V�}E ��Rz:񷃫KZ���/�X�r[���U�[,+�
D��9�t�v[zHo�Ժ-oH��9~{�f	��./�u����,uH�dt˻ObCTo�d [�����N��;�@�|�����Y���~�Luwޱ��]i�8>��k@ߒ4�p�Q�_p(����7�-�IM�P���>3-5�qL�#Œ��i�C��*��Fz3�%�1>Б�hBeNK�"�EN�Qh҃3�F0_A���.ϔ1�`�W��n �w�	�<~��h�ѸE}�S
����$�u����������w��p�N�Њ���8�z?z���<w�����p��0�S�c���d}K��n�N��`�h��=s,���f��l� �C��#13�>�	�J๨��_mX�o��{.x��b��T�/�׃��`�]��&�
�Q�	�b��K5gi����p9��\^t"�,�D��7�lS�� �Cc���3f$=gj��I��+H5�s�����ˑ)��l�nuH���a����Ie�P5d0���8�i��҃��Nd4�( ∞\�p�6V�O"���)�Lqy>�y�D(��~ ������1��Zpe'bV�E�dW��mmF���#����ovQ�@�۽\��iE������Km��������* m�hA�����=���;n.y�'���T�˯�&IpG�����vY�rɫF�W>�rK(��[w�6�U��i*�h�_Rf!Ø�hF湰��c�)��P���pm@}y�g�`gI/o$��\i�z�e+�R��h��1�ct^���\K&~^�t6�c|���v�� 7p��+��Gl o.,�����Q�  ���q!��z��E��2`3����n��={���T�]"zu|���2lȠ� ���,ji�I�A^��5 ���Y^�t�4KR�w���4*�}�dq="I��;����i�"1P���T�;W��D?�m@%�%�kɾ�C������3��n'��Tx�c�/Z-Ul\