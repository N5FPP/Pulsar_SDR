��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VYkM�#j>cSdw�u^�CFMr�RI��
f8�*�ˁM:%��lz��rg�[�]��hJ�-��Ǚ�#j��&v��LL2�N���?ş@'��# ?��}������N���P\������Gу��ހ���H�q�%��y�S����I�T}�m�"�:����nQOۨ���ߏ]��B��ͮ�8w�^RďBX�Tl���&s�,����-]�92�J�$b�!�.IL��C��zHՆ��:����`掌Sk�O�4;FUBTG���C�+��k�R����1b�N�I��G�W����|�p�`|���KPNs��Q�{�N�/IVy�k���C\��������h�Ϯ.���U��~�!0��":a�]j�Z�I�3������2����7��I�qb���.^���t��5M��-w���+��ǁC�2%��x��8���{b:&��E}i�Z�����=.�Y�q�b���,�{jIu#�q"�8_u��~\K��p��Ȧ_��n�%5�JH������Xϛ�x�7:IfU��8@��~ų��^rN'���lb��:x����ݜP4"mH��?M L���*uljm��V�I7yQwu_�^�F������b+�yb%�P�ذOZG��Wkֱ_���0�8~�rn'Z1�u�0nH�9, ��k��|����^P��V^+�^n�
��Ϛ��f��C��7լ%�B_��ڗ�v�΅���{~�>�BAA�"�p�bg�K C�8�K��e���N��,�W��^�b��0W��2�pXR �s��x��]���Z��'��\	��r�D�ZɕBD@te�ڠ��+�?%)�+މvX�T*������y���=q'7��҉��K���A��S.�BǙ��.�n�]�Ss���qV���S""�w��p��9n_�;��d{Gy��{���o��YP��K�'���S�5C���ł� ��|Y6�3�68<( �4�MH��qv�P?;�F1�����l h�#>���u��@�_�Ih�����KT�5���G)n�����ﶺ)/W�H'��Yι#�buʞx_��\	���!��ʂ�1Y�L�&�=��hD�9Q�X�^#Ɲ+���!}�Oh�����űԘ�E7�&����ç���4F�����W��6���ۭ�`1�k�ڽ��@"�Bh��.ϒWv>U�w����P�Z���� ��ٌ��e����:�:EXҤ:�xȶ�?��&&��i�Z[Gyc`�r���ѩb�Ca����c�˅�g���V��2'Z���&<e�{r�fܺW�����[{$l}��L+����p3�b�q$BEC�Z0:\~t�_�c��Za]
i?7�_�!��>$�s�,�(<��=��)Js~���5>wJg�S�E����dLx-��O��۳�{�)�h��/վ��5��u��``M\�gBzVl�����B9�{dlI`_7��U^�,C���]y�͸ܣ>�@j�� sy*�rҧ0Ǒ>J���(a
�M���W@Z�,S'52�o���+bnOOz��s��pw��1�9o��j��L��)سL��Ei�>�������<���KI��z�r�O��zm���f�@j7Nؘ[)[��[S�=�Z�QR�C��*oI_l�k���N�3�e�>��Ē��A��U6Bf�h{f�>��q-ph�?�ٖ�u
��~Ŏ���@W��������@k���3%��	I)�����c3σ^�CofhԴ$W�r��z�L@���ޗ�qݑp�NK\��Q;�]��?-�G�L0`��.�D��]�B$gut3�+!m��l�r�"��VŐ�*�W�g�����g@Me�Bx��Ue:����D�u��N��˞6�.λFC|����<^/��� ~�mD��By��@��6�">.�3*��VqR��f�ːr�s���N#]�{���#�Ց0����8�&;����q����J{�D�y�-��#�� ���>�s��C9貭��F�iI�q�J[�NM��h�i��G��:�[�U����̡�nB'V���@+8�'Z�x[VE�0�W��M^�����&����DClj֑��QrX�Y/E����E��2�ƻ�V�A���jӪ=�2�@G�L
��mJ��-�Z�ɻ��,+�@S���Ʉ[��Eǭ�t���ϭ�8ǖٚrxj�ag�4����}ȰO���/6zʭ<�]ϙ:�ٲ���¢�@tɚ��(��"E�w��+iO-s#g�qwoox��Z�'T5�]r�o�X X:��#�Tq"ΉIU�D�����������ې��JO�@A�?�yU֙佔����H�$�F��0A���o2��M��O�̿#� �qI?be3����;Ġ�/�f�r:/��g��$�oMr+v�|R�$�����r����#�b��U����F�"lu&�@W���w[���07&ͥZ��.I9�.��b����X]���{�����A�gnuH%���vJ	G���w"8��$}�zͺ����@�ԏ�Q^sT� լ�[p����>i��3�&/dI�W��%yW[�D�(S�Vc�s'9`��@_5}4�$��OO�n�acP z����;�C�iX2�'�3�Ȉ�����M|[�V�>��$g�d����W��w�B��J�v�[{q%B�#YNV�dKi�ִ����#�ǐA+A����(]u�J�
ۢ�M4�!�& ��(c�,�Vm���9�Z�)K�l��7�Ӈ!�G�3�/�A����%TW*޻|^���N��{�T�G�v�+��S�uU�4��w��P��i���<�S��]��㛐��?����0
�:#�Կ�SvF܉ax3L�f?g@⪹It�Ò���G��ƈ��}yۈ�j�z�C��>��e)PH	3�(�NxCi ���3=<��Æ\��kO8I ����ϕ_N���>o�fA×����T��qr�ǧ� pg��$�KQx�m[�ݱ�Z}uK��,/�(w_�!����!�j�D�z��)���'�Yƫ��h6Π��L�YN�Un(��H/�X+?�W)s<��H=���O�/�)��Ia�T5;~��P}P��4�?�s8֝<Y3DҖBﳋD�~���ez�v���\�5�����͢N�-k�>�'{�rF�L]����q�8���z�%l��$���x�f!C�U�δݣvpB9���r�O��iQ-�j�q�[�bE����"B�0�$z�Ti�)�F8:�j�Z̰� qvњ΁3+v���址O��T�\�1O-O5�aD���6�Cq�a��ಢc��7���i�L�%�H�w��j8BJJNn��U�f�ns_q�J�`_�b'=��(/X��14tmz4&�oN�T�����ρŌ�[�������TE��8�wBpBw�'l-��j&>)�Y�Գ��A�C�K�S��¥F���-MK��-�v/�\�U���ﯟm&�hWѶ�_���7��j�]lt#���}̯@Ť�����>��S�d�0���)0���25��x��u��A$wj�?~��uL�w�z��D-X�O�k~�:��1��!�w�1[p6������rkH:���('9��BK-�����#&f�����y��e�|���ĭ��,��hx!�E������it�}&�X�O�2�ۼ>Ѿ�`y��ɰi���X���^��D�~�lk�Hh���r7FC�؛AȪ�vVR&�0a�QS1R�Jg��VK��Zf����J�p�JysM� X�@�`��T1�l�x�j���%�HU�=�~��iOX�ZA�L�8�Z�E��@'#��ۣ�`��-��M���؏�bh?]��#��l/tvݮ%��*��Rݺ�+�P�n��9����t"���+����g�P���ƥ{(���z�V�Xw-5-I~�<R��cD=�W(�y )���ɋt8nιk2��2rD�L!'��-�5���i�h����E�]u922.�_}�vGa��<wy{u;���Xu��J](5�M,�4��Iv��87{G��J̑�6a��։W���:�+�\y�1
vXB���c��&�P�v����z���P��U����R��5J��������AY)y��!ҿ5G�~T���S7(��U<��Vs���oAu���.�_p��YtE�K��kJ��Z�
&������X��yQ�&�o�m6Y4�����8���U��n0�p�^�	Mӯk�UB�nvR������ᕒp���8� �QӋ<��s@k�%�:U�f�~�
۔P^���1�^����U���@��������h哄��/}��ñ��Y��9`앎�3йD0pȨ�38�oŰW�g=���M���Q��N�
>PF���epԊ�?��b�j��������	y�񌪚6��o>dX���&�g�P͗�Z˭����<A����8�癗C�,�x#4X��~$pA!�Ȯ�pf/��!�nU ��0�ۯ2�Cw	,��>����Qs�����v7�U�ȕ�+1KF�6�r�H�b��1c|	�������m7��!��ծd�X��1I��	�>H���W��u|_�I�}��`n�A�\Thܒl~t�r��2{�v���6�w�s;3��==V�YE�3��k�d:�OH�٘e0����w$�~��=�R(M���j����H(����l��ؔ��_�w ��D�T�?���A�C���A��k��CcP�y���zqJ�Gײ�����3"�t��GゑE�ׂ����+��-<��y/*�d�xC�y�r�y��gO��W2'���|-�Ɯ��y�I��W���� A��!���KVDΞ,s���P��m�y3.e�(cD*�+m�;��!Si�~�c�vB��a��ޤH�N
�^k���:u��hh�d�eι�ZP���GWB�et+�Z�(�F "���\��R~i���f�;�spl�ٟ4x� 5�ב�e�"�R�
���_q���Ԅo�:e�ՙ��;�,r�d�i?R�4�0e� ��]@&V)}�)M�h�z�2HDUs=P�P<F!�a\(t�e0:1A.2���"Uos��صѼ�����0x��epI�/����QT�>��g�B�
�{�;��O�0�{c� kp~��{�!���D8�rUe�#E0��-�(m,�;��x7)8����*��hj@z��j7!�)�����YH�W�C��]* �\�5<����f´��a�։d�}�E���JˣE��Ĭ�U����W��\�^!C�ܜ�\�wI�A��t �S�?��-�t�o:�|pG�e�-������_�;̮�2{�HJ�k w���#��lH��wDz~h����x(1p���j晿�slK|b��]����4* XG�u)( ��Ϭ��7���GZ�O�ڵ�6	���9z8��r��f�*$	aǖ�)��wF&�~�<W��T�4�Ba�̽^����S��=���츧�ˆUG̼����!�mzcW����p��|��Q�6��	�SM�=l>Ѓr1��2̽eL:;;�w��Hۗcc,�	v1�����.\F�K:pR���ڣ�A��
��6eE��v�iɞ:��/��m�َ]ܓ�!���@h��lѨ����Z��#�q��ml�Ό_�-�`�MR������7!-s��������M�"򿦿���`e���׌�iY�S�9[虌�	��?V"`?B��IHi�p���Т(ؖ=N�y �xg.�0�8m���9��/1#�H��W)���7ZMH<�rA�bz�m]F�.^�uj|�oEA����FkTT6����.Qh�"jF����[U�Ga�D�B��D�Y2 `����!Fr[��2�Wb.8K��$�<�Ʃqz��c����uWws��b����Lun"�:2��ٯ�F�q��[ʎNM������+g�c�R�,;���2�{nY�X�Ҝ�lM�нE��p�pg� ��"�W���A��Ǽ�� H��[�Xi�`͢9d"-�V"ٌ��.���1t�҄>8�ρ�i���x�(��f;���r�D�g/�v�^{��*����
<��U�NFK(d�/! ^3�ӴP����A�Iu���x�����bʫ�"?��G�
I�4��"H[����V�QOqn�AjL�,Y��P��uO�Ӕ��t�[ώ���#[�#)����/�-K�'��i��"�l�!3=�ܖu�YBpf�����W.�Č�Nj!:��7 �v�������Nr�*]7�(L+нRG�Ӣ�N%_�Sp��ds�.�F)�X�lh��J�W��0�s hAnp���O{,>?s����?��Ż�e�8��q2�#^������t�R�rb"��G�r3��>����OǨ	��I~s�	3JF�`Pgp�:?��Ӫ&�w��YIRp����u�!�Ijm:8�D����/&q|��-������@�)ő�0�*m��xՇ>z�8�{w�;���=t���[�p���"���3��9�+T�0PЎH�C�����__�5A�Ǐ�/���]0e.Cm[ު}{�a���xwR!�k��^h��O���>vf�߲�f�d2�*G��ފ�Z�ǟK�~Z�3\9�����ܘ�d���έTqy�!��	/!�d�N$��:�cyYC�p�y��ֵ����.ʒ�'�ql+1��U���<�eIv�SJ<rXF!�!����Sk<)t���;d����^z��a*�B�;�~�����4q��wQֵ�1WJv�n%ϒq7�Dk�Fɦ�c���e�3��!������*��:u��V�5�p�E�zE���l]��$��c�.���M�Fq8h�FQ��5�~�x�j.6Z@ɠ*���MC�K����8�)c��1T�����73-ط����S�KX��5��`(����j(�xN��Y��
�F����'y�vՊ#�ŸD]ԏ�9�q剹B����yT�P\�֢$��?���.�RZ˛y�,�H�/c��N6W4V��\l?����Bm)��κ�=���J��w):���>�Yl�1.����r\"��%
2��|J�$&V���{͓����L���t�I�I���m9���Uv������r#nzu�טk��Q�$ve�(��Ot5���sæ�n�F���a����βu39Pv�����܅<��!3��^Σ����j������)7�$�H��XQʧ�����q���t�6j%�����8��*Jb��ە��!5áT��N�S4$g$'G{���>3|]|�
�	!���Z�+��6U���nS��w�=q����pJe��5H�#�C�&���c';̄#�����0@�L 1�z���BN6λ��{ݔ���Ͱ�㭟ï�v�2/\� �e�"ڂ�l�Su�M.�0�e��F���g��0�˜9�P�V9�|���9�e�q`F�rc/j��)��o9��2�������q�%�v%� r1��5}]I
'S 5�
���؟�5r��Rv��)��$j�}R��ڶ�u�Ь���[i��Ty�8p�М�6J�mb�������1�+	:����9���@�{{�+�_�م$v�i�O����N5�`���T9ɑ}�ZW�غS��7���1
��a��ϊՁ��e �s/YӰʴ/���5�?I�|ah�i�&Q��_~>d���P�n��\���z�/$�(�?������4$�p�e��8,�=S�M)�>X��W�&׿�I��E��
��l�<�,y6��|�����*<L{��}
'!�ݫ��[_D���_;������A\�J���wķb�t")�{�ı���r����Ƽ�#
6�>��Q�B��vJ�{�Ǎ
asc�T���d?;�4Ĺ}��E*��$��/({k�I@(�iGֿ�X���a'	��Õd2
wՄs���c»ѡ��Yo;�'�=�.�E2"���9�^e(O�`@�[q�5ɀ�"t�Q@�a�0tB��V3kR'ܥf���y13�G��Z|ywK�qL�UO̜