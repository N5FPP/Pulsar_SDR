��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
���ۇ��������)��T�'�L�3*�51?+"�W������7���׷� Y�[�}nP=�PyW'���J14��qKxW�୽�V����+)Ό���-�o(��Q��`�`߱��H=%]�ȗj�u)9P��?L\�Y��rq�+W�||ꅡ]����Ҿje' �3��V�K��4���M
j�t�҆Pd�{�u�{d?������կA9�O��[�&�o��ʯ��j����Ǽ��Y;`�=���7B� M Ry��X��[�/�����f�E\
�`#��qK �T�PM_�?����w�/����S��Q}'�dS��&tZ�l�ϵ 5g���q�}�-ft���]�..pх)2}��d����[sH��;��D����џ ���AWBP�PJY؛U����6�?U	�	�0 ���_K"����_��m��T
wy������AAG��ӯ��`�t��"�r͢u/�4��wj�l|�>�h��㉏��c��#�8�g�{ۇi:��?
�P:
�ك��f$�F����@��P/�DH��;�f#@�LjaFO�`E��{ �]��N}o!��M�m[�~s�"��s�p��o��*#�q@��(��_r�����h�R�҄hb�U��+�7��p��ɚ���xWs�O$�r��G�$Mϩ�P1N���	k��Lb��V��y��Y@�

���͌��sa"��`&�X]!�'a������0Zepr��3���U$QJ��{�Ѯ��Z��a\F'l�;��?2��Y���l��c�.�2|�>�o [\��*#2WSe�W,��_��7l��u� �'z�<� "��.��sn��{��O�����^�2>( ����3�#�Sp����5�q��JpgQKi!�F/��̠��lл�-� ��]���6�օř*2kS��h�o��$�����p���Y,��>D�S��mJ�5�d��탮��ë�n" �M����]�j�Lk,�=�ȏ
��?Q��У���3��I��K���7��c���c�%,C��(L���yɶx�$P&���Y��k+�3_!k@��	�LK�Ӏ7��إ7�f�N��w|�!�T��9w�[�`g���e-j���⚡R&<pF V7tZ����w�c�ei��T>�D�U�I].�0��6�%�4���y?��(^ލlu�[����� #O�+H��{+�-aL�d[,>Y���:��S�-c9϶`�J�rjYoL�8�5q
;�G��bўf����7���Y��I�Y��7�ɰ��V]�I96BlZ2��E�]tQ�풉���� 
UAL)���G��Y�U%-b�4>O�d0+��Ta�-�3M��(�m\@�lco�TV�E;m~����'Q�������+
���P�W�������s�*;܇q���i��U���4�=z+��f���o �YO�^�\�g|�_Bi��(�� .�9Jy�S�=h cU�����Mw�7D��������A(�N��h��l_W�X4jm�ǔ&S(-7G�&�Z��tg���q��*�οR���q���a�jv~7e)�R�q	�\s��o�|=���@�Y��jЩ���hS��6�pG�N�*8v������<Ɩ�U�:|=I�g*%�1��X1��b���{�7L�aX}�z@��<�t��&�r痧h}��E9�<3�ۆ���?��`sn2��M8���qqNm�l��������&��mŐ'O���}��ĬCfd��uOhX�-
 ����;yJ{1�6�Z���	�?Bm�o
���Xx�&�<��yl����Ghb��Q�R�z߿�	�ҢßyV�ʰ����Bg�l���a���rڿ;��(����l+Z�q%1���'�WY��5��n����+��B��Uy��㒖�Y��H�՞eK�̔�U���/ B��
���}:%*��l��0�
�+m.L��Q�;-�zJ��em%�;�]��HC3		���U�@C��J{ޕ캋�@�k�ߤ��[�uߪ.tG�~�Io>!�t}�O��� 9I��c^�F��b���-�哏�,����p!C(T�\y�A��l0�������@p��/C�-��(�i�_4PW��c|�����	�|.�a| � ~�o��U	I]1��k�����J����p��I�P�{+G)(�)7k=��Mht��y��f��w
��yL@�o��1���ͳ0n�b��n	J�%:�3��U? '�ө�;O��bF�}�����V�.K�T�����S��RRߊO�]�R�C�Q�	��`�K JH�*���@o�U�gV����sUi�9A���&��,��9�]�)g���~�A�D��!�7W�����J&�@W&��L~����&?��H�z&�Qέd���D>�<�?�'��_�;����k��(�8���I$���3Ͷ�a'��0�u���W�|�g#*���a�m�N�맡�|�DMmR��<��K�=D�Sג/�s�	�KO_Do�_Ց�N�(�-ś��"&&X���F�k���l���An�?��3h<	��WZ@�WUm�3~r!���!_�T0�d,t:E�
Oi�µ%R��O<j~�����BЗ�ήNW	���D'��1[3K���R$��5�~�	�rY��&גG9��~��Y�4�{I{��`��3N2^ ��_�%z���Q*̃���h��g�5j,]|h��`a�sg�����W;�p�X[v�}$�����xoj:������+�3�8^�-�/��D��� _/T��i,�.����0ˆb����G8_π��"�N >�g����G�<��M,y���z�g�]^P��k�)�%���j?����%�%��aBOR# ���?>�pT̕ ��G����8�ʈI휄�����(j]��d~;y+�y��m<��_���� %�� L_��<^^.i��S�xS�Vwz�5{���t�eR�Qw��C���H;�����w^�c0"�� �Ȇ��c��7�zG��"���ү��^�9[{J��J�׈�V�3��W���j���u�"⟕�����"|{�AGW��EOL����#
fup��I�*+3�����E��W��T�ƮkK`z0=Ӷɫ�xM��h����>�ATAH2�q���o|�n��J|�'�G�v����4�����_��Gy�>�@�q�����"�j@�u�*�%�ҹ-Tuo"^��X���[�c�ۦI{,ڪ�Q�0 �Ĳ�}ey|~�5WW�q���x'�[�!8S`ˎLA�A�p$=�K�E.ya��r�'��R]ߎ���M�$0�rt�(�=���r���J��oD�@Xt�
2:��W���}NC�e��u��+[��*��7�yR�Yq���c�XT˭��
E�{jാV��/
�NZ&�&�{'q��L�Ó�3�ͭ�ŋY�41���{Ȕ��"�j:�����}�����_f
�5h�{�=�$JU՜ٔ�G� �k֩ضU���agT���MW�� �l�֏ى����½K޾~�πKe3_����eL�d�mR��wA�wM���C`���m@m�6F<)`c��S��D����@�\���	��o���8h�)�1�Wvd�,�zj�Wa;0ȴR��K\� JA(���J��N�
[�Hl:� �Ƀw>$�x�'��:Yj��EM��{�e-�{kI����Y����w�=���0ܝeN�;����0��~�\����A u����XhPd�ٚGf��e�@�]ۉc2w
>P���n��-j�>
��G�(�v2���e>F��"��k!�K~�Y\HV'3�͝�"�1�n]s��mw��!��mh���w�ZfZ�]<ۥ�1|�c=��ߟL%'%$=l���7&ս����ږ$�������EHt̀~��H<\<{:�!�֡�y����TѰ�*����E��$̖�z�Ոܶ��Q��f�'՘�{`�v�QB��_C)�p�l�}�,.�=���c� E�+��ǯO���0�%՚�k�^��b@��b��T6�F��}:��L�QOb�خ�c.�X�̴;��]��7���D Z`p����S(%���Y����xl�d�:����T��Ԯ�?]�����V�xZ���\�W ��Q�@��ȱ��-��=g���D���*F�t�ziS���u��	�Hq�����\5(�jY�1υx'/]��\����F84���p�xw�+����oXG������u����ƙ��HHj��Y�5?_d�A�ňX5��{G����lΆ�xw������ٝn�0 ���W�1��N����<��l���L���'�}q��4��0Im�����K'�)a�"�<��H[9E��ˈ.B�Y9K��1��13mGr�S҈M��5RKU���@ת�W����U	0 �^G�7�J�k��G��,�'��Ɍ�N�d�1��>R�[�*t���?�'(l������_i�'�5v���h���EB��R��V涸�< ��<L�=j��@�:���X���KI�-"���!򙅌�ϰ�kCv�G�S�p_��5�� �5�9l�@��D���t�?4|��L��B�p{�a�����[39b�BD�<��⦬*����M�J��K�O�3��]I�0�D�5�Z�m����7fY�S-]ϡ�����8�.�D����6�
[���}+�4N%��S�)��^�M���)�#}I�#���077@/(���R
l>�JSsL�{���%�b87�/9r	+F��ݥ��bN��B2��^k^A�U� ��Y�yyZn�I�pN���e}�{���C��=����O���Y�J3���s�`��}�ra�����]�Y�z��R썣yNL�_���¹������v� �Hmm�eS�Ȁb�pX��6[�ӌ`q�Y��;�H��HՆE�W�b�K8q �r��4ѕF�a#k��Y,V��:ib�����js������HH{u�8A������:��j�r�TH��?��*9{�A�'���OE���\��x?�#�T�� ���sd�>���(�]P#?��^�/$���n�8jF��� �j5�_S.OEJ�&}���D�sT�ꌉ渔���u ���{	W����D���{N�?�-�/� ?:`�)�	��gKn��c�z\g�kPK�%a�[�E�z�rR��d�!�[�/��Y��$���U����rs%�r�w��#Z�Nu���~R�����7��~ߣ�/`Vc��:��Qqg����@��'��k��.�C�����l�F��n9���"��e�#p��Љ������ůE�x;o_d�7��A���O����0��� ���7��/+;ǳ,r���ó��t-c�U߽*�k�+�*�R4�<t�	h����h�9<����zAwH.��J�����~��ud�姙h���^������m]*����E݊�IB>mj��Bd4��)Z~t�L�2zW���uf&�P�������u�T��N�
;x߉�;)��&����jPtG���Cq�5�L�]�&�Sw������
���q������p�*S��m��U|����/�'٩��Z��ur�(������0��M�þ�ǅ5������5��7��𺛶8�&;�鲼dn�*{�Һ� fbN�ZD�]��7��&���\Ρs$�N�R����q�biGrv��ID���\]|( ��A�%��Mx�j]��Ք�6��y����:�kj�78M�{���&����I��!.W$Z�u�O�� o�Yi�zD"#�M�ͬ�_, �S1�p�4��o{b��Ly]�Em�W������;H���G
�I����օ�A�H9�9� �=��u��}q-��S:n-�U�p�D4�Z�Ci�ɫB���
��h2xZ��7��eB�!�Ϲy����q�7��bNWDV��6<4mG��VX�y��n�`�Dq���q�`�3<��.r)��_��3�l���/ؤ��l7�����(a��T[2�\���} �|���-�|9/��M�3������L��K�P�`�������&�k�0
0N��Zt�B�/	+6�a��31l[u�hB2�d�N㶛Vy�]�ӝ��ѩr��'��oQ@p�1eߔ�8����� �0h?�f{�����@o�Tn�R�� }���ξ`��Zj>���)��������-�W��P�l�%�`ͱ�zl�k�C��=��8�@A�;�vfs����a�K��Ps:n���3!����?]�|>��z��&U�h�}��VOyE�h>�V�k�u#ỿ�h��EDH�ĵ��]O:#��MG���Z�'��畠55;����Q8Bt(�e+�>��N��t+��jL�e6{��e�����3�g�+��}�Y��F���6&�� Q��n.@Y��34K�^Nj��������_�������V�ջj�kn+lR��|��e�i.�Q�����q��9/o%�T=�`n�<|��?�k�vs�#)�TZc��Ki�S�'��w��v�e@�9��T%[�{�a ,(E��vL��V-���FN	9��L��F�c��	8�´9��CpUFI���_4+��=ᱩ��8��,��E�Y]��A%�.�X7��2\0����̱������t����8Q���ߝ������=J"�sG��a��rL��Bs��E���/��;at����<�l���x���Q/=���U��ǈ�b<�4��u6�̉���MA���1��8���N�Y�ʍ��������ڔ?�J?-9dv�1�3��̩��0]{i��=��V]���EU����cP�k_k-�!�G>�u�	M" b�X�N��kG��W��2� ��'MK3u3��8��C�%`Y�~���ٞ�$��%fYU�4�����T�ߖ������|�K�۪}BӾ��4��p������_��9�3L$'�8�|�Y ��e\�Kǉ�o�������/0��1��:����0T&t���Uz� �3>|�t�3D*{��.�~:�+Z�@˲�fRK�������i/��_͛[��9�l��͉4�qV���;Z��ճ. q�4}7�m�ؕV9Z0(�Y�U�Q3�V���U�JN
����pD�;k'ꦚ��89�c�n��c��tRts0����-
�ß�Y�G⚚�Ľ�y������KK�#xMJ�M��������H�똺�eƭ���w0��ay�4�u��(���6�r����\W�^2�w�_�����(<&�� �������uS�!l�b>���c#��29K���B�{�S^�tX��ԭ�"Z���K�U���h��0�ʗ���!H����{�Jc�A>�Xd�͑G���-i�P��̇���D�MG�ԑ�a#Jb�Fi��:�r�%`�)/N���ϯ�鸎��ߠ!>w�![��YGM�/X&�5�m`i��{�qw�K��jxY��x�+Ү��WDʇQ�\��;��``�֖[�Ԧ� ���T8��!�v����ɧ��ܧ��m��x�b3Fh�]e"'�[��u�ރ�,�>�.��AO� w�e�d�=+b�[�+�J1�#+Bbl�Nc١vi|���mG{�4y:/Q���$��6��B�����tӭZ���������	�������ѪrX�\�q:�)k��@�\9n(��s�!o�E�������|e!��ӧ����T�Hr�_�Q�k��징��j\F �=��|2����'eQv{Q�����WW;���O�RE	Ҡ����C
Y�����?p+�(}�D�G���)�g��}��w�X��tb*�E�}����̟N�Eh�(���=����4�.�d�c��~1D���/���e������w��]O��٩'-u�3t�0jy ,��gZbz'm�-�R4�m����tA8��I�r��}{��~�T˵Z{i�ĺ��ҫ��7f�#��������$}�L;˓V2��y @Q\҆���@�|�K�+��@l��M2(L����6��d�*�����=��O�@9GR�L��y�)��-�h�0XA�&x"F�-�{+������)�q8Iw}1P�S�'`�Ƽ��͌�a�t���Z*?R��V��8�}8P��nf��'�R`�\�rѫ��~�}�dX~�ޢ����^�Y�$�H��|�'���Rꬂ�h�vIr�����ۀ��f���T��0$�͸|6�Q�R8�YQKjf��T	���iAV�ҹ����F���4�L#����XɃwKΜ^.��+������X�7���_���W����*)��<E��@7�X�J:��.v8_?u%{�9�j!Թ��J�s�r�Td��w�������՘i&�+�,�}����)�;z��r���d�\��(��aQ�Q	����㓾`%��S4���d��gN�r��Nr}N�΀z�4�X�#TV{�Ǎ��h|�1C���h/d�(�f�kX���Հ#�n��Q�m�Վɸk&��<0�5�3�Q+�C�� ��
cK�:5���hv'��g����c�d@ q}�*�:�B7u�.pO���� ����p�f�3�K�
���0�lA��-�j�wVj4e��x l3l�����њ�[�"�kp�jb�̣J�+����0׸ ��+6A���uHC��XA���K���v����]-ϱڴ)��� ӏ��J�!��Oљ]ٱ~ⲕ��v�X:7���;E����5�!W@����� �ʛ�/ q�� ��A��`�o��
�\?��]7z_��uq䞹gǖ���Z1�\-X|wD�{�	5�y��� 0>�E�\;�>��������	��M<׭�]��j�R����A�{�V4���8�Ѩ��埦�p�xUG�-"� ��B.s��ѳ;+���2��,�
�U� n�os������ #�xo�zʩ��-c&2�J�!�ᩪ"�~j���fZ���kƈ<rY_~�6ƒ�I�7(EV��6�R)L�!8��4��u���!M����X���_Z�����I�2@�~�2�c^�7��L�ơhY���H>�U⊧"�b�Q��M����v�]�Ax?��8޺���jB I��
�Z�t����e�0i���e�f')qV��e�B�OZ�YH�o<�"4#����1^uI����K;��[ӱ��!H>�dY���{��wE���D��4�1��6o�MS�T6�joߑ?��p�G$�}ذ��<e˽ErO�6[ɸYt/���'=�"6�ϯ��+C+��{/-�����!6o� �p 6�8�!O��V�g�ٳY0_��
70PM�_�"�h���~\Uoo�X�K���d���� �;Yk`�����R�x����K�a����J[���u�.ԎΠ�Lt���8xEf������>[_@� 	�S���D��̖����v�ͤt	�|%�T}�r;V'�	�!%���$��+� Fd��Ҡ[`��q��j�c��k�!ݕ�� ���m��f���G�k,ռol��H�Ͷ������{�D��n�ة�ڞxoM#�Do�����ϱ�r��\�S�ޔ�����Z�n���k��~�����⸕Iz�ߘ�ݳ���;2*o�}��,�`�.B$ĺL�L'��lW��E)�ԇIBB��N����5�]��f��<�ڥ��R�^z�q�e�a�h������Zv&��_�Y�����xW�*�Zæ}�E'��&N��ǻ]@�G'K.��ÐQ~��<�kb�Mj*�?��@�x��蹔��.v���~U�1B�G����U	��V{>T�������VH�V*O:���Ìw�ɱ�,�p��D�\��uJx$�U���+��L��k���X>��R/���nsA��*��b|�,\��ǻ踬AP(
^�1N�>d�0f��V7���(j��UhXk�^R񆠋>J����Cı��%Fw����2���ۗ&��4�2�%njV̰���C?YaS��_�3s��2߳ ϒ73��=�Ey�)dƀ৬�X��P�`N|"K�S(��u��@g����i���b3�Xi��	}�������ͻ��ؤ���������҉P���rA�Ƅ���91�~Z{��*��OW�b ���ݪ�N�M!˧��Vz���v�<
���sl]���E@��X���ц�6`�ߐ�J�	���U��׃��f+����E��4��i�1c`3ٷ���ƥ��ǧo�s��|�&4by*��F���S'�$A��m,Q�!�D�Ur�9q�}|. (��f��Ч&�_��a�?�����A�/T��t������!p�������ʾji��f<&�wf��*d�~y��R���N��#c���'��У�e��@�H�x;�vBsR��G��\	�GL��V014�p���Q�a+��ƶ�ԡq���ZII6�ɉ 	�.S�%	�,+f�����C�S��%-���"B<�CE([~�N�����~T��������� �ޏ�Qr�f�t�ez�u�� e��C���@�$�,��R��J% ���A^���f�&w�C���=Y:��Я>���G�h1��� i�P���uo�`��<���!+8�Ԩ��t�4������w��Eʱd�"���$�`*����:�Fp�DXu�6�����,��<7A�KK�G|I�c��HN�!�{���'�t��kg�ƍ��Ӆ�)��6hG�Y7���)������Bh]��2y�V���ݰ���ʎ��o��d��J�UH��4���=ӜD�=S��K���s�(�e�ucK���{>��MȞՐ'��g*[����ȹ-�zNͺ$5�@:r���<f�'C�,�ۻ�#N�!�M˺�Z���ќ�_�H�ܘD/�c�����3�}6�ٝ��L���I+�O��r�+�����wʻ��Ȝ��߳�>Ӱ����%��V�g��oB"J�a,O$�N~b|���1Fp�IN�UtE�&��9�dR����ҭK敦��B�Xѿ�f)=o�%S���k�⸾2�A�19?��cTjO���O�9��f}��Qlu�ލ�)�Ek6%Y��+�8��?��f�!� ��6�1����-�B[ ��	�V�����^%���q F�~ܱ�C�`c���,�?� ���9����$nu�ܶ�{��U2��7bQ"q����~Acu4���f���P#��y�4;�v�ɥ_S{Z�1��s�t�.�`�
�<�?R�#�J�����I[�0�m%��
��|�=�����ެ�+��Ġ����{�`U�t�W��\n�&��h�V�+!Vv4�)'��;s�����l�gC�����b�iA���),w:{���8��"ay�Bur�g=H�`R̶��L�6H�$��ܒ�-�W4�u���%pK��ָd?���I=�⥰�^�ǉr�K=��?W�����|�]���V�E�o�0p��_3�U�i��x�3��e	�
�Y��D7$�g,����6���132$�m��F.ԩ;l�e�K�Uw�Ҏ���k�OeqF"U�s^���bmM�+^��X[��`f�E%&dݱMW2'J℄h:�Jdҟϛń��1n��yT���+�Ĵ��K/B��H�?R�g�KaS��&3��������\wv���H��L��:w�pls:r������������˒��9T_�mɰ���c�Gw�}ߢ�YwD�L`2�Y�j�D��x[�8�?HV�8�p$Y�"u:��
��L���T���8��_�,Z}0����-�e�ud�� �Al7�Ý1>t9�S�nT���J'n�C�;7}�^K&��$��� rnӼ�n�2��
�>�_��J�-�/�M�W��,��\$�5%��FJ�&�H\�����[�9���_%�����ă(�,��3\��E:�J����}�5|C�!���kFQ��ckews�O4coǛ�ʑ��C:��/������[
�/��fśl����/q���%\��i�Ƹ��ibf���d����!����j��`��.��8��	��p�������'Jd��c-D�bn8���t_�mw�	j��zV��&<8J�S���Ԕ��7�����w��f�im�FQ9��=���E gX���<;�ܴ�� �R̒y���祜(�;n�DŶ`�����0h��D��+�D=�������\4i��R�	��Rh�`2�2"쒇e0��x�ʩ��GOFDT���g���.�T
"��؞�I���>�D'���Ǻd�5<~\�P�&��j�SR�	R�&ۂ�ump����X��p1����`E`=��Ɛ��f�Ŵ�����~W��]ȦcY�6�N)Oc��jº���2��n��G�i�xa�qoL,�^�(�µ6�y��V-'�+��n7��J����4~V���� ���31�b{��Y)�"�q��SYq+���b�ƒ60��Up�^���֑��'��M|6�7S�,�d���l��=�y� ������,ľ�D�l���~x���
���_o}�19��9s�05��py�_<�9�)gB��4%S�$[��'	P�AwG�gK�Ř��@L8ZM����CG��gZHX�w֬��P�
�h���Ei��#��?������rɄ(��8��<h��2lDC�w�Ε8js�hH��c�]�?��;�Z�}5��6�8 ��t�[B���4m/��i��kG�d�,�l�4����4Ϻ�2b��F��I�լC@�q@m�ݰ�"&hme�a������I���M��n?Źi����7��us֌كcd3�R#kޘ2+B�}��Y�i�rЌy+�'`�;b�/5 G|�;�>c3��oYA�h�b���Hs*)Z~t���N�VMR����`7�����̤�� ���,�[(
�&u�2o�HW 8[{�O�)����?�q��̧�>p;�x��)���ǲ�KP�Ven&�:�v��"��Y(QCj�[>Y�i���.>	�zͦƂ��(P�?�Qu�{�Jċf��X`�(�燋�^���峮���ɹЅ����Ʌ����s��$�{n���0˿Xj$\zBް_��"f= 5�c�f
�)���^��#Ho��p���3�PV���͸��S���gw~5�tc��D0�_�}!2����a1N�M�����L����Pz˹�Ua��*��&�=>96����ߎ��M��#�w�N
�a�{_҂�h��F�f�Z��4������Qx�x�l�G	~��5��xc�L*�
Ґ͟9�c����\�dQ�p�!��$?���<U����}�B~�ЇǏHZ���:}R�x�2l#�VYc�F�|h��o���hnu�Kݲ��a̪SM7o�ǽ͟�u+���]��$��³6Ă�+^
����7�Jjj6��2#o,T��@Wx�1����'2�A�U�Dh�؄�����#�ޒ6ȝ��=u�^��$�Ak�*ջ�����v�%m�M[@��n/�a�M/N��m�:"C��㬼�3G.0NG�'r�cB�_�����b�*�@�"�Ե�zg,�����:k�8<��gZ��+�d�ч����0\���
d�>���$����n���Y�e=�?G}?Sj\�v�l��I�Z<VVs�W�`�}��E�&	��>��3jL�P�(�i4o!�K"gS6��`A�hWӆ˰�m�vH:Z�\v)B���^O`���Q��{�ֶ�'�>adq,������Ρ0� 9����B؊	;���L����vJ>��`�a�U�4�Xv���i!Ďƍd�3! *
��/U��)��q����lAՑ�{��Jj@ X��Ken�\רʠ�>[�I+C}����*�!D����X	���Z��^��@��K�ŋ�Q���˰1c�(a(Ii���Pgo ��5||�95*����2L�3'R����V ����Jb7����<d+�V��2�O�D=[�B�{��/E=�Bs2jX`;{��,m� �ܼ7T�n��O�,��`�W@7�R���>�HU����\�Z�V��E�]n����_!3ngN��|6Jޤu�&�Z�}2?_�Ҟ���,DV��?�ȶ�N�:�n2�!�D�56�ӓL{��ؠ�^����
����ܢj@�8�"�޶� ΁8B;x�ɼ�9�^�tB%�$���bb��=<m���S�g�w
N�c��ۯ�4R�Lْ�=�E���t����������ք�)n�*E�žW���{E]�<'nu���
��C=��*�M%�ԇh��0�`�Yv��x8�	Ez�c�NE~xcRaJ�*7e�)&��S�\1�C�����o�b �n��s��}��!�6з6���r�A7
=5mk�;���0�9�*�ߞ;vx�l�]:�Sd�,���h�ߛ�4d[|��w�G�{����(�d��N$��a�W�fgON7�K������#�t����s�c�,��/��L�+�lg״!ll?�gz�O���ZV8��X�<̍��7ʆ����n4�`��+#u�πUY��9�aLXO��(XU�N���0�=�n��eP[lj���״��`A�>2��k{��gW�rڑ�ѽ�¥�9�n�~|�o�wL���k��!UB�eqU�Ib�4�����/ĆW����!��<�ShKC���nȘdc��뭈b�#Ĳ
�>���U'�����N$�눟@ϱ�1�`M�x��Y�YI�&i;�8ƨ�z4e�M�vHj.38�!�+�^$� l�2��Ĩ,�C�9�#B�~7�Bŵ��Of?�&ð�h.mm�qk1�����)�I���G�ҍ�y�`x�v'gp����U��e�ͲӋ=�3���g�ZG�Å�@��)G�e_��r�fNI7�L�@����ə;]v��v�h�5�p2.�{���B7�� ������Y6����΅��89�'=d���a���cDJ�&=D�Z�rh�l�S��tr����a�vʱ�k6V��{�	_�X����PI$q�Q/@�FJEpuoB����=��/xF��<#YF��;6v箧3GiT�ɟ��P`�=R�&t�d8��#����o��w�-7]ǕNΖ6�ΰ+���#�����&��k�P~����ݑ�H!�d��K�mX�Z|�jN�WR������d���r���П<H�{��z�t�0��4@�$"��Z�;l�K
�FM�MJ����N���k��Q>����Y�"�ʈ}=�Mc��s����fpj�N��8�{��G�vJ���c��NR���n�]���]L:�6���H�S�L�#���>w��x����G�TW������e��;.6�u�)+�{ޜ~����ۇm@z���U����8󀙐�+���*?DF�Bb��n��4�eM��c�ݤ��s��:�`���U�Hq��2��Tb��K���՚z�van¹�&�c>��(�w��0�5�Wf��;�~�DJ����r��u�C��g]� *]<����u�\3V�Xk���� h��vڐ� {�MI��7AQ`V��zR�'N�c��ן�{,"�i3�O	���K��T�bF�&�G|����c�8Ⱥ��|P7�8�y��c��D�`��s�N�Ո!Ƕ/zS�ɋ��3<� �A���&�1��8x�{��c�އ�4���t�����i���@un�v�b���ɧ�a��Z��nW�=5S�3у42K�(=�����8�~�k+Z��,qk�:����QMƉ��G��uo� ���st�K��	kUD���¼��vSP����1<64��/h^��߳o�q���P��E$�}@�� ��)Sd��	Z_~[�����n���0������~�o�9ŉ9:�欄��>B����� a�t�s귾2(3YU%;o4�]2����;P啄���*���A���>7�MCU�ZHh�����v���q����w�M�3�����
�-�^հAV�l�{.�v
^ɵl�p3I�K�&4�}�~қ�N��q0"��ǖ�5����{��?�a_�׹f�� 8��D���~�6z�Q�D/2�������YOi.s��� f���u�_MyW^`�Í9^�A(hܛӹ��vx0����?Ϛ9)X_�0_���-M(�3�>,�c��=�R*Qi�O�>�@ny��/��)��+i4��ǫ��Gno�ͬIv���-��n���,�8�S%�c�h#S6#�����\J�)I�3mFHP�N�{O�d���'��|��џɺ�/Y�4ֻ�E�=[k��[xƘ��WA�W]�#�j4�I �Tb�w����\-���������%\s���%\�"����u"J{QƋ�?v�o��?�*(pqr=;�9^�T����HWM�){x�Y�7��,o�^Ū,S�wh<%ol�w0d�薌��~�.y�ƥ�K�O������q4�d&#�j7�͡�8�'Te�I OqO�������$� �U:1DǸ�Ԥ
�l��{v����Q-��@�j� R�珤�G���Y���>��f
X�6zb1�k)�@P=$�U��4EF@]�٢0�O~0�0]���� ��`s
"��$�M��M'�P��T#K�7��4.|b���?;�"p�gD$r�|�Wa�"\�S�J��\{t!Ρ�tk6k;��O��F\��􈿃�i�n�s��:������.MZDa�M�]V��r�����v���c3򺌭�U �p͍J���k��I��׍_"�+w���b�!�i���q����~~�u]2�W�е�f);���V���5���'�;tz�䝒Du*/qIE��X�:�d ���V-hRB}\R�Ov`���5���K�Ċ���c�F��v����E�.�p
����r�BkW*��GJ�GB#�>��~5��qI�Lc����	M�jI�.�O�e޹�[K�������	�E�o2P��d�4�<O�uj�4ܴٸ��k5���/p#��O/EMÙ�kM����(�w!��񶋱
2E�ˑ��h�׎ֿ�B�f��p�G�N:�|�?���~�k?C<��k-�M��H�	�V��^������GJ)_~��:-�#�ʭ,�깒�e��)t�cϫ���,�=OL�V��1�����	��� ��뒓餐A�Ven,kK��Vm���� "#[�fsv��LB����U����2��`?���֝%�S�
{#F��I-�m誣�P�'Y�h}V�&E��=�)F���.oºb�|{�����x}aZ*�A�֟�H�_�h�p�1��C�[p�G�K6J��5{{'3荋����={k\�Ș\IF�v��A��[.9߭2N,�]Uʉ]'?c�����������U�Z�#T��Cc~exmx�r�x��EE�G��1�Vڴg+�Ƴ��n=bo{X�����Iր2��{T�����{L�|q-�菁2$|D�ۭЛG�浉;	݀�A��iɎ�N\X�)a+#�R?��@Vn*Y��B�F�M�]�����p����,�&=D�^���n�V�?��޽�����b<"����e���;-C4:Q��l4#�8W�w��[�Nil�_s�o��3L��(!؏�qFt��<���N� ��.<K��&����y�P����g+R��S��7��h���M���ڮe��3n�ѫ; ���y��}L�(��[����3I�*���f4���x��]�Dl��[b�@m���^rgn�66����.��J=����uQ�UtH���٘��)���?9g����̹���V�*v/)���^I���p���W�ŃI�Ùon�xfL[9�p�Y�B�D
��
�9�5�3"��
�q)%�t�����б�@u�G�C��yi"V�X��� �h�[޽�W<�S�Cl��֎fo��f�,����!u;�Q+�#q�H��Ss;��
�5h�)��r��Q���Ձ`�E�Yfyts�-C�'.��kʜ b��b��In��ց���)R؎f�f(X0����v���f�����>^ɖ_������鍷�B	*WhnZ̋9� @k�&cF���|�~�l�<�"�Ή�s���r{j�������MĲ��T�s��m���ߑ�[a�"UbX���7�Og�z��s"jb Y:6Ɏ�bm��4M�j�)+҇�d���m�n�wTc���3�֍��c��]h��e�D]z��vN=�z<�i�����.�_M� ��P��I�� ءh!|�]Gu�Oȶn��#�}&�N�]+���wk��q��SR�&ϣA.���($�a�s�"�(��VJó������!v��*�:%�+��&ʍ�?,#�F���m��-A^���B��zR�-R����n`���_͊�-�{�	�4�n�����j%ؙ���T<w�Jο�@m�A��d��^���8c1Vat6n�is�5-�p@n/|�{'e�q �X���E�鋱��h,�i�S��(Lڱ��t�)^xl�I�܁���ؾ[0'_>d~�
d4��u6 �}��&�ZJv10��<�E�R j�-��E��D^	� F��ǃH"q[�0?���9�5&�9c��rv�(8��	U���ac���؎O�FCG��ɫq߁�[A�f�ؑ�|��3��Q=A�,[�)��_I/�N,�5^�C�*_���~�����O��Pl��4�$��	`��N����OQ��ϟ�B�׭���+��\��8�G�q�:�A�;b�,���-r���������gb�}�����ɪj�G.V���a��w��d���Y�^���=d�����uF,����5��톎�F���6c�`��X�� ��lFˠ�������τ0D��dt��\>T���?��WA�j��/�w��W�����x��m&�&�RE���^��U��]�^�;���-���vu:'ZJ%7�������Vm_��w�5�e��8�����bI!V��Z��p���E������~�������s��GDʪ�zS~D��%'>��y�-[E�@��ȆZ#o(�>/�ɖf���'�ޤ&�D�\\�"�odK�bm����Ӱ�=<?!1p�SPKrћ���É.��̳���X�-*j��z��`�p���&�4�z�9��8�t[[��_U��_��俨�@��p�-�L���!!�1��
ɍ1+y��F����.�E/�K�&!�O��Q�!/|�^��WJs\��Ny)���'�i���%e�^^�<�@y��V��E����`�PhylLٿ���΍U����h��]�r��d�S�[��yO�@6m܀���1��6 ���z�l�ߑ�T�g�m�����v���Hn��(}� +k�J'
��xAĎ�<
)#�Z�7�y�«��Yħ���65������Ӽ��,�Ȍ�����0��A`�e���m�����-�M�e��Ak����&W��l���,�@s*� q]ئ�5���"N���+U���>? ]���9�9�UK.@g�����2��-��=��~'n�-��R4��ċ�r||',އ Z������a������v ����y�'�����7�?HH�F���o',�x\hoTo(�CѺ	č܆M�������i&��z���؜�p�E���UuOԊᒳ��0ުu��S�#�u5�`{j���! d�MƗO����f�P�;��5�6ԗbU&+�[~m[����< .]
P�Х(�v#Hծ���&6�a��w���k���˕�����UYރ�Kӽa���خ7��좋+d7N�����1���ѷf8>��ҭ6~ɋ�pfZ��r�nhb�z���%��8�A��U'M���H悵/�_ٱo�h����,#���+$�b��z���Sm������}̰�������Pk�k)�yI`�i��ܦ/����UW�o�$�����f�� �2u�kb��7A�9�&�l��J7�%d�U�	x������Z��y�=;1¨D������٣˺�¬� �m�7��Η�6b����������F���S�R!�b�X"�w7�\���蠕���#yI*C�H��g:���%�=��Z>�{��l
�\�D�?����L[^a}yr$