��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ�V�P����W^�o��K
͵h�����h�
�;� X����x�Ep�*���'�p˂#gD�4H��fZ��"4��V��6��cq�`�7խ�:����%�	��H��\	516�K�W��K�����T�Ԋ�MBUTA%������Gނ�E�)���!Be�N���3�ti����'-&�y�QIG�ϯ����mSwOb�2�a����9�h��t���Q�u��U�m���J�=,���4��{?��Z��%w��0M}�6�X�CP��O��E@�j�M�ؑ;���+�$t�eS�xc�I��06�F�n.�!����h������
��~پ@���eps���4fL�G�F�9��dF{�p��4�^��Q��'xI�x8���\���#sG�0�ǉL�Pʻ���2В����r+w����U�n��V�)�O��x�g��{qj7�ݼ�t�9�
��l�����a���,�[�;_�����z!�B<i��gλ�吙֓��u���V��
w{��<]24��Qp��ce�(�ЧrK&`�8����#���$ǏV6�m���҅�32��lZ����߷����G� m�q�NF ��f�V���M�<�/0�����9ո� �E�E�يF�ד�o�&��T��V~�HQ��9="YU5��H���bV��sǊ����1���W8�ĸ�Җ�R�|���ȇm[��(���q��Tb�8o�w�7�e�� N��\^�7v0B����K^��Y]��M
�"�sd;��x.	3�n|&#��>D@�_���t�zJf(������.n����a��>������z��?ޑנ����g0�w�a�d(`���� Y�b��zJR8�O�Da�}!�u�D���/�0Ԛ^��L��Iz��ҡM%T�0O�G@����R�g|?NN\3G��Li��h�'������条�ձ sc���`�I���^z&���!�w�io�w���53h%�7qKy�cK�3�=�8�]&��
��:`�8��(�G����&���汗�K3ǱE_ 	6"�(S�CQ��Z�,�A�%O/s��R%(��c�6�����p�ߡ��;^�_�@��S���Y��&rS3#e��$��\�^�U�7���+/�먒?YxA�#����i�eӥ"�Ê�-*�`u��nd&�8�=����l,G�fN0�����u�����Q�83���b�m* �}��<�r
���^iS� g�()�� g}����߃��<(D�S�g�%��1�o�M�l���A�" 	>�A���K3?���QpŴ����]�8��q�i�L� ���"V\��
%M|����J��	;y����N�ѱ�o׫ �l1�]Cvk�[�:h�0We�4�4ںNd�
B��ܨ�	g8V���� ����c��I�� �@%�X&��(�±�\�26�Oc6�.�}�M58w7j��.v�cn,c�Z
�_߭j� U�F��ciFz??!y���H�"�H/��-����}S�U ���Ma�w��_,4KA\O��4^V��c)����m�xG��ڗ-{6f�P4n/S[��
��C�D�,��Dw�jG!��9�x��6昽N�Ck��BG>^;��J��~���Á���|A;�2@Be��0g�|��l�u6�D9�O�f�aV��4$0��@U�+��/Q?�2��~�){��?�/kg���%W�{��%G_�S� Fv�7�4�;&�L���9�����-}��&w^!���a>}�ޚ9�>&߃��X�8^c�c��_���"s���V�� p�k�L�c�F������Z�_pԶTf�f�뛷�kL�#��8Ǹ�OБ�hi�������:�l��ݦ�]�S�);fC�`�e��Z�EP�������� �x�7~��I�.�`�Pxo2/ESY6'���<C�}Q-�v|UU8
=Ț�Rm{������H��3�[���)�'�w;7ReD���K3�v~��.�U`�!ӳ�"ݗDx���06��}�A���ڂ�Tٓ����e1�w�˕̹�;�Z��>he�ԫ� Pi���vap�󐲦���l�x�׎s���i<��F��Ӷ�������U?�m��3�D97Bܔy����S9����c�i�Cλ�趁z��5a/�`m?� ��>�G��SC "�s�[a��_ĜJ%��M��U�V7e;CP���ixU��H�i�� ���@���Gc�	DL��Y��2�	`w7N����f��5��C����\!贼�O̞�+RZ%=�k��W!��KC���w�q#�)���.�;#�D������=_Y�A�Gu��ky>yh?��'=�5Y�ۓ���g/2��M3Z9��jEQ��ǩ�"dQ�ܻr>?$��E��?�K��^9ȹ���/>y�%��mKC�����m�p�P�zP�O�]�[����<�>�$��7�V�Z���t>��.�� Ҧ�1�����"c�-�J/dY����g@SR�F#�������{��}�)�1g�S��1o���V0r>,��@7��K3߄QH�f��6b�s��&,2��@G�Byj�xita��\��q�����;�X�"�&��<�T��'D�Q����J2�BQ����82ZI�~�D{��Z�y�w~���6����@֩��B1oK�����ȞG�FH9����)�ې���vF�$�O�l����"P��o��y�=�/�82�	�h9�J�����{��2=bC[�n{�k�9�	I$���b�"���o���ɂ���G�=���E���mB!}U�NV?3����0Y
�����b������(S��ѹ�H��82W�#��V�[�����Ȍd�XHsX]!Ujj��9}�ĸ.#�>��3�d�iU�J��A&�Q��һ��u!k�a�ug%.���4�%{,��n}�N�S
.�k�|x�,�}	x�����q�p��(� ���)�W�2�z]6��}���rJX
�����g�s�i�L�H֧����I�X�`�%��jW�k>)��9o0jsP�* /]�Y`7`�V�H�4[�FF�/���$h����Zo�9�<��}N�V0J�b���v�v�����ߤЄ:���uH���ʩ��;�0Һ�ÏUo�עb�uM��]#����g����=�8�:���a[H�/�Q/#�����
d��>{e���bxa���>ԫ���"��*>��c/m�l�F8��1Ң��B\��i��$"X
}D�\7����Π�q��R�*7��9�*	2v���N�h��Z% ��r喉���Iꖿ/�"�NU���
5�ɖ-
��w,*x��E���,uf���B�LY���K��z�6�²m�Ż�M�AM;��;
��5>R
���|�j��cdꠊ��	V9x���㪢;@z��7��f�f(E>���U4/���E�+��"��{\pr�)��k��g�,FB�������� rR9��(�?@�9<�7�qw'g���/v�i T9vZ&2H]5Q��#�h��23"r��#����i��Y�m��ԬǖS�lq��sD��fb��#r�ض�%�g�� K��o�o��K޺FD��_���ԑI�c�t]cv^tHTU�����l��[ھ���O�ԧK�,�e��痯$�~�Ul=��6�柃RC�_*���ɾ�����myi�!�1<�1et^v7��,,��Q�:�Ϭ�}b��v�1	ًĻp���p��;�LB�'�D�v�n�VVu�=%Ͷ��6P!�Xq�_�z�7P^y������RX=���Y�?���Y�n�G��.az��@spVx�ٓ���d:��t�n"{��������j3�<u�u�us���L�|�n�Q:�[�zʬjiK��i��BPfa�3�?�w�u� ����� &?@�V�R�}�FЀ"b�����K��p"��Y��	ޚ�n�M��'���e�E�@������mo�a�!�E��:H�6*�� �fh���;_�[(�i��K_7m����4y���.9=�j��%C	!����\Y�
k|�ә�f򍌻�����'��B����kH���O..����:�J���|�J���I��{�%k��T_���	)���s�5���.�~�"��:�v8L�ݏƈ�s=���	I��8gRt/�) ڈ�S]��q�t��tY�|�Ԣ'PLf��έ�w�U?�2)���{R^Bۭ �\%����e�Ѐ�8�Vw�����Av*���M��7b{�6����RMV��.�f ����y�d������W��&�PT����iҎJ�+�+8� ��&d���(�l47Ôȍ%��Ay[^L#���w�<igi�46� LLދA.^Ϸ �z��H�q'�N��� �Zq.�p0���J�`x ���@�D#�jܼ_g/�,�T���ո����f�ka��k�=R��M�� �d�J�l#/u=�376�ɲ���%�T$Rv��t�u�
�b�6�Q�?���Sa��Ṑ�sŽT@�X�O���WJ5�OV��T#���L�~�Ҋ]#B�x[e�)��n1K�0�z�.�T�/�7Ad��i&Q��!�y�d���nc��"�k^�����W�>� ��͐/^J�u�gi&KHjz�]$����g\�uTO׎�5K7$3n��j	�)9+��$��7����p��a�e��}t�m����b���Θ�t�	��5�L��\���u�ג%�`T� V<+y��'#P;��h�ڢ�0����T���qN��sFé������+P(+䠨�@�}��"��ܐ�����O���[���5�f[����ebq�?�����$��ƚd��<ƌ�����exF�br��E��SKX��Gؠ�R���?��え��Z��$y�|���13�2O�R�s��U�#5E�w���v-G�&=�g�I
V2N�	A�0ǲ�v@
�KzwRבP�����S��ݰj���u��o���]���<�N�h��Go8�jܯrڈ�@)��2ߠ�N��Y$	R� x�
�B=3ӽ~]��nN�u1ޗM�l��c#��C���?;�u�Uͷ�n��ѭ;�ܫ�홱
後J���Qp�ϔ�[���/�d^E�*���}�	�Y�;V��1����x�_](�6�d�qQ|Fr(] �a���~��Ҕ8-�]�6�&F��L���G�a�A�����֍EA�sp�Z���]0�$�f��zڍ��mi��Ue�UK��7i&���UT�C���Ȯ_��	Gt,7(	P���y�٣m�����<�6�],����܉t�z,+��Ł�	�>d6��v���|��~|�~v�-S��n9�/u��u��e�t·f�>$ŋ�*�T�q��i��jW�d���`8�<�i��x����9���1���f��E����%�AG�t<�Q���tB�|+���yi�͇X�i��~��r@�|OŏV ;@Y�y�U�i�p����"B����r�(<��C����d�D���{䮓J��-��\��ߨ����ȸ�V����2�Ԁ���(�bɃ�fK�o~\�#�����T�~�Y]�
 Qn�&�^��Oo�Ue->AIT�����ҰW?<?��鬠M_�4Qq��f��(濑��''��|��Ld����:��vI8W�H#e�ܬ�\��(�i;�Z��z ��k�X�1���,_T�����3$uxҔ���+��ة�!Q	a�Y�ʷ�͡j�>�T�;w2#JC:�\x?%L��?�`s���|vIzh>�&���`#��q�?۾!�O��i{𤀃5�uPd�}����ޟC�m/�<ºE�_�<$B��t��k�
w.I��y��4�:|�=j�mi�@T��X�Ĵ���r��}ad[x<!�f����"����t��|���;tL�j�C�O�M�`?g���a���<gL>�l"�Ԁa�L��(_�j��W�_S�@��9r�eC[��	��j����sd�Y�]75hϤ(S
�mk�Ao��v�(�%W(W������<}+:tV4ގ\"�V�ˮ���#��3�Y�����2l��� �%i��Kw��mq�+̓(�:W�AP��L	c��m�H RD��0%�Y��ܶ�͓7e~�$��u?S����Er�[�X�a4>�LmC�[k`���1�׼&���w�3p
@.G���1�����ї�� �
�Y�<�~��I����h��yd�!B��K趴T�m}TTz����a����86�)k*}ƧQ����v&6�\�虯 DE�ʞ휛���Ȁw�����w_�����J�rʬ�X��w��=���ѤgEq	��	5\l]7��(G2�IJ��
���|#�8�E�=R��W�Sv��ܣ�B�Y% M��E�ͱp��k �v+�P-ی�y:mmK�q"�?M�@��Lh�7�O�gD�nl߆�]�zX��
�jS��#ڇл��'�}��Ks½��.eE��q�S�w{N�����qDc��V�8V��Y<�op�#�.�?�,.�_3'U*��,�m�\]I �����$Tw4����sV@�m�t��˜���̌����_�+�%�G�MԔ�A�Z�ޙ�Bp�v����=e �Ѳ�?�@$�Y�V�L�82���7h�}`7q3����N�f�Q�,~ޑn(��K��q�Acv��[v=��Sj��?��GiRQޖf��6Z `���ڑ(���ʢb��X�e��:Qw3�4��mw*�G��>�K��0ɇ��a���@g���g(�X#6�iۨ��!j]+�>R����,����(0u�&�ٱk���Y����%^s@���	gN){�2A��X�Y��K��G��� ���,�-���x:��X6�o���.I��s���b`b��QvM�b�iX�,�/b�F5��!�@��^���]D�����O]�;G��\�s��G�~O&i��f
e���ي_&��-]?�U������i��['sv���|�j���%��óx]�ӫ��kG�遍���7&T���Rҟ���H�`xw���C�=��ș�t�MJ�uza��' �ߓ�P��,+�L�.�o�IO�^�Rچ�*$�b�"_���C+OS��/%���`
����'��[���1͝B˓�ԝpT��W�����0�1��6Q����ӹ��w�7���|Gz�N�����u� ~�dA��#��MU�8.�x%��z���߰
��v�Tl���A��`?'��.�t�Z��m��"Vm���b-����L��J��Rar�����|dZ�FAC���̡�nfݩ�Ls�c�>T$4=',zT��p7&��ϻ�MC�_��p_�Xg0㽋=|����J
z�|6���Rƀ� f�o����_:M ���;.;��xJS�"�G�����1	�b�,�/P������K��PM??خd(�9)�<���[����S!�޿V�.�D���5�)O�b"���G�G10�;��5� �`lĲQ���l�ȼ��x;�IQx�d:�#Zf�c���� ~��̤��w���?,����d�]�1����&�dz����wYx��l��׌��|�Tt� *���+�@BT~lw6q�E��(Y<�	*kX�d]��Z��t�����\/��8��`%�n���ra�= 4��@�\�$e�كg��mqU��D��p�����O�7�*������ ���R6��A�8���oBiCD�MTJc��Q��Da�����l$�Bn��>�����=�-�]E7�Z�6���Ԗ�J)=����g+��jPS|K'���ɣ����1~0�[��FZ�S\C�[R�և|v����E2ߣ(�_n�"�M�42�]��4z�C�r0��aMbx �$?��A	J������� ���(��/1�P_�R�u��,a3y�-h�ױ�}�@�:�I�n�7�7�LXb�	���q5��j҉#
�_W�d�}H�a�Y���i܂Z�}��r�3�Mt���y��U�I$���<�x ^��eG6���f���v��,����S�5U>=D�ԘV�/Q�)����=N�#0Ad␙�5�m%�?詉\��k��u�Q*����U]��#yK�F�o�@lA��|ȶR?N�0lIv#�b�}�$��}��R��Z+b�g$%�����H��a�BE��;w�Tލ�W��F}��p1l��x!���̈́�bD���?��b��B�ߩ>-'zO��jlᒖ���Vzq���P渆�JyE�����7����cl�m4����E��˅��9w5�V�$}�O��.nEF�]N���꛿<�~�\�&m�Q�)f���,l��ȫK��6�u���!��dތ��ŪE�u%}pa�E�'���jih`I�8��giX!��R��]ʇ�0�&��Y�]-� ��ptX"*�.��e�4�JY����s�=�j͖@˸RTC)�4K��}{+A$���[e�x�i�\�0t���!t��]��N�����J\fk:��vRe�Pg �a�8�{�d���%�W��1�~�0BU'����x�?%Pǒ߯/&�j�K0P׻���]9gV¢o���H�]Q**̈7���$�ܟ�3�E�+����EL�tT�H�<8!6��/����7e�V$�,�p#B��2Km�7�]��8��%K����C�SI����Ҽ-��|]��qK���L@�:Y��;��+>�št��^��2" h���KD����4�X\��W^R�J���M�	s��7B����K�#�+6���q���ٝ�0c�M���Nf�r��
��mW�� {�>i�Ђ��~,���So<Y��@L	�	��N�����x�!���,h�.��@��t�1t������/�R/8]"�h!nŹ����&|1$����/�e�|�����4�l�}�,�ri^���fG �����7`�egn	ʽ4�	�T�"�m�u$��������v�Ύΐ��[4�"�Ȅ�N5�_H��蘤���W�uB�T�T� k1ׂ����}����9%ߦ�1F��X�-��Β>��?��<�����h|���@�D��:�4�6����Z�<�`T���A��51Ap��%1�O?`{�3�*f��4�5�����BK��^�g���I��o�z��H���Y�3��C�l�*���z�
�y��A��������d!�tj!e��O�� �0����ֹoG���boʉZ4�S���~�=?)Y�֜��֫�e�W���6��C�60�х�-E��K+egy�B�����8*Y 5}z�\�*��Ķ��3�ǽ�w���'�&d������S�#�y�*&������jF/*Xo�.A���GҶ����<r�|H��v8��Z^" �p9�T{�J���TN�L��w�m0�l,��*�˴���������t8��@~��G�J�S^���M[�f�-��`^�z�[�7�c��T�e{!Ɂ�y�auK�Dʊu�����(��v��*Yzޜ�s��
�b2h�j<�I���C�&�{��p4=L�;R�����Oۆ2tJ�K���L�Na3V_h�P��j�L���yk�[�|�A��Kv�n���������nU���o�[26s�
�[��^��U�����C(�QQ})i�r9>����Lj:��T��^b�J�N5�%[{�^��k�;�Vggr���^.��}�$c;��L�2�ջ�*�F$�1�
D��l�+�是����0���8jM_5�'���-��:�TKS}|�<��/4WA�Mx��gԷ���q�
��K��m�ࡊT,q�蘊�;��b䜈۬����M V�ˑ�Z`��{<T)���~ѳ���cvv�²�+��	8��a�я�+�׵�N�����!�%J����	Œ܇���a���J��%P)׻��^��폈a�d��P0@���J(��7#t�ډ��m�!���Td(�Q1T1�~�������(D���9�v���։�;�l&��d�'ɾ�~0��|�ʓ�
��O:/;�q�U2YwU��p��;ֶ+����8׫m�k8�@�dAT�RR���"�vc���A/p<�Þ�1��)���?N�5�_�TX�����(@�"�	�����A�~�wOo��Z���,.��""��ֈ0���w�'lT��h8^M�)	i�y������*��\�
��s�$"Y��G/����?��N� +f'���	����h� d}j����B�`YN�L>�2���ݩ�D���U� �wW�s!��7`өp��3
��.)��hRz��.W��)W�!I#���~E����Ҳ&�=�����j�H�X���j��햤A xU�
_`��
ಒ�q2%��+��9�|U��)������VX.w8.�Vm�GқM%\ n��=N�M�iDg�n��{���Ky�=V��Q�EÙ��"U��T���Ф`��|'M���E�^:��2��!�b�3�s�3�W�SV�rv&�����)͙�A#��&S����|��]��hր���� MOM���Cc_{�V� Hϭ�nT�d��t�e��������ځ�H�#̅jl�����Q�f9��@�ܕɟ������e#GM%%Cud�#�X�c�`�.��`o��|�Ol�$�1j�a]Fn�W��6�<,��U��#m��݁/oѤ@֝Xka��m\eZzĉ��h�/=vi8�G�`;�0(�C!�>FY�3�(Z$��
�uT+���?������s^h�:U�7�P���b���� �kٛ�t���6����̱N:ƌ�б�I�h/��T�n�wϳ��.�^�k<c�)$P_�s�L;5Q �� �#�s�A�_��߻���B3#�V��=q�	��������wu�d*�:�/�+�9��A��R+���w���w虬�Q͔{�1�Q�F��9$:�G��՛c�o��[��u�;u���e�3����lV��l~#a���=s�<��� �w׸�Ԛ]"@�/�a�웘~���+����v�ӷ�F\s+��C����t��)�?x�LR�mwߠ�l����zc��ʷ��0d�{�~��9bxx�E?�����;�5 ��E����7ֽN'����5%n��LI�ϼ]��L�u%