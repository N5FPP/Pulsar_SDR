��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�۫k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A'xin�XO�v⨺��sZA�R4��g�psXdm"�d��Q� N���Ǆ,{�]򢖮��@[P{d?A�lc�R��kH�̈K1�������9G�b%��}���>��vC�).A>l�<b��������� �U3Ӷ�����n?&�ON��<��sC�d��һI�3rs�4��$�I��пԨ�
�v�=�`�QXp�?}.щ/�'��z�F�O.Sh���;�����Ţ4��虲������oS��7Cz�4dyu>�ڑƘ�Hdd]GU���a1�ۚM�ګ���{I�]b�x�j�-�����Kc}w��z��\�MW�v� �&1M����a��m���f�v\�2)���dQ��U�"��Jܬ�Խx��6�nc����
��]�r�	TT��|��kq�3��
���*ų���o�Pz2����+C���s r�p��h�k���:�.>@�����q���%�K��>����5Z���R���x�j='��G � �o�2i�=3z�vú�nE$��t�e������h�d�J����v%�O�r`k�����t��P���0�x5go�J=�fq<{�wY��U�����4�nF�S���O#��z^��Th�'�O����m�Aג�SZEjC�G�Z���x9�L�Z���`�0�Ia�w�� <��*�W�C'�`d�񥤤��c�S3 [=W55L�� [{�e�U!'=�;�!s�X�W^��j�4s
p/on�j�V裁T>*�?�G;5�,تAh�<�m+2ϏY�����~��r�+�Lv��F����Zj���(T9'Q�a9��qJ�+xazT��	+�I�N�=���ch��.��EL�>��%��H>1��JI�Ĝ(�{�,��# ������2�h6�nL��@-X�oz�ϑN�S�6���~�.݋Vi�����G4�B2�m��P 0}�4���Crl4�Q�ۅk&jTg@�
�ҍ��;Zb��a��x�+�4�.�?9��#*ۂe��C ��b3�&�����vTEk��g��l\yf�؛(#����!p�T&i���-�Wa�W'�ս �k@0��3�n�������D�X��0��r��p4�4�̊��E����Y�}��1��N���L�£z���
S�������\�����C��tgZ��O�f�V�E�n���������Tyh�-��iﮦm��;F�^���^���d��/�O���a�-(������0����J.J�͝��n���7�n�1���X���b��n��o��<T�A1��q:��A�8�|ѧ�jL5@�5���/�6�GZ�8/���_J�!�s���%#�J-J>�~An�������t�w��VzE�N	�"q4cr��Mg���i7;e#��6�I�Q�F�w�P|
2M~���TAQ��pCC�&��:���t��K�^nP;�;�X�ՐՀA��p��_����R�I�R5�e֧��se~���x�/,���۾���!�{�J#�~�S��/�����L� ;M�$�]Yt;�03C��Jk��0	)�\������������kpijV���XEm���3��nN�@�ܕ�.}ǖ��Q�	B��|	�G|