��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>�m��`K���?�]^�6�,X�B� ��dt��\�<�bT�AT���*4�M�!�c@U�v��:B®�H����u����w&��*R��Q���\���h�NC[~��p��/���']ܑ��<u�˜�Hy�����#�������D��*K�x�����N���^d�Y�iZ;���p�g���&m�däB���1j����Ơ)ק�Yto�{9��{Y? �Of�P�1�;��g
��`T�Y=�����5�و�-Pa�c,���n)���##�r�����a�9d���S�M��mOFZUUD4��C�@�Q�q�Q7�Lxy�{����J;8�wq��yI`��m����LR�6���%��UB�e�&vY�t_�l>�{��p�wj�S��0���vMTk�t^T��"��ޒs�d.�1p-yk[����3�۬�A$^ ��&A��<`��!�#ܞ;�`�>1�(�L,���	L��D�"����#R65O͜=R�i�5��/��[t"�jZ��}�g~ �q��a.��o��.�"�1�O3Do���g�=&o���G��X�q�Sq!���}	��G��r�H�	���6��nPo��^��d��g�,�e�,&zv�FQN*��E	XҰ��gY�9rk`����\S�@���]`�mܺ�I-Ti��=`֒�Y�re��N�j&���g ��zh�����Ej�e]:c���r�9i�~�~Ѩ�Xb�La?���Ԍ[�ZF��:�����c* P�
]h�'��q|�	G��-��x�:��!��432����c�3n1r�5�rs8�\���$r�p��7p�+���ٰ��T����b��g���k_B=��Y�c�}N�ѕu�4�Ra�O}���vH��>s�m7�H��N��l�}Z��ȬOuk�Jҵ'~S7ڏzn)޹QQ9�Y��%g�~����,����Qwp8B���� �C��I������_�/)� �z������R3���)��7$X�@�z�KX�?��+y:;HG{��xZ�C�����NZ���@�~�+PY����ޞD4���]�3��,-��X�����?�(��eЗ/�X7�w�oߞ��T
\�Ef!�X��]q����t��.�c���8�X�þ��.�:�5f���{ܣ����O16����F�w=-�����U��jA�*Y�L#�]I����K��D�7�;�����*�l��7��ֶt����
�D������.� 9�K���SCs�.L���_(�腕�k�d�|���`�$�UT�M�KR��K���+~����4�\i�)�:��G��aؤ�`����X�����s���_9%Y]�2fAd���,�[�Mz������r�mU[��w���_��!��|zx2�Yw�5:���6&������8��{MD�"�$��[?���|��=�O�����q���N�c���	F=���.�k��1#w������=2���i�,$���A���%�����?8%�cs!'���i�����x�$8�j�(E�-u��(��uV=f�{�l�OX��
�.XL]�� ��U�P'������3��i�'��n��u+��A�#�q[jK��dݼe�A��'�S�4�N��D�ޢ�2��>��tlr����D�ם/"�J�e���k@��/_*Zh��9�\���V�LU�cd�����λ��Z��7!0�V���3[�ݨڠL׼=_JC���}3�UYËIn;�<���h>�Skw�ĔX�	��[�L��_��#��A�����I���b�ɦ��\���E+!��{5'�gjM������)IF����V�)��C.�똰�Q�[��c��h<��Ґ���h�T�2�{2����=?�jd�M0�7qg�A��sV?K�>F9?�Q�FNamJ��B�̒~K��:���o�*�Ӳ�}�P��05]�ј�N�)���$�c��g�H�x[<HL��֗P���}��M������p�>�3�gW�4�seV��F��^=̢�dKox�=�:!!.*�vw���P�p��Z��>#�L.E��םv�O՗<�}��1�0ZQ'��7�
�i���Ph��n�=̾�`��<�t�Km�+`�'�ق�����-����R���I<�陓'+�j������`�@���t��r�,������I<�" 	���K�t5@��(�>oC�wr� �xF�����>pe��:9��nr*�f���-�������d�^�0�Nᜢ�Y��[R,��&`��>w��r�㾋2�o˔
	��=��g�6���Ö:g�3w�D5�̶�`�D�5R*c�{������n��t�͠f�߼c\%l�l�	z�aŁ.�Đ�]Fde%	���1ڭh����G�ᾯqh:r�9^�t+��J�ƅ�#d�eJ
hԻ�<_�W�5ʫ4��\LZo��2B���+���}]��n�}$?v�Le�[�
��|8��//�č�����䔪^��XC1�]�&�x|̽p�gx�O�GA�0�5�3(!;�_7�5����*ފ�y��c��9d6�J���eyj�~,>�H����ĸ�p�;K]3Q��ѫ$�7�۽}�B��'���핔Y�i pH�~����C�+y͐���i�%�U�)��S\h��[/�m2�-�w�$ ��It/ yK,�5�T1h��$]�ʖ�N�z���hV��#���@�6��nt��:RP������Ok�B�1K/�m(��.HCd֤;_'�;�.�T_�ܑ߯�����Y�4/�Q���@�5?�{� �~n��?�n�����x���Gzѣ)�FO#����Y�ʹ>?�:~+A����#ޱ]ޙ�8k�t��ɳ���3� �(��`]��o���"�#{��4�`?�0i��;��f�8�aC�����'�h�[� P��.յb"[�J��3�'�`)�'y̿ܲ����`mt�(�	�g��ϩn=:�*L:�r��
t�9�)������7���>��T�T+� �"u���©h��u��g�Y�����ǎ� 1=zP���}�H>�o����j�#<L��.�3�z��m��p�~��Q2�Q�N�O%����<��fޖ�lГ��4e�z�e/װ
�6m��$�n�-w��P�2�ے	Z1' ��$��D�xy��h��A���`���2�F��T>!?V��[�P�?�ದ� ��М�,\i�4?��W�m_V�Eƿ�I~�H����K�#��B0�����L���ӑ�4���s���6����Z�(��rU4pJF.ٖ��]CQ	�h����.rgԈ�6��?l�5z��T�����/��-@����^x�p{3�3}�o-ZYکF�����2 �JrF}��c��|B�2*�.H2�