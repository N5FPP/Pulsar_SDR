��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY�Ɗ����2�H��4!%��wLv��*�����"�w��2$ �e�Ҵ�e�gU\"��u䓹�!�Vn�T���'���f�=���/�<�V�(A-T�;��I����ń{k~+},E��{g1X�Z0(;�b���=5u���^�o�J~���.O�������r�MU����c�C�9�@y��i�n��"��>jȎ��@�h�T�$�Z�J�>&�����-J�aT�z� �Ө���W��c� ���S��]���F���B-���U����A��D�"�׹����/v�P@jb/�"	+���jI��ͨ�v��f@���-1gٯMvm����|Ao�g"�Bi����{���'��^�W2�̤Z`��9�	��?Y$:,V��w1������b"=P&<�$����d%��L�>�%`����,e�r��iOq�,^����ݙV�C�����
���������/�^���L�jq�6�J����X��i$[u�?{GV�^�61��-/�����]�ĵON!Ń�yJ;&�:�ލw���q�g8����xJ|}�<�G��ڼr�P�:�,d���#P��"������]̢��D@���i�=Ep�P�o��j���j��뷧Ⱦ��&�P�[�cة���Z���<s�P�i�]`�x�neR>�(ybK���g;�"��ꪯN x�X�^����B��Bd�-��_`�#ދI�����\�lǝ����.s���Q��u�<��n+� 	w��^1
1�!�p��mPQ#�ڙHӻ]������ǉ�+�%w�W��K�����ӊC����w���g�dY���(�p�l���c�O�'c'�s&�(%�QL������v�����C!8+X"�:!t��&�M.rzW����4��"���$��o4Q�����Tmf�NDr^q���?+�j�v/¿�c��(�kr�u�y���z�W:���r�0�]���x��آ���ޕ����o�g�[��B��Z{*E]Te��LԥC���꜏?կ�Sx&��m���ڦ�b�߃Bn��:�H&�Q���6���R?q�k���ٙu�6��67|��%��ج�s݀�RK�^����a�ϳ�EfY�շ�{;��Rs��(5��U4�çF)�ex̮��$���ҫ��d�l#�����0BC
ȡ�3=�'�&��h%:<�\�� �@m��U�&W�da��v��}��onW��R�x�&m8X7�"��TeCe���6N�F��6�H؈� ��1Ѱ����ž��'�)kp�(�����?y��Ds	��Ï�57$��cz4��w��!o3di`��+낔ت�G{i���+�ǃ}{�\�ݧo����]1�����3��:<-y+�3�^�z#.�*9DmH:��� `��[+)3|l�(s5m��	����}k�Ӝ0J�փyl��Ҙr�*�zDe���bs���T$�SZ=�Ƥ�c٨c�7���և-���W�_�Pԙ\ #��ؤ�TE"�YD?%�$�����'z澗X��Y�4_�b���LN8ߘ�s�{M�ڼ��i/����IT�H ����W�I��vC.]����[�1��������HN^���\�9M�m'���r�t��̱��s�QLS�.�J۲�ҿ9:�넾���R����W� �D��Q��ɜ�3q�#.(��Zk�+b��>��*?@�6�<K\�^�>9�W�ρ�	5����Qv�Y�;�O�$��6�LL�8\��rg^āI�ΫU����aǴ��J����g�B��v��Ica���f ��)G}Ú��.�Osw1%̇���+��dG�q#BCZ��y�C�� �>$I�4�"8lw��ִ�yy�UU�o@�U�l1�O�/}+� ���CCv\3���e*o�������w��c˴Vu:�@��@��:{�9�a6b����tǄ%ν���d��no�Ĕ��-�1g7;>tU�1�d��r�A���� �;N��;L�Tmz��m)Ĵ$>�@����[��W�(͐k5�u��W}a]���Sx�������T{T��܆o�h���Z���i���)p|��ɯؽ��/��ً㮿|�?����Ľ"�'Vs<�
 9X��nw��V��v|��M�F�H��6���X��M���5v�F�f�%��R:�(���o�7�Jh��}�N�k�*]3C�;*�2I�5Vt�.D쾪Iwf�_N�b4Զ{��[p��dx��(bn=d� .��v,3(H��	�JO��,�U�H�g�<�	���C
���lM��1[�����������+d{���1���җ�x�8;T#����y��4�������k�h��MyZL�M˼_3���-��+S�S!��4K�[��q����O�һ�S!�&G�����P�6��,F�)�S;���>�B#?�wP�p�FX,�>�����PS?�x�ro�x�
�PFZ�hP]��a,[@�e�s?�����i]p0wJЪKѝp���e%*�7bIp����9�����hw��у���̷ 5��Iŵ��V�����h�Sbw��8�S�a�R`���6�7F��r͋9I6Z�%)=�|��z4m�e��j�FqQ�,��t ����>i�x�� ����cU�>d��#_����[~�|�X��px��m�hK����#��g�O�� [�Y��m����Q�K�|}�{�3�ŸI�x��]])��)Z;<������������J��=�g��X87=��Y�tT���bͩ$tSf5��Z��\�4ܗ
��Qd`C}K��)�@N`О��n}�S��'Io2���q2	�"�_�Q����l�jߍ��l�t��q�G��`��f�X������r���"
WG�b)\��l�'$r[bQ2�L��t��ފc����x��t�͐�K�؜��@�U���vM 0��WR��I$�K����FPaI�"S�?$��N~�k:dl�׆�!tI����_)o�ۍ �ݡ��ae�&U�o.��7��P�h�5E��aT�i`Nxު��f��ʦ��$x6���0;�j�%�cc�����V���ޖ�����Y�b���B�u�X$��Q�:�#g���r�G����3��6o�y&�F���u���Ƣ��s��u|����U��KJڼ��SԹ.`<w�2`����d�6��.Fq'��t7vfʬrUy����_�!.@������W�f�i���I�<�>�v�q��CϽ&bɚw�����|KbE�8�@i��p�6��EE�XX6o���~1��y>��$c�����I��G}�T{#Q������}�wHjU�g(�`�~��V������������/^#���G=%��w^n��/��)$���V�O
�`{-��N� ��2*�]��mM�o�<H�MB�Ŗ|�s��e;/�T�S�u0��/.��&��fO�;��1���b����� ���Is2��ɱӊ�:3���]`��)d�b���.m�A�#�s�I� j������
-b�Gg~�n�[;'��qc��l��a��.�E�48G�
�)g٦Y´ƛ�����l��-3C�H��_�aW�ad|���[$;{�*Q�MU^��$a�ճ�Ե>gI��P֐�~1��<��fp�w3b�� >��a���F��j�>�Y�3���Do-j�����~�<艃���1�?�+.m���u���FO7��/��!��/�g4�P�� �12���!�����O�s�a��fn��h2'Ԓ�螹��X%�*`���Zs��I�ʅpQ�թfF4��[��K��^��VE��2�7_r�b��T�g�Sԩ�C����f9�l�;@0�F��&A�1`���gX��[��Df9�$*�Fs޽&[�ZHȐ��m���
Jи} o���f��Y�|���#�G\y��xUzqt�WM�iþ-'��}q�/�ジ�w�8I��k�%�v���e����S��K�X9@���]�sw�>a$`�ﺗBw҅��0
�F����`$�7Rp_=!��^��u�`1���
�fz�j^I��& ��xR#�$E�x����ck��*Me��m'�oBWn�q����T}��8K�莮kU)օ�N���9��>����| 
*3�2=��>���$PD�y�S2��2�*=5��{�߁Xǘn��$�4��v�.{ҡA�C���2&.��	7�|��k�#A�H��9ll�p2��sULW�b�\dc X���l��@����x�H�)���c��-�撣�OwZ$΃�eS^��o��tI�{�)%����Y���d�s�zq�*A��+y��g�S�!݈�B��jG��d�:�j�,C��D�2',3�&5�j$�?���������Z폌R:?�5 �������hV��[Y	���~>TK�+D���	M��p�:�2b6��0��Wb�c��G�{<�CΦ[�e���T`��w���v���2�̐*�v9~���i?*1I֌�y���~ F��e��2�Σ%�Ȧ��n��)kS�w5�[�+�h}�����'Q�t'����3�h��Ft�B�겗$4@JtP]K�-2���q���ߡCBZ���Ɓ��X�a�yq���|4+ǽ����۶,Fa�л�@����ɨ���mY?ǐQ��a�0����ѰH�B�}�l��|avɋ'��?>UD���`��M��u�Uw_ ���|��M{A��NB����/�}��w�0$Q�)��dYnE'�Z�܌Zd@���0��X]�BD��r�BI�E����GdHb�p:�%��4��s^`�u�9'��d�����Ѱfɛ0� ?�O�dL���5��L�	�ip�J�T�	�c�>�B5�ʮyK����G��{��:؋>Y�1�/��g��l �J �y�wp��eL�/�'.&�S!�~���D�Ŷ��bw�.:�`����%�w�R�>|�n��r�#=F�zԋ�A����c��FW���v|e�1�^���ʣڠ�"wX�K������RDd������:�ծ��n�=���~� �ZoL8�D-ciEF@���d��'�j��3A�œEM���1PN�=�s�J�x��&� KAG��b�h��޴�)���1�s��t���bhzq=�(��^��g,X;M�`G�-?��N�W�Do��ȁ?a0Y0}�fB�:O�Y�[�	M�n�jӿ�j>�A�+���|�۰��w]Aڲ1�v�z
�e���P�k�X��v��y��3��,����V�~#]a��n��y]ҵ޲ݕ�}��II�C;D��߉]��%���N%{�7����n�h	�_vP�{���
O]�K�i�C�EMS�s~�j'xU�C�C}��K�`�ic�'�wx�h@�]h��w��uWa����n�Kd�Ț?���Ҿ���:�x,��Ϳj7,g,��4��t1_���?gu��8-������{� M��B�0��� ڐ!~���Ó6ZP�'�Z�!�4eyO	�� dK�V^��%���b�+ػV�mp�b� �s�t�r������+W��I��:)Vw�pb�{�;���è��:��f����s�Y� M�h=SE+�cX�TS=Zyn��ߚ����j_:�y��	pf���o���r�g�����9�§�9i:JA��~D���M�b]"Wڔ ���̨�+���2+�ٻ����5���&�T����,v0w��
��.l�_���JHJ��ǈ�YH��bCP�s)�B@�{�3WW�;0����,�^����Ĭ���E���f�T���m��lD�S:
Q���2L[)G��雺��ܴ�g?L��d)T�/X�#�� ��h,�3��UrO|����]22�]55�UZ�h��.g�ɸlDkX>O0����#M<7�L�@�wW��TI������֪�>�����5A�}�KJ� .�P,��^i��h���$�zA�Iȵk��� 	s�F��ڒ�.��uN�rW�p�1t>2"���3��n�2Zݛ���CM������yV�+b\����H�?�" �!��%ӓ��_�z��=8�a�0{=D]�/�j( ���n����JL�D�{xo�Do��J#O�O8i��� K}�F��{����$�߮��O���
���5�4脎&�`�B�[ǚo�.��`zx��v���Ct��>�̖��nﳃ���>8��9����Y�I%
�V�wڧ�1�{{[�BoV��Τbl��N�Jb�<�*��%>�Q��;��L�^�ֈlߘ�"�JC�0��: �|n)��YŮ#�Z��k���� �t+��O�.=
AP��0|�-�Z]����6�aJ��;�݋UM'�^�Ɗ����ka.S�u����Ը(�������bVo�p��|�oښF���%��"I�>�#��Q���0�ϟ��V��/�p�AT���N�G��;9��dg����\l�����k������	L!;��i�#	��6Q��=|�Wc!s�M��\E�,K"��LT}�c�ROesL��p@V�K�~������ +@�ADOc��O5�Ew���\����"�"�&9��&���㑪u~a�INFR̯�1�{��,�=�.��83wE���@x�i��]���E;g���ܜ�<V��%vDS���~M6I?yͮ�^�O)�������<Z�h�b��ٌ2�\�������r}�נ���6��/��?��$�7c8+����ў9���n��Ž�GRi�Kk+�_�||�g��qA�׫x�4��]�ws��� T����:mx�>~: ���rh$M��$Է��ǇP+ ��ӽj�7p�=b��,?q��݈���}��N��e�i�����uS�;M���v"��+���K�l�G�z�"�"��/;(��{�H`�-S��$D�LI��
��AG�c�$;�9B�
��Ű`�2(h�]e����=�!��TKe[�� �4��N�Pk^/6��*�e�EJ`o�hKG���vN�e��颾�P�����B7Z�r"�K�*�����Z�q�XyG�_�-s?��t-�3)�喢k"B�AawB;.@�HY��qt7�U���*"9z�eq�1_�(��W�����s��	�_���,3���̡���U������h�A�Y4J{T�K������k��ʽv�_�;Bz�ea��h���ߙ��Z�4D~�������^Pۛ�߼J����ɽ��(��T������w�ʔ���h'�0��v�� ��;���M��q��u��&�Z*�:�#�C��R�Gori�dlClKq��2�B��F�0Y�!��9s��G�@�'�5��3k���ܾ�JB46}�[�Y���ԍ��mI�\u�i�:"
�;MX�B-C*��3#��UCz�~z
Zz�wd�G�D�('�o/��輦�
fA6��xq?���f0]�{X���p�()�F �Ў��M�s�ݒ�wߕ�,�ۧ�����E�-�>T��i�IA�)A>��)�D�P�(���&֖c��;r�P�p�
=mA0	�vOjc�;�h����*n���1Y�bw��.�b$۟��3e�N�����~��r�̪=Y�������O�C-;��L3�C�F�W`��(�:�A��r�<@������T�� �\�ѫ���<&zd�|���k�& �?`h���[em0(џ�,��t�V���*o,�E��Ůe�U]:�,Q��n���#'�x�:OJ>��^H���i`�o�.��.r{��(��t1�W�c<pU�16��oҐ@ϋ)��� �U=~�L(͚vѲ��闔�@��\���85��1��[���"�FTn썷�|0�p���\aw[�暾��!�(Ƭ��aq`;��0`nG[�"U�-5	UW�����ͦ���k/���ENY5�
ȳ|9q\�)^Kq�Ac0��k�gD�%�jj9:B�t�a��Y���֤G�>%�q�tʵ������o{2ᜫ�*#��3����I GdLځ7�Y}D�� ;T�>K 4P�AM���zv�*c52]�94d���={ ���Y��Oq�.���P�C���_��0(,{H� �8m�~T5�9�E�)9F-��nP�Hv�T? .i$® �1i8Sd�Dⓨ���DP��ox0f��Vq'a��m��C²~�7T���� �Z���`v�G
3�����]����+�r_DA9JL��aـz��w���\G]�����	+>V8��VR��A��~&������f�X�h�A���&����#/��X"	2Io+��z�����>��PU3N�c㧶�u����a��Z�lF!�u9�Ը�8z	8��!�Aߵu2[~���TL�xA���]�*�~l�㳮��	�z�G'/.�Qb}(�v��Д�*��`rk�ba�Q��u�t�|�\>Z|�$�Pw���fG���������J
��k_k��%�eT�^}(���oӦ��B��E��@=j-��H�V�K(��6TI����$|�ٹ���Oq���i�VR0�ǫ��JZ�1B�