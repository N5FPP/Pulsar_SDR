��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ���L����ѳJ���ף�6I	��7�"�D�}ے-��KpV��s�h�n]��[��;,��*��_�H1mTu�<'�M� ����Z�H�H�#����*ծ���p����*�R@�>���Vx�Cl/_G�b)�z)���e5��=")D9d��R�d0�� x��Ġ	\�{���> �Ueڼ{�g�_ˡ����T�x�\mB��޿8x][������v�	1)�X}� E�� �_ð[#�b�$Xt��C�
w��bGe���ʹ����UG٣�ɹ�~V��e"ѦΙo�ɱ���0�-�y�v��CPܼ�Fڀ�2@�E\1l�GN��Ϣ l�iRP'�ϙ����Y������ T�*�g���DO��� f1v�\�w������Z�2���8.�QV,���W��K��� *�,�J�6��jH�;�B�n]��CKxv���R�i-IJK�vC�?K$�Q�Ai�L�����I��L1�Cɂ��[�������x�9ئF��ty/Y��Tdto�	�^�S���/C'iy��^�,��)�:��K,϶>�e4��D��#��#�a��ÉB��� m2���pv �Ah���q�ݩ#��?-����A�1	�)W"�"Q�T�y��]�,�V��~���zZtˑE�qv��C������+	�i�����Kc����|���F���o�|B5Q�L�ν�!������q�"��?����z���AL8����B��<�x4|��<I�*��m�}��E�r{���K�B
�8� ��p�P�ĥ��X���@;;%lcKrʓE���Xȉ+A�|�7q���vI+@���dK�K���.B!xW�����4��P\�T"�8O��y��_�e�d��Y"D�k]3���HK|��@�u���`���Z��3���T�eY���@������z����
�fyW�5UIf���0>
�!�>c��n5�N�[�)��@4�X���ኺ�4)8\].շ�+5�W|=O�1�	j!6�mp<�0�oնw�z�����\ �8r�n7�D�텺"�l}���G`�V� 3�$�I�������~�=G��R�S�B�C�ը���*-�������W�'�ƫ)`�l<�v�1{�й�H�'���p���g%8��~bwӠL���k0SzXR���J$�/��EsW��̂��wQ)�<��9{�� ���w��'{�X��&"nYB�L6�y*S�TH��0U��U/��G��k�?��˛ȹ����a`
n�zK�[�@�{WO5r����n:���������(+�Pj��[�:H!��Ύz�� z��F�0OW\^�s�
��! �ĺ�b�!~;h����O��5��q�� ������XN��w;i}*�q8��]:�Aahr�8�hH0�fR3�ӈ	ࡓB�lG�ܳ�H�Ͷk�+���#9Ҭ���Z\B(���4�.�D#����Y�v��qBT|�Z��G͓��B���h� *������b�UL�������l�J� PƜ"���ϣ���biʣk��� 8T���Á.�o�0S����
�s�����5��� ��ő%@�n?7J���z\�,E�Ne��Dϧ�MC�h�}��E�/~c*�XϦ\�gJ�	�ڤh%<����T4?g^�Oxޑ�9$������j�t!�D]�Fgq��M��{8v��$�K2Ǡ.�|�`1����'\�AC�	��< FY,�x+��_��꽘�C���L��ܞ{v�S'�4k�c�{X}���R	�8���:�}�&� �T�@mΕ�^�TjB� �5�U�T6�x���,�m#/B�'��~D���bO ���(�ޓ���E�dP��-�%������r�`V���wU}�����"g��u�N��{�1z���Ԍ�"��V[ж�E�9>Ԯc���#B9����)�_��B5�]]�iY�<.���:�F�bu��^�Ep]����^�G��{x�<�*"�k�y��Q�
Њ;��d���pn�S���劦�i߇�п�A��`����X��:��EݼDa�O��|���g�h��z��s�E|����;T�_�9M�@!�l�?�D�ـ��y"�[l��yL��1��-�7�+��8Nc�-�wr��^����(?7�Q__!��=�y���ס󴶲�c��m�o���y�0���i�)�5l�/W�FQ~��	�yo꾟��k��`��m���m�nS��|~n2����X@�#h��\�'9PV6��sj�y؎2Q>�_�d$2T�6����w��0���9��ѥ��z�pa �4��8�������Ki�BM{x*9O��bj�f�|�7�w�8L8@��ć�V֮w_����g��j�����򄮘��%B�ޏ��㇮*).�Nj��,�~�� �8�����]�j��B�F�X�I��-G�$�eB�K��N�@�S8f�V�آ�H	ٙb��P��=J=p���:U%*�&���A�f ��5h?Ϥ��:�du/�a՞*l.�4ԧ]�0�<�Rs�<��q�)URTI{�T*������`�ގ�����K���ܭ�ލ��=#<E!^|[u�za�*�{8��� �$h�T�L�K"h�O�0�d(t���-R
0�Q���E�Q�l�ԾHL�W�Y�HZA�]�i?���hi���;/�ta������,n�4����������W!V���E��e���4ډ�ǣ�/,Hp\Oָ��7̉�
nS�b|j]3�m#EWZ�_5�"�bk>Gl��P���?����#8n���f��/�+�Ts�?!B(�:�rx7��")Zn��PD��3ۣh���"j��z�6�B=�^�J�!�_�� NT�)yt��2B��b��%U�ca�fAԋ�j�j8���J�9���o��Ǌ�Q�=ݰZΪ �<�+R���ԇ�HEF�)�����K�vW�������˄�uϼT�F��_@b Q���#�Uka�8��V�@�S}�G/�J��Zo�����bMU��+~��I�R�5��/�~�5��D	�\ ב��k3�B����)� 8]PɌ3_���(<ԫOJ�B`q-/��.�"��4 ark�x��`a�D���_���[�Iw!^{�1�l��}j�@��F�K���EMt�˅�}-�S���VI'��>��"�-��P.N.O��~K�]TN<*�WV+HȊe�{[�����5�؈���g�����o ����-KF)�bHH��Ȟi���5���������Mr�7W4�����^��<��t�,��?�ڜ�@|�5Ș�bC	A����r��k���	��H�=/��O����T9|�O�
�ȣ�b���� �px�y�Vt�S~�_rq���3��W~C����<K?2Z����0���#�S��p ���~��H���dCb�8	O�F�dm�/�߾c/oN%q�oh!T��ױ?�m����툻!����N�� �kZm���6<������v>9�Բxv���!9,]�Y�G��t̥}�~����s
{]���&��87�Fg	�X%��I�=��کU/f���P$a"�h�8Z�Z���F���� �'�mZ�#/L��an.F)&�"�M��i��Yb��(@Z��rYkI��3�p�ٯ�|�3��$m�P~����!slI�@�W"N��l���]�J���FPR�z�_�kD�x��Ϳ��w>��JY�����!�*��z�ujC���deS�_��;�Q
�.�[��7��?/t�WF���V0�"E*����ǜϲ��1k����ϑ�dKZ;�T�[���;��Y;d)_�����O&t���[q)E���<���ɽ���i���MH���W9�r�Mﵴ�
����l�~4WM����{^��ۉyy�+���<L�E��!J��r�v�to��j����#7�T5��Yf�;�u�6��(�q�o�k���mU5��G7���d��j��!�{�j��w���h���xN��k�ASa�!bBD�����=M��/��'����x��f�p���
�t�tb�qB�G���R��s,#ޗ���1ZO3���mӎ�,VC?+�9(1*������C?�Y�.[��z	�Cp�S}9�l=hV;��h�����Y��?�K9��E�Z��D5���1�#�����*�� ��휨!�� ���@��nP0S�*��<����b��z/��4�0;�w�|��P��jt���4e������6.ѷH8"�v1���%���?V�0�����[Rp�ŝn���vGu���()��/P0�Cç��Q-��p��zCR �%��]�5phT@+B������cT�{�<~q8��:��9 �����i;��B���غ�7ëX����-.�,�n���,�[�Y�}z�H:�"iX�$���q���I�����`3�I�>|���nN-���A�/��JǮ�ʏ�(ب�7'�Gt�Bc���i�;�2�4���A�V���d���vKL�y;��[�]yv�l��,����{:QO����pP^d�>!�/${I0�%w���� {<>L���f�����p�������R4������铦˟�<�-c��'��{�����(`�~?<~�����r���E#:rIU�9�%?��YQ�O�K%W�2�	���5��q��Ĵ�D�0��:H`����o�?�Cq�~����*��JM���ڧ�ߝz��B�����gAq��:(b��fU�5�Iߐ���l�WA�>:�/#k,,t����7����v�c$�j]*�i�FD9����윞�Q�FYKI�6�N�]�����K~v�V��¶�oNvM�qU?��th0�/b;2������y�>��°�&�(��#@S�%lC�GuڕǍ^vX|3C8Y&(U�qNi}�ߛC��K�8� ����F�+��JZ�� �����ni�yB	Qw��z�'E�#$�Fzox�����yxw�i�����~G�v~2xf�=�������Ցe��9؛�q��ē~��S����P�	��1Q�̜+�ZU�����p��˦�a}�i��b�������D�c��Gk�i�v޽��7ܶ�M���)oLe�	ɧݮ�~�c)����	"�Τ���p��m\�d��/-ȇ�MA�0)3	A�쟧Jt����4}����C�ɡ%r� _p�g��̏SC�v��N�-�o~�ykPp!]��]�Ǥ$R�1�G�L���͎���?tx��`L���Zo�g�T8�z�"T*0&1���^w������=�"�\���Og@9��l�H���V��t�����ަ&Ө3@٧8�e1��"�"[�)ar+��l��^�4�������~�Op, &	Vx�A�gڼ�A�J�o��sjg�s@��u�� �C��2R	�����x碐]+��r	Fn�����=��͔[B���� ���̣������ܨ|������S�4�Ww�4��=��D�5d������5���d^���^���^)�:�C�5��|�����1*t�M�Y@_z��q���,��ۭ���lז�G(�`,+I��P֯�=�%��� [�N9�=e���}m�l��w}5�Q^3�����Y���5Ͷ���g���G�{S���G��$��Y4��z�J8��&%ޡ�>K������Ģ����,���������R��Wf���nZH���M	�� n�:�iÿ<~$`����.| �?;�j�%Ui���&ֿ��t�)��}���'[�c&h�C�����Q\����U��n�i$�X����R��� O�3�
�:�t�x7�ib����}lD�Ç�'*��5�k�G}R�!^b�M�K�rz�2Ɲ����*��-`̝�ɏ#la+�y���@�Rx'M��U�pOW(׍��K譓m(��������D�7�����,��=;C��יAW�U+�yz5� ݜ��y$2�#�i�nݕ&���f6�`Nk� �#^�G'I�����-�w���["jB���
C퍼x� ���l��y8,��i3�E�|�k�<�)zc�0|�����$I�<6��t�Eϸc��Uv�[�] +�ܶ�	��<�~a�P��gl��_q/~�e�#/tUO��wxc�B��|7��;3%�`Ę���vz�2̠G�Wt�:���`��{��_���v4�4單���g
j�;]V|�pv7��;"��U�D-��0�ҁ!�Ѡ��@!r�._&= �[#!��/o��-5 _ɳ!���#��^z3���c?I]�| �� Ne��Xa�q�8�����So�c6�����땧���T��,��@R��8?�0�25�(z4[7�C��V��X�{�r�/�U�
�zp��mR&jc�j��q���?���ȋT���n������dk�4ō�'�:P/�E5�i�Z*�׹�94��`,[��8gPX*��q��[��Q�+J+�\�/"S6�w�-V�Nx�VJ>�%���Y��!N�]4ں�%��pd�Z���$j��³�,���V�
���9�s�l�r���L���9�"l� 7�	����R�FS����ILk�:���j��P�����rH���T1w�C8��5+A���缜�i7;�F��0B\i��"[@�^Ҁ�=4W^�	�1[`�d�"6��v�X_�NׅȊϜwd=p�����?@l��<�16�KZ�ֿN�˱^-xR���qA�S&Ř��v,�`ժ�}~"q`G0��j�x~+�a�q#�^<�>z"�㱏�Ǿ�%�C=�`�Щ��"�D�rܭ�`f(%��
h�	�dG�S-�p������uc�Eq5ݲ��V�$.���S;�柁@u��g,Ȋz
GU��m����k�?��'#��GX���q���2���x�<El��Zq#1��Z[e+��YAN��L���Q�u�9��k#[���/O�p(N�L��0ˇ�'�-}�����b��(��:V������l�h�����![;2ᬵ��k�B�0�e��"�!VZ��cGt@Fi�!Ӈ�e r�q��~��?�+Bh�����yf�I�X��K,��B[g���"2U�֋oCv�������p�u���Q��zvHn��C�گ���tU8F�*L���
�u�O�#�';V�2��a��0�q-��b?[����q�d�]��=����K�
������Y�k���i�81�t�����@�ƠG@�i�+h��Y��)9^��ʽ��4w�W S-2
_I?�/b5jh����o���ڐ�����ݍNsL����g��+[��N��ע"��H�n+��"QM&��iqa�}��vP�tyx�s<w�{��d�7��p�)S�թ�:8���úI<����V���cB���i�����HB5^��t }�a�U��/�,1��P9�S��&�1kQ�U��UEt6�t�P�;߭��<���z(&�3�)g6oz|0�(�:�贈�-��ġiA�Qf4Mˮ�T
)X��C�b>��
\dc�~������B��~�0��G�=kM2�Qg7.*�1Be������ɕp�oWB*�G0|�=�~��0ۤp|i�t���n����z���:����3��~$"���-Hʵ?L�dĆՓQx�������	�]qVy�#(�i�������E.�H�g_�a�Q��]gxu��~��k����5DSQT;�����7��{����=�\�+�c�h�[�g:�a|Dݶ#i�^9\ �#�G�>8!嗽s��WCV�:��Ɂ�u�kʋ`��"৿6R��-�������*��a�A�v���v��T8���wa��F����y^��	H��Y;w�
Q��	��*\Q����)�;�Ԇ�%�>z���(�����gL�y��a}�M����Q��MkPu[�}�V23�P͠�6.d�*�]M� �M���aS����
O\��9�]r��+�>�-z�!�N�:�<�Ny|G��&���m����VJ�x7i�E>w&i�3�,h��(0զ^��Fכ��|�lL�`ʹ����vc�*[�&����n��~Rz����Zʕ�qO�h�h�,���N�V�_Fn�Q�mǶ��:���+�b��(aʓ?�%��CG�R���Q���w��u�q��
aE��H�g��S���	c��D���`��QƩݏ��bk^#Wz-�[Vӌ�����n�=�Ix �
�!�{w�H�;\���P���i�d�ַ�Tc��f�)&�&�׾�d���q�L���Z'��A�����m/����c-�u̵����$�E!6zEd�X1E��j�� WD�rD�"���2T���¯�ޚ$�@�����k<pj�R~A:�X8e#�(j��S��<Heӯ<H
���t����䬛acqG�TK��F��h�q�*C�M6si�DFr�#[!5��Wyv�����]��u�z�o(ДB}���o������Vgsߟ�������L�8J�?�=a�i���O;�d�oud_�ɾ6�By�JrT�d��VEi�$z��1،M>.7�5��z�;�[��~׻S��g��
�x̐	�q9"�4�%$ ]��'\�#A[�\�RGP0�Y`�āJ���L5u�N�����G��U��$�A~��ރ��B�c���b��%T;�f�"݀N4P�&DU�Ҽ�?�w�Te0|'v�����%o�7���}ɦ��G%�W9Y���Ԍ�<��"��"Q1ϊs��['�q��K�}�.�zFG»p����4��&�����a�izIZŰ�`f��U란�2�ơƭ��@GR���h����B�p��2�g��l��zV�5?l"������dr�)4�r���īj�|e��u��]#�<*(cȣ�弚)���d���g�Ʉ�2sJ�+��ȧ����W>��D0����m21��q�UѦ�.ZO���t&�����+W�7�-��fG�D~aL}�USA/��e8�=M�x�"��烪�w��
^�`�������,A������c�8��NWK$5���{Rp0�kem�����y-h�ݘ%(��"AV1��u�7�οP�e��Z�A��s��z��������l�@�լᰵ�f�
�
���=#�;�~��-DM�p���a�=M -��vz��cۮ٥W����`獢�
�qU��2;��%t�$�<�jȩ"�,����hiB��H�v��g����=����8(u�\�?�i�i�n튈|��D�2̎u�Ȕ�/��1��_e�OR���>� ����=C[*"�UǷ��=��;�>���%�1�_�h�s��E!�Ɛ����n�MA�x%���¬W(�����t� �"h�m�V{�]�/f�W7p�F��1b�Djr ���QĖյ��.�?������~��"�s�'��V21`T���wU���s�Ά|����x
5⎬H����2�2��q�
�$����n�@̦A~7��M�O�"n�4Q�wfغ�:��o̉�pe8_$S�E��Y�I:A;V'B��N s� '�����a{��<�!5,�t�c��}��y֞���Cg=�U� .<@r˰�O�4˗��i��y����KuVӲ!�����xO��!W��,����St՞-6�#K׆�"���l3s�������a\�1gY�O7+�УY�&�^V3z�Ŵ����U�[��ۢ��a�!h�S���R>�aP<�n���a5$���W.bu8&ր�!
S�I2�/�{I7&����HM,�kI���t^��96�Q���LY[�8fSՇ�z�fwJ�T�h��6�=��"`�*��j�1�(G��"��:m@}!�����]��,�r���Ψ�# �?����M�t�����vϠ׬�`�Cܩ�ˌ�U%A���z��("�闻o��[������L�T�A���sN��bT��P�ߣ��U�R���C�����-|:�+�b�nTI3����xE����{�k�;¥nFiE����t��%U���i��1F{���Gw���I�c!�K�cr=O�&��6�*���=F�c�i�x��{��1�K�Se��s�sJ1��G�,c�O��xV�>�_�aѐTOɶ��k�!7�m���|W7�Fo�7��絟�9s[�&n�o�8[�l��a �e��s����S�������� ,�����'nGP��=����En��Uֱx��Èd��[���bz�{G�����A6�cO휟]Y�'���o���i�9|E��o��_֣��KW�7���|\�1R��ֵ�����Y[ ]�檞�Q~cRà-v�gz$)�s��+1�
U�:r�4��Zo�����-޺�l��EE�{�b�C�-!1*�xD}�����G��k�x����ka�0��I��/G�@ňѐ%�5\0��U�����L�L���p��^�C�
A���[����0��Q�fH&����i'R��n*X�U/Ɖ�'z!V��P��U��qd7۹y�)�M�� �����=�9��Ɩ��ˠa�ؔkYKY�Rz�C���'o��&�aF��X��_]�V���Y� ���]I���.�1�3�D�Ǔ���F��S���0|���E��W�X��D��KVn�<����h���(�2w+���gH;E��[Y��[ز-/�U�?���
�^��(	W
ӄ9Pʁ�z`1���l�o�#��Ǧ�?�+��o�ޕ��tl��/H��d��A����Ƌ�KHA����* t��4-k�>E��PQ WW������*���q��bb��A|^�AΠ�ܴ�G	�*.�=�<L~��?xN�d�2'b@x���A���c�-඄V&�����M��
�<^�?�=��a~��a�B�x�>$���	�ղ�T4�|�d �o�׾3IZV��R]�'���
S:zh�`!
��Hj�:�8��0�������"�<�Z�v�j������zr��F��E�M	4��7�L2PSd�tZ�ꟗ�6s-O�x��O�'dP,T��	x���.N^!�<�ۮ���,���o�sU����C�_7�Gpٰ'#x�o9^R�'=	�3�T�r�\Y�M.���/3�a�G�̣8:q�a�9�!|*9�R"A���H*�l��nu�E�M��k�7y���E�d����Gwk.%"ؤC��U�"J魦#�y��V��l@u�N3#�����ʩ�U���>{�x�ې�,���M6��Wt�P���/�0�\p>�����_�S-y��
���;F��r�ٰ
�o.�S9�0��6t�E+&�:Il4t� !5��5�a�����N����A��.��kZ�R��r%旲.C%�kv"qoy�!��Y�C�����j�|l�q�e_9�r�E� �9S�b�Ӥ��v��(�e���O�	x�F���v��'7V����Ҭ`�sѳ}�C�#��m�a�ȿ&���y��Vw�f1ŋ���B>p�W��6�fp$�cS�*o���k�c�<�UUeeU8�<��Ɓ�oW�aV�([����3q�I}%������zj�k��	�b����X1�@Q�0���)���4�C��N�>=%u��J�+"NU���i�=g �2Us�����#��})R�&+�W��9&3��)��J�k����p�5qL4��B^~{�n�Z[+�i͜������c�:O{9�L��^g��s���3pyb�����z8Y�|v1UA맖������O9�[,ݮ��K%���.$��~I߲�����5c��`�q 8�[DtD�9�����A�`�47��Y���-�B��}v�{��=IM��?K�S�:�ڋD(�2�	f4Y��3��$���*Ů��<u��tSe�sX�E�ŮGN���h������ ,��f�gv]��?6�ϑ����er佁�{�rB�uZ�M{u�	���!�Y}�`�aP�����ٮ7�z��!�w���<IC�3Fiv	 �AԪ�l�eS��n"��+�On��'�<:��*���	{���\��m	��`��},_��%aj�u8��OF��e�����)�Ru4�B�0�R��5{&��4��>�H"6�Z,~rU7w5֨m�?��6�C��a[^�͡-��t������V5;��7�C(J����N�
��2�d�A~�筌/s��T�ev��^����G�	{�P� ��Ӝ*�nƵsV�q}�џ=e���w;$kR�S���@4>�IAЖ���=�Gv�6���ү8��g����ξ�۵��Ћ�L:�>X?����x�$@���5\���Hˠk����t�vt�����_ζճ��&�,Jb�!�)���3*R�j��pBl �ß�D��D�=��7(
��?t�J�lFT����^�ʤ�K���Qu���2�~���f���f�sc�Iã�`��-w/?��A�Jm
Q��Z����ʻ����v������E�?��:��{./���&ʁ�{��ro�LځĨ�����FMV��޶�x���7i���t'��k@W����@RY`��� B#ڹ�<��e��,=�^!�|g���P�P�������=�V�WL#o�Olq��JaF�b"���HR�(�� �@͏,Y��v��į��m����.��`v���~��J������]t[���������g��Q���k��]��u�
X���-7���d]G%��aR�A7�_�$�L�8?C�������[-j��N�P7ᴔ�諿)�F'�*PKK�@꘯��9Y��� $�d��]mD�v�ͨ�%l�+h���J��q�ҕ���$w2�j�n�fx'󚕶�����B�g}>�{�T\[��GY �0��̚"˵+�[a7�m1�8�F L��`�?E���3@��=e�L(|v�|�Q)��hR�ڎ.F�<P�(0D�ه��Ө��h?���K~.i�_�L"���𕅹V)�8��R6�M���Jt�ބ dh�-4��gNQD䜀j���� 8����W���>�s�g�i�9�}�)Mo|�wK��e��a�w>�E���I� �I�1�}^`3i�.D@�QS_�D�$�?�<a�=��̨��+O���9��]���l�π�_;�H��篖��6-��B^�p��W&�/���m�i����Av��ڍ�,
 �]�/K������#�Q�%�&��z�ڛ[�c+7����s�`6�"�rx�&�"U�3�5�Շ�'�D���0�1�'������:,¤�;~@sI_�R��d�r���>F�Ek**n���(���2���J�z>[6��y��_���K�)	��[���A9�*ש��^�*dMN\_ J����̇�
�Q�U�f����`\zY�vd%��A�ꈜ�=ꬓb~��s�ve���n���ߏD>�^���c�4L�O`|Vj �9n���[_?�+(�{F}�c�Tm@Ol���uVS��������Ebc}�/�qIUk	gkcs�KV�I�\��d��g>����5���YY=��|����� B��*�Dk���:�%;����o�Gw��m{`�`�Έ!57��M�n���F���=��J
�`FJ;�M:�B�x!�]H.��/P���R�<^�^���(��yZ���e3Y"���_�gJ?D���݄��b�܍��轜�F�<�۩�3A�\���f���?D=��6~�97���`�g�xZ����H�g�� ��Rr���iMT[���}�>u��l�-X�u1i,��O�v���"��z��=�n%i��I{4�C�' kqJ4h$E�tuh�2�ƭ��ﶟ�w������� ����L@�����G d]r����]��%Ke�վ��!�f��#%�پS��Y��ʸ�q�����|���z)����wl��C�*]��I��1J �h�Y#�&F"��f�p)�bT�5A[f�O��
�N=fC�r��z�v����������U���wƥ���ߑ]c�h��S��2/�5׽���$��Gc���X9D��@�}B0�sP\�̠&��~3�S������;����?�����e#�����-4�:����ΐ�x�[�Ћ��p���iÏrՙ\S_��<�i���e�N4c����F用.���J�p!2^��_�v}:\D��;�Kp�XKQ�AH�L��IUI�2����J��#
@�N@�y��E�$�$A_}B73Zցg�����Y/@4E�K����w�$�W��o#_�����;W|�p T�则d�;�ӳ\���>����h��Z���]�<�K�:P$A�v (��n�x7s����f^+��k4;�Ɗ�f~q0�<��J72�Bםs�76��O(��ʘE�����+�����ޕ�c.����1��ppcR8��Wq7�c �˴[���v<���Y 4���D���� ��CL��b��9}�P��b���B0�W<�bu{��SY�3�w�,��<���? ����"�w�� �B��)������>�+��;�4 ��N֐�W�O%�ǔ��$���ӫ(�ؽ�ɥG4�un�¤4�F��^顤�rk����w���͒�jW��¿��<yU�u?�g�W���o;���Q�uAZ>���xW�

�f߇h� X��G��o��g=~���jI�pE=��f����14,�ɩ��ܨ�۵�&ɝ�jf��KH�M���)������w5 ��
����z2X#x� ^^3(�%�z����Y[��]�5���V�Lwꨄ'���4��`=� �3��r��~8��u�s�&D�,�����IP���A��=��xǩ$w[�Ot��=8���������D�ߚO[N� g��;��Z�ß�+<�6�����#WE��ꥥQ��3��6�0��q��5'G�ߜ�g�C��u�%:��Id���V-	9��<7���u�S��B�؃p%�4�ĝL4���n�pu,�/���-�'k���.�[^�ݑ���v�Ť��E��۵���5T�u�x�||Ў��0Oz{84��9�C]P&� -O@�*��G`G���jЀ*��Ìki�_f�@�N�]�;��Vx���/�}�HR����z���a �bn=���w�{b�ح9ӌ)sT�s�tB^���� �υK�z���L�|3��$��{�X��K��Jk�ـ�����Y�fr��P���Pn;ڢ�u�x�����{�u����3vBJ3�!TI���u[ߛ���;�ܵ�`�r�6�{X���
4�dr�Q�!��R�@��tx��:�%��I7.]4�p�na�L�٥+�򰟏/��u��p��k��F���%�*d�B+�.�C%+~��E�Е'�<���픪������wuG����s�*�Œ���;y|��F.���`�N�����ƭa$!g@�����u� ����N [��4�l�!��'FT0P���ꋷB�z��p3���¨�9|�1ce�h�p���G������6Ir�<4Jڥ�#�p��a��k92��UAl�mKhҚ�؃o��h�ȶ����N���O���w�:X�qۘ����*�'03�ҕ|�q�몀��y�5&�L���e����KZ`�/|���B�����5G�	Lq ������?YN(��(:���15>�Y�Oq�>�hǂJ���Py��I���MZ�k��/�&��9��A��eg��� �\�&��_,՜KLKZq�7&��č��_�gM�n��@�5��_���ѷ~< ���<"���U��Tk搁�޸�N���4k��ߖ������5�]�qw���T���}�;g��r^G�v
>st��6���:�幪I�n�'���\��.�����g�H=g�k�V�mws.^Z(/�9�`�̺��~�X�2�F��^ �w�bI�]�kaC��iu�}X;N(���9!![:���)�J�x�5æ\�}9��a�������r���1�CŭX��>*&�]u3/6Z����G��	&	�"Ŧ+�%=�X��Y~�`F�z�eӡe%P'Q�3��r1؝N1L/CT�6�ՠ0]DR~��� ��y7�Nő���6�C��@����[���������x��\���	&C��[;�-�q�&����ݩ�l�u���!�g�+}K߶eOh�0�N�L�A�緎,���e��~]-�v'�S|+�5N ���H���p+�Rd�Ŋ�	>�b��`S,�w�3�0���9p��F(����y՚@s�z6?nC�y+}`u�p��O@96�QŋܸD�b�Z�So_���; c�1�q?>/x��#�x>�mjf-��_��A�r��g��:DQ�]�����>K��b�r�#�A����P9��	���Y m����F	q������s^���� �
6��	�O�%���;0�&�?�R�M���'_G�$����]q�)q�KN.�g����lz�E�s��v�;�� NK�TCʥ��(	S�F��ۡ߼�Rn[ҏ�I���_�sIǭ���0�G�c��-H�A�T6�>O�Z�^��,Xd0�q�o��}ר�&z��3���i?�%��v��$���(�U���u��P��W��A�eG�v�@��|�[��4�H�p���a��^�������X�ۈ|Q�Ѫf�5�|�	�шa1�pK
)C��:�_-�
����3w���t���g�
B�;f8S�����6Ҥ\��S%���a��,Ca�Q�ࣼ�#f�O�7�~���e(�Lz.噡�ٟj֔3��W[Ԏ��s��zR�� ȲW�ź/u1|s<�IcO��G�]9R�v}E�c��$��/��lQ�\�m%����!�А~��;o%M��8d��T:���Қύ���d_�S��oUN��#��&�!y�ڋS�@9�Ġ�	|�
��ĀI�����CzS�uOjT�Ek�L#�U�נ<D�b��8��%&�R2D�dDF�lz�6y��N4Zɍԁ��~�E0�?�@)t�e�t�&e��M��ڬ���iM!�4� 4U�T��di�{0'������k��=���M=��v��OU7��K���wH�#!���Z� �ӌ��.��0��~P)�a�t�(M���Rf1�Nc��]F㡴 L��$�z��K<�[I�9��z����E��{�����=3�L��o��^!g��;�qV�d^v������]��kS59�4�lz2A�~��B\9��H���}zͦ[ f�}�������ѫr];��"���������:o�)Uf�*�vt�*�[��(4�����S�`�p����t����zJھ2/��*ܣ��QY���T	u6���.�Ĳ�r�B^S��ȱ��>��qT�o7���.CV�&R�˓g���Elf�h�~��M��ٿ
�~�2�Bh�����˄�%'ӧì����Q�`���,�.7������ƚ� h'�CA�~���,鄵[4ⅼ�y@HXS����3>MPWg��e�SW+�Gƈ�ڶ�0�ɀ�Ā���>��'�@�"�[{�TzUR\�;/	����i<�˫ԞP���VڶH*�j��2����&և3�ʛqq��D�65���v�I�h�n1�E��
���c�NG2�)��H#�f��C���ꑄt��p�~�d	zL3�X��ٰ�:�<��I�M��:Z�p����]�j� �2�#�����}�]�٥��̰�/�QUq>,��+�)Y��M�ֻp�����}͗�~��x!�z8T�q]�ʀ�?-��A�S%����A诊�e �\Sd�a]kg!�{�0,-�(.9 Tڎ�)��-�^�ZIT�|��+��)��}qn��.�񉾅��R��m�I�6Y�J�vo(�?��$�
2����x:d�s)��/�k�R8�n��ןA��%�-��& �>��I�A(�A��>���#���fMj�/�����8L�`�pja� �]w7#T�����PvH��qǉ�?W�_��U]@mm�M0��ӉЛn�z~^�f}kM�eO<�{�
V�(��7���j<k���l��Xi1d��,50<��:��S�CF����;��wčނe�wsFw��Y�ꝝ.��C�&?U�o㼸;��eidq\.Bѱ��s	�@{*5+6FF��d5�� YTH9��W��Uh�Ԭ�����!��	.H�7��KW
|wC���h�|���U�B��X[����U($���\I��tz�_5,1Hd�" `ߌ�R6\Pl�u���uoWW]F��u�1�J�?T�}�8�(Ы_)�z�����L+kƞq�R�������`�����g�c��|�~��ɇ�)4{ӓ�c)^��y��}�L�|�꠩Ӎ���}���y��23��G�R�q��]��a{��@?���HX�"=y�OQ5�ѧ�
hĦ{�C-ll��j�o`��k�(
<��y[��Y��_��D�-�ퟝ��arlֈ2c��/�&`1V���m�]ԑ��x��^O!�!�ر���)��e?&e�~H{�~A��RO�6�Q8G4q%]�m���:U*x)�͊�;?"F0�-�������<��
��.�v�J��8�s9��T�_�8�0(�"�'�
"�5�)0���d(BwV��0��� �v�;4b���$tk���k�;��� ��p�F����~Nz�v3�@�jYTvb��B*X�+��8�����VpS�#�ޏP�ZZ�L���=ȣ��{����ճ8l��K3�+/������U���~��l[�'���f� �I5>�'�L�^�U�;Ś��c�G�Y7B���Kg	������ �	���l��A4�e��]bT��t��r�e���Vb�\=n��`�2ș��A���Y�%+k&�Y���!#̩�_�, �\Zܾ*%&͙M�vn�\��KaY��D�o<�����_$��J����C�U|B�W|zΈ�7�ӕ���!�M���:�&�&�Dp����:2ͼ�M(֍
�|��+>�o[����|9U��B��|�"/�����q寙~8��Z��n MX]�:��9�&��ayf�t~ko)�\/��`{j�����z�j��Gn�p�~(�<nu���ɯU2��p�8r	�.bߞ��?y���)E��&�KY�ô���<J�q��Zg6ۓ�|��d��f��Ta �y,�75}�]~��/_#��zs��'>.	r���9C���������(�B�[/�8�+-�[^���f�}���t�J*C�����9�x���Z���k���\����Fww�P��)��!f6
ǁ��T��S�&3�kEY�>d[�t�o+��G��� ��rɡ��)S�g�|�۽���U$�a���;=�y�|���8�+���W ?�g8�욼v�Z�ar��v�wEJ��<��E����a*R��*��W��;*Zhå�b��;�h`�c�ŦIbR�0��j�ф��,�w��f�L������ʽe�a�TWh�0�@��O�_I����d%c~:!�l(>���b�:�uZ��o����f%��^hWF��Dx�OU�ֳ��YH���g��h����ذi�������_�:���;��_M�`y.�jH�Ļ{h�&E�M�dL�s\Q�{+/u"ܸLY��^2��#�,dyF��W8d�$�RZx�����v��
g�\��*�� �6��Ŏh��h%�'�<n�|�����{�h�g�e��jx���kl"*�/!;����@�1���,:�ڔ�����Z_���uN!�+0��8�v� T�cګe��	7=Ơ��م+G�"\uk�����E�7��N�!F�4���X�r�e"�(�ܝ�{�(�#e]���0G�aD��"�)�^���0��d|��2��gԉ��>���C@��İ�!�3>�0�I�t�����P3�6���ж����wG.�		V�C�c�F���ȡ��V�U�Z�k���՗	��戌;�H�@+)C9��G�}�*���ޗ�j[E�'7Kゎ!�ip�:֬wn��¹e7�������\*ҽx��(��T��e�>N%��B.3���;�(q��Xb��![�\.%.��X���X�~��x(.�4�Nu��Q��˳}G:BI�=x)�7�ށ�39����]�2�"V���a��=o)"�棉i��ϻԵ"��K~�n^+�E�qMo\�B�4�R߇�U�n�=��c�,e�b���c,.�ٴ8@��?�X����1G$�����ל��t+9�A�-^�sF�D��K�|kF� �[��g��� ghr�2|

;���4��s���r�x}�Uo'�K[�*�G�$/Iڊ9�$<��B�˥U��F����o�o�^c�Fl��('N8W�*���txv4aFJ�L�������˕$�H��]�+��^Q~d���c�����a #-޹��[lo�)9R�XْW�����K=מ/�g˫��\L=?,I��]9Xc��FI;��4&���S�W'�Bҗf
++�d[�j~Gsq�j���] �[+8�i��X
�<�Ƨ�z����8b�_�f�%��6ب�N����u��eZL�c�c  ��2��; ���(�����Z���V�*o���~w�Z̰S���&�n��=6�0{ ��޾�-!��`���}k51/�5�U�����х�N&�a{�c�|��ĖY��W�8�7+���l��n2��=E��I���p��e�yq�{�Mٽf�NA��C�#�M�{�$hB8��d�����d��꣸�9,���@�?-�3[߃���X�e:"�}��ԋ��&(�~U��IK�_
�������{cn������nQr��T�H4bPW?Pp����r�ie��nz���y �\��em�ò�0;�V�kb�Y�]�L2�S�o�Ci;c���=O�u�ȳr�]��{����,y<�T�
��^���\�{���$=�ݵu������2<j q��mlˋ�ڳ������I%^�ֽ�_M�j���G=��\��4��p����������j��UJ�d�A�|��?��i ��;-�/�8���{���$�O���i!�.e����#Д8	�!��t�E⪆C�&��P^8�9Hf����O��S����P���]D�1}$nx8������E���:�%�g���D�\�	�y��ޜ\j!G>��Nz�]Ff���!�j���חKP�^S����-B�{LL`Y
J�&�G���C����z�	o�=�}�i�ˮ�'����0Ѫ��u�_�0n&�V�M8�j��2�&�:h��]BPtX����3���~HX)�Z&+���t�#�D�~�6�ВN*�ǭO�
Z��c�
�.����v����hnK �n0�蜾��{�0�g2J=V��v���ؤ��gٱ�]���`��ҏ�b��Y�i�+�����EUg
�I�R�a@4m�ek��KX����_ޤ�{{!��:�t��ICI6~���k�f]��aC�2���\�8�꨿!��=�.�}.�cs��K
S��;��^��˲�܈)0�*he%�e�����~���d�øqr@�^�JF�J1��я`/R��+�6��F�k����%�������7t�]x����53fa�c&CK� :�T� �W��Z!��сB xp�����an�����0*��,���:#jQ�tOA�?�y�@���F��I	;T^�%�Z)X|��Ta.�;ؚ9�g
^� G�q�X�>�Ӿ0�4��`�rJ.�� v
�I���螫����'u���a�i�����c�� �|:�\X-�-����{a�T�*�$df�����J��#Z����d"2�}W����Md�ܿ�C1�7����X��d7��1��@��M��%��".U:�Q#z%��(g�90B�!��}mN��E�6�|���rŖц��A����b��j:����p��#-�%��4���QуF���6��[�gi��+M���|o�!���q\��5ٙ�dsBz�f}����zT'?��l��9�p�)\��Y�U_�P��923\!�E�S}L�"��1�� s����6y�yFF�x�M���RM�B��6����g��8�	�+��j�=$�u`̈́
0���K���MI��|�7���r���
B�]�aE�?A�b�� � %�}�#aBk�O4U��>��{3�$Z~6�n$�0��"��`���8�;p<��q��`���j�Q�a&�.>�7��~��J�+{��wp���EoL))B��i�����w��G�REU�e��S������2.ɵSF��)p/����u#�`�O��+	��Cyc���GuH�D_���]�NT��'���w�.�AgQ� �| q��PY{�۱�O������E�ji��@������~�h�Z̸F�f����@#k.��2�L<��`5Z��v
@�0Mq��5��f�T��SZ��64��z����03y�˔��"�[m�/k�L�c�y9$Z-L&�c�'�?������&�y�ٰ�7����	t�#@�z��  ��`����W|�)�ͳE;t>�L����OW�^�z�=��R���WP��d���=9ek�4j�4j�/l�^C\t(�֘j�|����CɃ�OwyFEbb`��g�ޯ�]<���Z�׭���
�P$��UC�ۈ�M�y��/9:��Հi���V�g����f�.�����E��'*ަ�D�؟��x�r��LD�]��a% ɟw�>$�4+�kǻ�������뮡l>ɻ8����H �´�>��%����q��UڒicQɵ/����uo�-���!�A��=�m{;��@���aa��~��VEaD� gH���f#��>����_�3�
�G�&�}܁�!����܅��=�hي��b��� �ˌ�=9��
2mڀ���n�,:��Yj�i2��SD����-���SY#�F��o*TP��^-]hK$�V�ߙ�MM&�-PԶ��5^НT�]��]�>��d�Lx���E�I�v6jv���GG@2"?9�k!�V�S�c!���{�&�?눾��f������N�|XpvZ�됸��Ro���Z�~N��8a�viv���I���`�9���e����S�\�/�q��i˕�s{g<6��c �����5�b=���,�g��ޟU=#>����s����<�-��M�(�h��|�:1�	A���s'Pm�d=.�S�?7�����qPnD�o�,�6L��r�v��f�Z��IxY{��T*�I�5����"B㽏=G?�} 9��
;0��`�7��ٶ�n���Ǩ�P���+�3��s�U�N�KS��H���9�_VGS���=��P�Vd�Z�[g�����v�V*�9]_�$��7��s�a8Hk� �A��8��y#d�5��l@�O�u�;W��[�]nݼl�K!:yP�����>�����X׏�J�F1x��)�m�/k�Nj?��x�2wlP��W�akm9�U��t�К-�|3Er1E��+-���N�N��g� �䲆��+H�I��PK��i�0�/�Ӂ*3ie^�y�^��i��xq�eM���:���vM%F������*��!.�V�&z]s�vj��-�IffTIu�Q{�ir%Gke3�t�	\�U=����u�t���2��bC:��[#(��s�����ј6���͋�7<�w���H뿬L{}�?#s�����Jk�{l͏#��ƪ� ��r������T�-���ذ��w�&J!g6$������1�_���5�I��K�<r'Ľ��ä���D���c���˽	4lA�<�<�8�<�/��ûG�������[�	�/y��?l���G�cz�`�"�A��{��)vچ`��>�Yن�<�V���B-�@��2����I�����������+�� %"blrN�sW8�w��D��6�]� .g|Q�9AS�PYʥ�����E4��S��X⧠��K �\N�3&�q�6#���_�@o?	���\:	��*����,��p0�ûq�H�k�CUS.r�/)�������!{��A���s�S7.V��+����y���[^To�Y�V��̃XP��e�&��p���[��{&���5��I!Q���,22��M�L+�_A1��x���J���xCU�v���4���޵�q]js<E+8t^�`���E<]_=>D�8F�<~x����m\����`$��<��a�g��s"e�Ѓ�úf!.jgag�,O�[qM�������}?���|{#A4�z�v�zj 3H��W��MӞ�Y��N�9�L�=:�"E���g�h��I���X�d����j!��aI�z	�w���;����4V�y&jB�[�^i�jfTR�\��e#w���Y���Go��G�%��q�v�K�V�����D*�~�K/|�Sг�Q�b9ƳA��K�Ij���S��I��خ��������ߢ6i����������T�� ��_E��RH��pk�T M-�2'��НV����d�t���Hb⨼	��|��~��gc�~O�D����S��0o���1�m����M�;���]�C�$�>F٣��j4:ن�U&�˲�jS�h{�ȍ]� ����K4)!���qq�-Kle>�V�JsŐVKݥUkv���i%� �B��z�c������%�u�0]>���m��tf��b��K�=n[]&d�DN��&-{Sv�ONl�!dk�4�EDB3�%:��0_q�w:�=Y�q�n�O�?���zo�{=�: ���m���3��F`(y�m�'��k����f�EP��l�Fw������o�.�����6���:���n7�)ϒ���ύ�L�h0V��7��;;���Iqm�PTb��ݕ	�L�0XG���i,�>�w���ĄQVE7��5���@n�#��3�G�Ñ��o�J���6o���Z5�~6�m�n�>�iPjA��^�蹠�zo����=��	Y��U��1��S�L�j��-bCI�I�A<�e�M?e��/�F�ZF�+�M�K6w5{sࡁ*�|Yj1�kl����uq���m��c�7r������/��!���~�A�Jo)dI<B_�W<�V~x)�!�̺�7<��:�<� �gF�u����^x�2�)� �s�A�3W�.�a6�Wӻek?�@Q�yK?���R+����/����>L��8�`�4�f1߅�:P�\dfa�w��Z��P��x�`�_'�:z�o��v�Qc�+M��wgd��[� ׳ct�ެ���g�ۨB�{=���颒\�qԤJ.߿{�bK�'����@ �~l�W-��d
�'"��1	,N�"����F���P��֟Wl�4[/h@��K�ik?��]���n�D�!rͧ�>ޘ<�ih�ޢ�#���M��'í��x����j�����ʟ�f�v��8��'��u���n�8	,P?�|G���	��|���iܲ�w��.��s�~ȩ2�=�k�#Y�/�:;-�.�����L�t���^�o5��|�:��zՎm�cUϘ�]"���|D��Փud�&�-�RH�v�����g�8,f�o�g�g�e �����qo���V~+"�ˍ��#.�!�Q����+��7��S�˵�;��*�Q'۠Ńv��3ӫ7��l3�=K�����Ґ2�-Ո�O��e�K�}]�Lu���~��O3E�1 1��:�X{�fL�-Yb����rۓj�Ȳ0=�le6��:4!.���#����=^P@�H�M���'}I�R�1���YD�0׷99��%pZ�5�q���>�.�F��'OGܛ}��1��:��2�#�x�S镐���j@ܯ�}c�Q7�OE�g�j8�BlKׇ���S��jk��|�E'����(���!&��{�E�\��l���j�f9����T�/�n����-�u(d�4����Չu�xۉ�
�E/�aS���K:�d �A�����j#��i�B�әwʊ- �mx(*Q�~=I0�w���W� ���u!�!���m���y� �PfhC�#)��u����K�	z���S�\MF9��7���b՚�)��G�2��E`d�B�٩�Iȼ��Nvg��H_e���GtSloGdJ�p��S@�b ܒG���~3��έ8�������WX�;@�7�2橍���:qwUR�F��Iɠ#����%�+R�H�R�G����vf]W�/�G)g ����6�P3�#|w�ʼ�&�>�(�Ѵ���<>H� �;�������
!S.����sL-�F M�
B��5Y���P��#.j���A��)�֊�\���-�X�������\ˊ�]�3\�ן��E��d���7�U6����Dj����f��/yqK��]���w;��*rfА5k�?5;�5�'u�!���_����~�m4T��}b�n?�r��{��?����<!Y�/9���x,�[,XO��ʪ�]���l��߿@�� �zk!F[Vn�� L m�CWӤ$��
��ny:��|1�i"Z�K��`-�Ԣ�|�;�����P7�8Z���7C�����XN�'�����������U�!��)JL'�*1\�o3���q-$��CN#jΘ5i8�g{_���ъrr�tm�5�ׂū\�{�k��6���)�YE �Ҍ��(n��6��tP`�Ւ�`*he�=�y�boz<�Y
��1a)ޜ,%&��h���[��{|��/�c�>��Rp^s�O\��/��f���s����E���TO�'+c�����i�a�
=��ٻ��	�'���d����aRO�1X|���&��k��で����P�X���r)������t8�XpR88�~N)68!kdl��<�=I�ے�/ǥ�;^�U���k7U���0��|�V����ce�D��/��|ǜ"2�H�/�F��[�	J1�t�g!�J-*TU��H�#��u�~*�xM�s�~p����;��2o���VD/{��ӣ"a<��;�h��=3Q�6��r�s���q��~#�S�.+qS������[Z�)7��C�.��X�R�{"�}��f8���a�|J���ߖ�|��c<�8d�L%pO韵
Ij��8�8Cs��ѧQ��׍ZUd�",��@,�T4!�X�%ծ�v�y�rM�?ڨvl�0��f��S'��'ؿ��A���_;Rs?�i���o
�<�Nw�Jtw�uo�y� �ƫ��W��"�S޾���<�ؼQ�_m\:	 �A��ƅI?(3���q���{��������"ew�m5�T������NͿ	Ti�)h#Aɳl��Yz5��{b/lTng����k�
���lq���뮏�U�C�5A*�)��~Cr�u�wx������yi�"b��2��Z��ڧӼ�,͈�k�v����=���t�s���=��5iP�Z�`�e�S�T3v<Q�aV�
�E�9z�!��4xn
�f���5��#�����!�b}�ꭅ�ն���{�a@i�����{��1�ސrQ���~*5����Y{j�}y�Oy窙wi��B�Zcu�$ˈ��mBG�v����\$��H���8O�앺�̵��:B��,��N$��d��EN�at���u�MRT�K��F�����b@�*O���B�e�@��@l�1�ڏ���RV�xE�"V�����i�?�;����rf��%?�T�C��'�����,%9=�g�\�����eQ����t4����=�@����i�Q��=�n娱s�Ӫ�@�D�}�����7����{�~��e2��`c� g�/����C��u'�Q����Ժ��*Ng�/k=��f1�d�����/G9��.�}�-jmQ�r�:����MFJ=5��i�8�^��vW=����by�������y��|h��l{���Ie�XyS (�9Z/��ӄ��j���pe�;�����z���	�_� A�j�5�c���� q_�EG��R��S���miT�Dat�yOv���;F9�G��z�n���EHp���_?��^o64�e�n"��[�W�u�f�X�=��v�RѰ��"��Hh-�:h�(LUH�zl��Ȓt�Ǩ�޲���?,-غ���k��]��֠WDً�2f������S�:�׳�f1����"a���j�uHE�tM1��Rc�]�ʛ,:�<�ߧS{f��Fq�,#yg���{pı������mtg7�T�?�����6��_�"L̝tv�\n/�pg�\���+�W���J�r��<�򰺜a���a��3D��
{���+��G0��we�;��J�B�+�Q���P�K ��rW�o2<l�EJ��긛�� �f�@��0,=���٘�S�*�D�ʹ,e!�B��0�8�1�`%�"Px;a�ts-�}vmR�G���)cZ�����t�"\�Dn._����f
��� ��E�p�$���]`�R���l.B���g��p��Vn�o�O���%�!��ѓ+�$�u���\�o��1X����4?��4�ed#9�A�R��K��j��� ��K�!��(r`��d�����c@���Z�Sx��f}M3X_���
�����?��<l��;ݗ�P��^0�%���z��3RYR��L�2��yth�>�?C-06�k�ǢRٲ،�.�F����[&(nԱx��"f���E���ȷ�uG�8�p��<� hy)#}c�
(|+п'�  �$����̓{��u�Z��`����J�|)��1���v�Fi��*O�r���j���� �X��[O�-k.Ҵ팳Y/�󝤗��I��3�A
�at܍�~�K�U�%�rȗ��L�h��y�6R]�M�gzew�R�����c4m��H���&/��Pː�S6�T���VB&+��@�6Νv��3s\%w]��|�5��)<��J��[��s83�rb��m��$E �O�;��2�,��G_ғ�,����]��h������83Z����8���K�8��ذn�Z[3yT��h������6٠bQ�[���Ѵ�¬gMz+S:����h�r���b�i?�@��%�5�Nԁ���/0�G�b���z�HVd���������U7|�L�6[F���8�P��~������������>z�P�� t$�ј��|���>&q0�e���kI�}l�/&�Wp��1ha� ���?@2<|��Fl<�CZ
��C!�2��.�]vT�G��O�s��K-M�Ak�\�{PL(�&`�j{I5>aj���j|c�3T���'�����/V	�0u$�*��1T5B!8��sہॊ������b2�e��Z�����!.fP����E)=4K�nj�S%��Lx��Ê��������A�P���W��l���q5��5B��v�߆J0��`�V���p�SQ*v��b���x[���Fd�=0�������!y�l�P���JU��T���^�����ˊՇgt�*om�a�ɦ�z���.A�م��E�LlL�K�- q�;3�^��K���E�냦��i �� (n]U�{�{Bʞㄙ俅�fn�(.�1�R�QЛ��U3���vFX1(����Ȁ�+���)��/ ���	��ꁊѢ�'���f � ^̍���|�ML���U�b�n��G�i�~���	�6���Ѥ�ɷ�
�D28C�g�n� �?G�󻪯����N�P�o �E��RE���ʕ�`(��� g���I��Ds�{Ds��-�z8-�nD���n��D�/����8�s\��ɀ��A�2d�����'�Ϯ�[ˣ�ѻ��F���#�	�� }FN�+�4ߤ_ħ881��Vd����	93ڏ|a�2��ߜ�*9��qmoD�p�S�� ��r*Y�^WK$��:qoNE�t���jKn��pK����2�s�˫��k���w����1�X������H3�sWR��?��?�$�>�̟b!�����������T|�3��B6��=��f|
���MJB`�n�X&�$^	�O��؎ n/M�
L�cf��N%��չg���Z���da�Ȁ���u�����&f���&��z�P�a�Qg;vh��M�I�T��H�8z�q�!\P�E�k����ęab����Ԇ�Ա�D H�VyA+A�wQ>S��qW��t��{�#)����D	ˎR�GĞ@n�t*���0�~�;��Z"�(e�9:�鴷���OyI�d[y��;�q��p��Ɗ���$�*���EJ�r�ɾDT7���]�?��(��?ys�|��N�U�E�b��|�@]E�S8�)����/nI��ME��h�r�0�u��\n��P���L����if�*&e�^5xQ�*�8gn���Fe�ъ�ʻ� ����bc���-�VXÈ�0IA@a_�/��q���5�߯��{��9v��-*���o#�*�X��U���n�޳�5�����q���{�����ŜkLP�����H��Am{�ƅ����3]��V��{������dҏl	2��a״���0&iH��2*S�䩗&G ��Z�eS��w�f�x���p���}@غ
a�|V�%@k0:%^�T��Ʋ_z;E�2Q��ٴn�\���MUo��:CΉ���z�Ǿ�x���u��K�"�a��\s�rt�{�+uex̜�ndР�3��n�s#��?z�S�Q-H�抻6M{~̟�n?�N�Ϯ%J�¼�'�#r���;6ݗ�1N�)���6�?��[�,�t�į�w?�p(�9Mߠ�|�Y u:� ���g���Ļ��(��EM�/��������8�Ɔ�<����%�fx��v/��꬧ �_W-�D�Y)Id��^�?F%�h\#�~G��A��g��3,��;�T(��8r�8E�H�/;a]2'g�f����fo�΢���s1s@^�U�&�,�b�[h�U��@&��#��}y_3+]9�'Ei��\�~ ��߅���`�7��kFaù��Ļ<6�W��2q2[:d�ҝ�]�YK�#d��a}�1v��{bn>�C���(r�{�1�0t�]���z�N�[z c#F��k��`�i##7N�eZI� �^���G
tRB�E[G^���kp�@O��z�u�X|(�7@[3�lˋ�%(w+y�d���ϖ��(���?����55���Pk����/����X�T��(Xn}�*���=S���1d�NdP^��}Z������^��zs��Ѓ�X
�r3��dx���63��R������_���23N��$���#���Ϛ��d�������bB���������h>�Q�Q3��0M�d�[E�V<�6�V�Af����[8ZX��~97%DhN�)�#��!��
wz��bY��.jǈ�{�G_��*1_Vh��U��������ұ�Β�1����#Wp���ے!OxN�
�F�F�5��h
8"����8kx��T��;4H�M@����^pOz��e�nP�����:X���`b����.��y�N�
^�bv>Lz#����C�ߏ������vv�H��e,�uO,�4����M[*q̦�;�ӽU���-�gc�����}�Cv�1�����%I2j�C4���Y�9��r�;�(t	9��h����1>$�̒MN�Q�V3Dw{Y�^w��|�z�>aњBޢ�{��Ì.�0�p@�\g��.��,�OqԊ��t�QA?2��^�X�V���9Y�٣(>�-s� ���O���iIl�m� p�%��>�&�>g��W�ځv�@O<;�-��
)�H^.@�G���j��:��jM`�\w���_�M�1���� {u��)������bY� %��D<�G��'C�z�ʖ�/�Uΰk��
�B_ ����犭��v�0*���sV�s輛��i=
=�M�%�P�����~���g;����d*�]ӡ�7��Ȕ�ig�i	9X�!xsF�������G2;�%��9:[��5�LZ���6��k�Yxa�t]^�p/��
�)o~�X�N�Î��ْCJ"�Oc�EH�.�7�H߫���Ǭ��Z��VG+�� 21kg>���6�c�4��C�7�Ϲ�P9�n|벫k�nJ�n���GX�Ĺ�n �yD�b�}��S%�8g^c
6�cΠ��h9��A����S��'��t����p;H�|.������h�R��;��{3@nb�ؖآ��1���$�i�=A���g�K�,�]�xZ�x-EaҾ�I;�����v�S�]��_�	@�1��WBl۽�&�����6�(�J�7G� �U�>6�+�PJ�����h��<��I�6I��Q�d� �k�w��
����x�R�8��i��	�Pθ�T�!���q��_�ѥq��s�߻�r�HY�� ��d��<���@�E��;�_��֖Jz3V��_q��K�	Q=��B'4ژ��RI����7��ej�h���>@�.+�m�륁�M%?�a.�%[�ΖX:�`V�+YK �ZP׎-��'��ʔ�<�	�T|?5�u��|}�(onj6"a�&'|.�y
�m�J�y��
�(���?[�k�*��.�{Kn.;�,,M��}<���Xi��.��Ğ�� <
�kx�`�d������3�rY��nH�5@�e��j%p�GI)�4pK�1Wt���n���3�Fے�ɝ�.����ϰm�e2p(0�l��Li�\S��u��{�<ЮEo�g}��,
���@?���-�X��xNa�������T�>老!i���Q��O������0��4X2'�T�{��k��0�WX���Mi"�����C��E��p�A��5P�OR���ƨw4}+�c����H
��(�nO"��� ѻY<�O{3�o�LC߾#��|�Q����	�x�\���ݨ�'V�#���*����z�q�.R�ľ��س�7��c�4���%�ڑI{J `B�^4������=����,�9?H+x������.�_��m��&e[��尬=��H��g1`��r�c��H;�s^��I����ҰX���ؾD�K`:�v��U���a��&��w?�#��m�۶�Z��Q��ժ�w2
��՚� 0P�������~b.�`���<�ǡB���dl�9|A��^�u������0�G�E�R'��� Ez��]Hq,&e�+���Cw���`�+�Ũ�|9n��y�q���y�G�b��7�`��������] ���Y�� �뵽Ԥ=e�y�i��a=����T����_�jS[�)��L���3��ͬ�f����݌m�A/�m3cn()q+�4m���r��o-�m�T���!$��!xT	sq_C����\D_:q����t��^�؍IC����^�p[Ya��(��{��ŹX*+6cO�'��x��Y^����G1f��H+0���E�Ϭ�H��4Y"��t�
Gʘ^ml���\��H��9�Y���HT�vMO������뒕D~^J��O�ZH���`@��S� �\�	���A0#A�|=�Mf3�G���X	��
�b{��]A�#Gq�z79��F���c��`��2�z�Z'�*��
����:�uV�8C2�@,�B���]-<8�Vdo�����m8�5^+�!߁���C����࠻���q
ֻw�m�[�O�Ϫ���*��8��P	7�ǆ�<� Hd-ć{	�p��Zgj���`ۅt��M��v�������vx~�h�A�
$�68z�gZՎ����f�#a+%�S��1O�v�C���K�@��Mvǜ��ht��єjR��ʂh+��?�ƴh�E�0�F#)[���{��C�CҶ��I�}����lNس(S6�i$�1�	a����ŉ�W�F�"��g��\)�3�����Y���oߠ�P`Q�?N��X
,?k�Z$��c�����~"qw$��� gg�gn1�0{[��lm|��<J�U��Ϗ�&�t�i��S�O��=׿n��Y9����Vb�X\�Q	�&Ѹ���eM�D���!5�t&��,�-�����I�M���P��&"��]��FZ��!��w3�6�c|>[ۥ�/��G۴�Mq�w�=(�{"��t���͔��^2!5u��v��/;q ���0�d�������6^<�ۿ�ࡵ?���Ԙ��I�����u��Iݜ|�D'Y�� �HsMT��q��u)a�,l �_1"����!%L-�pL�����)���`� ` 6�����$���?ZS�H<�X�Dd��Q����E��mt����|UE7���-jY+hᢉB����v��,^Z��H��ܹ�^��^
�d�a�ܦ�\�Gu@]UU�DQ$/��`9�
��JD�y���'q2
r�a����u�s��U*�n��Y�.�d�����M��&O]PP�jPc��`��T���w�?s]zv_u_]��^՞K8���w>�JYA�[?t�|�漪�D'�ı1���Xo�N,ˇ��v�z9ay'\^�C6rx���ܾ狺o�N�4X6�胖ޢ��������F��=�|���1C0���_m���I�x&αHq�P�V.�65p��%���6��	�d6��'��پ/O��y��h�z����QJQʗ�*#<�0���3�Nh��׷�FG�a�XH]w9\�RUJf;�ӪL��H��+M2/8�����ZnP�ɩq0{x���p�r���gr�{�쀂�j�,��v�k����p_ 0��C�KG�}��kC��C�<)� U�t`WQ���2�U?���8񴘁��� �y�L�@f)gVฟ�8��2�+p�,�.��kAI��*��uY��nrW����������|[��N�9��.i�F	<��JTX�	�h)W\�'2�X�����Ś����ӤW q�f*�ϲ
v�K�CДz9�A����)\l�I����]��\�I���[ى��y�|�ea��p�b߽W#��𴰘��W���ĺ�Dl��^�(83�.mR �-j�;İp�7<���9��Ҳ�����~��(��n�$9�WY��sc�����P%�ȭ�݊
�.��M��xI���<���'����O��*�z�̠��&(P�ӊ���O�����La��2�W� 'W���c�� �������<O9��p���EU>]�6:�6��
�a�\3n���cV�`�)���Sp���XSv��� l^,�7o���T��M��ׁ!��uޕL��s��2�E"��>�IA�yHQ����3�-�~ٿ\X��Ţi�-c��;s_��>�18h��bg�ҁ�6Hja��W5�GF���M,�9�٦,O�0�E��!̆�O�����I�GM������**��Z���m3Q�h�|C~![%��u�^_9 �x
�?�yn�;^3@��o����^<�{��v�X~�)]	�E���)}w4^R���aB��Vt@�%�!&��d"�z��_*��=�6 +�[U�k! �J$�H��6T�ҴlIp�&HAjm��N��a���g�`���Y=�S	T�����
�t�|�B���<�6뙪�f�?�����BO�m~�'��ʎ��}n�}��;t��Y����*7$Rcg�i�Nj��]{�G۰�4�b�<�	:&1G)���:`vo?��wH�oy+�;��C������7Q?~�)�k�O*�ՉB<!M@0�s�G�m��nO4�:/�˱�P;��*�/���?��2-�a�|a?޺���|���xGȼ���f.��oY�����aA�=ĩ��H�}Ⱦ>iyI�l�v�NR�J5�|BDx[/Wb[�:�*���w�|�չ/03^N�������}�^��o����$C�D;�d��x,�Vƥ��&k��>Nߩ�;
����f$Ҏč�K�/*.M���!�B�	���o�0t��/��u,8S8d�-���g9���� y���m6����,<�$oZlǟ]mK5�Yӧ��q��X�M�����9����o5~49
�'S�.L(𛸥�Ԡ��Yۋ��|��O�o���7�H���bp4�*�W1A�����E4b�h<��\B�G�^�'U�d�`@�x$2�#5ֶ����氒[ȹ��;u�h+u��'��!Ǜ���i�/"^���H(��N��b> �
����/� ������Pe�t{<$H��B����pm"r�[N�Y�dîc�� �(klun�O�Y��Ԅ$y����b�.Y�<�!|�z0DA��-�[ٱ��9P��+�7����7�f贃����*�H(a@ݣ�h�����V�h[9��	�jX�!�A�G&P�������$c��Sw�y�b�m��A�6� G��Q�0i�?��ث�T�~<ݧ�;�sU��y�v�������7'�Z� ��wռ���K�1"C�vWa�4]�9�us�,(ę�d�O=rfl��|ʕbt˙u+86beV/�WN�p��p���w�`�7��'��û)%1�j��w�/�~��؄I��^���N�qѼ�����z��I�����u�'��Z8�x�d�����:84� �f*���	p:�1��)�#�+��7dI�e>(�/�f��!+�-C*Ck�)13H5�v��`FR	�\�nH�C��zS��W3�y��c=�b-7��ꚳEg<�R��8�o�b7S����ȧ��!���Rd+���yT�L0W9��i�|��{��H!?N���Ѭ�������XS�b�$��I!,�~�}�7�����iM��)���iݫI��+����s������*�U�z�3غ�y� �et!�U���Tq��a�ꃍ�b���J�U��q��OJM�\�(:(���BnU~���\�I��9V���6�Ok����wwj�I�9A�#�������ho�k��Y7)X
����Z�tT���A�>���
B��^ݬ��0��B�\�Mfoh��N	�sً�@�ح�M#捊�������2{=m�~��F��m�,���d�!�^?�YÆ�b%b���plK[?�@ia���Q���a2$�Kq��Û�~���`ש��qת�����[��/a�D��K%`��Q�UE�G�xC��2��%n|�@��Ky��[J����C���g�����:+b6=��D-����t�OX�E�ɼC�,�҇�6���P�X�*��N��P�/�
�� ���ký!��xR��*�#:kq<Ϝ{����`V/U\��4����B~j�~妔��ݤ���.�s��q`�%u�kJ��b����-@�oc"��/�E9��fș3�1ױ��\�l��_��}��,�ͪ�w,��6��4���]~�[o��w/��J�k68�`!�㸗�Q�R�\`�䲬����0��ֆ�R�IF�/���#�a�_G0p��Q*q�g�*���F�q����-G�Hu�N��Q�LE^�^*`c�L��ʔ���f�����Ϩ�?c�����T���L�D)-�Ĩ���_�6�)�b�_�\L.�ܣWf��	����Y�C���R�K&q��������!w}�e���N 2����4nU�.��j�2��
ϊ���i��՝�~���_��@�Y�^�2j��J�����5�9���a���#/0�%��E�Br�G5�3Y����QW֓��ц4��֐*�!|�v��Ͳa`�����0&��&�[;��]všѧP)|]i�Wdv~Ԙ8�V�,�~�l��.d����^�5��.3cHՙE5T�<~�X�}H���Z�3TK�
K�%�K��E��������}�^��ӽX�t�b���d*|�O�9.��i�+�P�,��Z-�e���2�<� i�-K �*:�Z/�B��<���Q1|�t�P/������Z��y����;�/�=�x�0�2n�=���{¾����2��T$G�!��I{�����1d�y��<ٷH�P�H���S\"BV�-��,l2�Omy�F�����/��%�4S_k���4%ec\���#�n�XzU���	��#A��/��9l�|	��)�-'��� ��hL�~-��Z���!��<.��X��Y�Zb�8ꗮ���<�׸�}����gq�S�u&dk��[�~X�fb�-�(h�g+��N@�4�x>M�*I�/���ւ&�U5QO�D�}yB�CɁ�?w�"m��%(�(�l!sn�B��N��e��9�j�w�.�?���;�bo�~��+cOQ����������f���'k����)�1��.�����9��=����'ˏ���vB�A��/��CU�v�kV������+�4�=,��6��:�ٴ/}�]�V�ؾ
�%�r�*��N�D[�_��u/n���6�X��Y��L�ko6r�
&k�E�Y= ���q9��IT��P��=J�(ӱB�'�:
R<�;�J�蓉Ȕ˿�IHwY���{�?2� ����6ú�<ߴ8��$Y�&L�P�A$a)&���ن6Q�!��`�:>pt�<��|5��1\C��g���#�꺧.��jZ�a���d-ʒ�%j9c�,ל��?K����U�x��A��ҸT�N$�C�F�}|�ph��u�_Ɠ�a�8D��q ����ϝ���Q
�{�Vc�z�b��%%��|�vr��/��L�j���Q�ݮ���b2cE��M�L�t�B�p{�����$mۙ'��~�5LuY�C�{�4��Q5����^�"��n�
 �Շ���$��͞P�,��J+~]Nz��2g��l�9>k�"�;�"���͜J�d���I�`<Pe���@:\=�Iֵ@��ܨ����My��c"SsE���QO+V�X.^�a#�j�+�Wh�������^z[n�;s��1| Lvw�o�����\N�Qa�"�8�?�8�T�I}���YmV)FL���^&��E�fxs��3>�I[Y~�K)m��8��/�o�eU�������71�H �GG`�zYհ�&�tN+`8����d�^+��vJ�{�/o�܄gD#�����k_hA�I���r�~��Qc���*��Ɇ��<��[<� �Smnb$��Ơ��U�촛?5���@��TO�u9���QE�u�Xq�'�s?]AjY��
�R杇��:���5@���:G�Oԛ�{�X������&�b��1�'�v����w��|���k R�@�;V%���w�����
���J}�,�..3�/�x������!��$`�0���f���������۰��x#�T俙j�̣ܴ�:^�ٝs�9ϝ�&O�^�����J��ݓܲ��Do3v� �wL��ٔ�{����-L�\?dBʶ����:6b��V]sW.�蓱�d�<���� /4��}=�X���S��\FV%�'lpu�d��j.�O���2�Pr�>^���`�8���}#����P	'w���u���K��W�y�q��D׵�m�ldT��/���0�A�0qO�e���24�Xƕ�amע���" (���ۧ1x�k�m魈��_�a3Ǻ����x���!�K����/�>�8º�k��Md������C�J ^!4�Ϫ�ȡ�rk�_���'f��"��u/v�Q� ��P���|�}����	�b�W�.��Q�$6+、���R�e��{�P���^LLg�wV����%|R�gᲝ���Txy��_�0M	����^ћ �8/�>����}O�$+8C�o�z��V�+	�B�\pd��\����#�PA*�5J�n�����l.��n�'sU�w�	u#� t������\o���ZDG=v��-ǡKI�K�t���\j�sA$�:[(�_�Y�"��M��HZ�.�z).�����.�x�f1��$���ŋ�G:392`�
҆���`#*g�ڝ��J�bΣ�;f 0���vN��PzV���+9, �k�*�L�����[��$�W�@�:�@~����������];���1���$Hy0C�$��n뗅�K��>V�$�N�d��Q7Jڝ��ח���v�6"��b)�k��
e5Izd�8���PG��e:������}T���\�ϳ�/��UD&ŢU�*�}1��f���)���#��9�FK�1�V�sWgi�P���
`��_C�nFP��� "8*ae3iP\�M���EZ�
�HT&�.�m���&E��y��n��OCmh\O�m
wʔ#T��%i�i���Iv���d�3P
�QP%��m������_!�N0�>;�#�me��V���frOg⼅�����HHX�Ĩ��rO��S���=��*�����+��M�g�JX�hC��1*a^���d،�d+��#��z�+��X\M��NM�� IJ�55f'�xPe��m?x�r!)Lz�R�,3��=#ȋ��z1^#���mj�P9��}��m������K�q}���͘���}�R���d
�D���^՘۲�v���p�l��w*Ţ�e���?�f����]���� �y}rLb�΢0�^�ы�72��*��b�f�A��W$����q#t;->O
&��-�U�u&���u_͌��"��c�[�{�I!�܄���(t�nG���,��g�&T%�'*����r�@������(�HЊ���o<�ȁ2U��K�������p��օ��=����9���R�U�0��}_F\n '�&rfI��m���<_��`���6d�Rֈ|D�T���������Is5��ᴥ�2>g�ێ�{�U),|�M����3��;1t^��D�e
 h�f�wv�vXtB[uн�6���_��J=���[���C\�gM�1����l���T�' ��d�8�LؑW����D�o��9l/ĺGJw9IxI�>kKV�ɫ ��<ڡ��3�r/�4>RPY˶�����<��@J����ܝ�^k;g��޺�;�\�pR�MH�_�Pޗ�pi����,�����>VAZe�-�c�T���NLV=
\}�؟A;���7��4X�cl\�uͰJ5��ȟ�U>M��j�RUj�Y��daac��Y�-�lR��dUF��RE�y��_&�sUv�+�w ?�C���8l�?���z���5x�P��Tc<B@vh9�NL�$��Rͪ�󡋺i�|
Z�k�D�&q7_��o����1n}���U���Ơ��:�_H"��n僼D�tuӎ��\��w�l���
>�Ta��C!3�{�/9j��}ga������_;{�.^��sFbE���U����vGfCƺ�m��&�XSI����&����L*3�/T��`�Qrf�},�ѥ3��8�}}��F��7��
��٣W?�l�*d����hA[^:>�`ߨ֦��,�/t���D���Ɉ�а���6d�e�Ê��x�t|�sd���r��)J�	?r�� ^R�Q�0��pS�v>�'r�.22gW�<z��EOv惊@�4�^gR&�Cnf�Y*��S�~��q��ȳ Rq0�ݘ�5�+��4���p%a/�	�d���q��$XP�Jl��Zd��(�+D�]�Ś���?�^����sw���$jarrhZ_�.�AF�#��N�l��!�9/��?��Ձ�ߛC��^�sS~C;E�Amn�V���]��<TN�r�C[-��.�/繢�eҧ	4��O���r�.�ǣ�3�Fv��B�G��A���W�S��AVe��}�z�D���ƃ0�C�i>Wz��t	pW����V�h~�F�.��u����\�AKfOLh�PK�{L<Z9aD� ���g��.%��a�(�P���=2�CV<��`˘%+�w<�\�qދ���g���F��h�����H��˄���Z�AV/"OE��d�S�\N5����m��_-c���N:���a����.��"�8��jB�v�����(�|����a�ݠ�j3�P��6:����}�O��nAG��r�L:N��D�c����>c��ѡ���=p�(�o������ߑ͛�����9pP�(��T�*l�h�Ξ�WA�y�mF��7�K�8���^@,���c$>b�*�iV�6�N"��6^}�Oҕ���s�j���6]9�GW�4rH��?��(�>X�h*���-����V:\5%�ck4J��&/l®�.���L�d���+������F�İrtM�?����$^��%��<�c���mLz
���>�-���%A$u�Z�تS�'	�G#[y��e��а�ɥ��W?$�xW�_꽐�	(p3�H��HF�0�2�%^�/ j��'9F�Ȑ)���9U���w�/q�32����3�D�	�^�S�v۴ϫ��N�)�mH�7OF��8�f���K��,vm)5��m��t�����x��,ib�=-k��]��^d��I'�G�u�C�R/�a��|Q�I$�
p�5r��I;T� K]*�G�Դt�����$׏�~�IX�p��.%����q^[^��H1� +<��ǲ�%��$��C�SpOW��k����N�	�4K�ci�����S���,����?���?�nK>�f^8�Er���j��dsD{�v�����m���A��GKr1N��!�#���"���?B(�G��1]Dϐ�'�O�JQ(z'�L!�O�,"�4��n*��S}MPa"��v~.�;T�2��]�>���t�H��H� Tǌs��W�|7�-h�5�/v��$��6�~��)���>�:HƁ`�rX+����'��_�4NO�-�K(�v���QC�a(ԕ4��09.8�@qN�`�8���k^�����,�f����m{� �����u�`���Yhϡ̷p�*7_�À�N/Ô�q�Lb�Ϫs
�ƨ�_cy�I�����e?(qc}�]�Fr4�9��E��<�<����.jb�#��J�� �E�� .a��e^E:��|� Pp�K�N�oC;������7�]ǜ����"O�l��L��1�b��K)�9��I�u��-�bb]�c��9Y���ù=�ho.&6ėƈ�Ag�ֵ�ݾi�+|DOP�w�[����퍴�	�Q!{!["�{W.X6DK�2N�Ԕ�`��{�8m�������B����e�l��`�TS��6P�#���	�a<�*C#�I��Q�^N��M�p8"��g�Ibծ�ƅw��i������B&dO�~	����_o�LB��4��ە�t�ӊczx[9^���Y*v|�.n ~Џ �(hoF���$/���sK�[��� ��^p�s!�Wx䠩��o��ȱ�k����:�x)t�C�d�7Q�jR򺺆��ȴ�����vx�	�#���ߣ�k�m)���'��pq�fOA}�?赔-p*mI��F1SK��'à�<5�t���h�q����U����r��,��%�`�R�)Q��ڔrB-g��.�)~_�u-HT���@���>k�u��rU��E�歚�;��������Z�U�ɉ}r����~W�2s�@Vh�o	���~o?�/��ζ�퐦/�TJ��������:�t�z��t�2�n����щoyv�ʊ�O���u��&7~���3��C��8�l��^'�����^U���&���H�n%XJ�R����7Vٹ��+A�L�;�&@e����~ah���b1ًg=`��И����8��\�����r� �Ǩ%ٿbN�z�:'�~��k�2o�R����'��2w�}J�J|�}����Xvr_�y!�0����a���1s�ݲ%L�&�� }��������k)"�ًiޘl�`*e�i�(�֐;O���.�v��/��&ϫ��(' v��zKb�%1�n��2=��t[jg�Hsqd�k<�� c[c�µ%Jz�=6��I��A�)~�|�U��Ϗ0g/l�={����f�"@��x�hCx���������(���+~/���䖓���}aR>j�d]`�
{��Zh3�{'V��.��F�3NοB���သ���Z4Rk�{����ߚ�8u�$+!�c�<��"�'S�y�5�e��"Zy
���i��4�̩�́���|����>�5���.7�_M��bB�fr���3Rhp#}��e'�lr�AOM��W�&
������|�Y��J���Om@ۨC�����|���<:��,�����3,�h�5�~.���9-��Z�����{�C9�����ygg���f�U�u�#+A!r�3P�B&�
�8o3�����@_<�b���tq>h	�8��ѧ�k���r�u��1��\V�
U�� 2�7P�rvcX���1Q�5ub����G(e��TDͽ�L>��<�	ڞe	H̼c�����Q�`��i��Z��{WH�'-��Ŷ;�+�����X�U*󍀲�1�h��E"\e�8�����l��ȷ���E��D%=襀�vC_�ًfWgωJ�:Gj���AJ�&R;�0�C�z��g�:6!���J{�q��6<K.hi�����f����Q�w�T"%i�1+���d�F�:�rG�ّ-��as
��ڊ����&��Jbу�2�X;C�J8���-�f�*L�n5��&|�拱M��1��@XK�>�(�?Z��B��`�ޯA�^/��"�ZQj��wZ���tȰT�@\(A�=��J��Z�.��4��w�C�&�U�J��nڳ���9��mt�,G�a�����_F[�;�f�k�sO��.����5s�,����8�m���Q+ʊ�87i��GCs�k5��E_˓}&#�){O�	���%��}\쌀%�#`�x���S�#�a!cn�\|<H��!01�� .hae��o56Yp$8��;	X�k1�ŧ���Rj�%s�  &O�執����RV6*��'u�����_�u�̭��������1�t�e�!JQX��ƚ4��AOa�vA�o��^5�34�db��d��Ȼ�+��J�7�g)&`�vMm���E�5b�Y�W�� |�Ý�_u�{��;��|׏PCƎ�AvT��v}���QH��Z�?N< Ihބ+'X�i�m�J'Ǳ`<#9���Lh�y)�Є��5�>����:;m}y�˜�����۱���nA�M��;ͻ�������V��3
�6y�}��p��P&�\�ƭ����_�+�,�;O�h���xgp�uԐ<�pV��b�}QƉ�l��j���-s�'�M��^}`�s*Pβv�0�>�@X��(RU�^D�l<_�L�(�-b���m���x
�jҴ���p�3�k�u�;�,O��2��pճ����"r�.Skϐe�^V
H�v�o�b�H�́;+�_��&>p� e�[[��ٯe���=��xӝ0���?�)b�#7�[�C%�K�G���DH]8���$?*L�� ��f�P����d��	+��}zD���$�SݨLА�am�����>v�P�L� 파rį���rB��7���f�	�;5��* �%I/�ލ�R;�UY�{�	A��5ɪ�fխ��x	e�r3#�"X�k��]X׊����}���A ddu��n��P)�����G+���۹�
�7/~N�����j��^#nF�'�o2�[<'���@��yY)#��������{�r!&��L��������O�l��5f Tύ��������=k<*��p��}&!� ���Hi����H��v�Q��L�a`[&���Hn~0*���������H�A�de�~EPie!P��*�=&/q�����D. ��2W�����f��<5���@	��qI.�'�gnL�X9��C�TrcqS���M�R
��%�?�X^�������c~�����m֮�����s�s��r��P�r!�YU�S8��[]�FA����WP��B.nS�T�@��^��.���ӌ��_p~��}uOVK_�OJj��������W��q8�5NO	�����y�FÐ��]hI�E�P�B�f��g�S��=���
��?6E3��Ȋ.D�뒬�$�f �Ehђ)�d ��\��`ج<�BT����QsB����jl垂�J����a��s�ɒ"�}~�윮FK�yұ#�W�;ͭ��+��T��A|�}p?�9pJ�%ɰ�3���+�ү:����ťK��r�3�Z��#^�q��8C�����x�3!�:�}��	h�Kl��2���Lá�L�Q�T�Wi#��,���U�T��j�i��h*��|o��}l���++���������QA�\j�� ����8�����P�	�� L��
��1P/a �c����l�q�uR�����ہI�k�W�.�N-G�^���Xʘ2��X���
�E28a	b��v�>M��j�rO ������m���h�c��3;�Ƥ���g��|f�E�{O������h�B�+yr�(�Ι{���Ț/;�`���b�[`�:l}`�����75�o�I��28�9�E�ؒ�HP���5ȑ�%8��j��f��K���Mr��d�N������{
n{��o���Z/��L���
�k�7�QW�A�|C��]dξp u F�/l3m�|&K��T�\�;8J��l�s*FP#Q�����l+R
��+�H4��bsj�!s�V$U��K��E�������8�e�,����;��S��\(T�7�a�(���Y/j TT<ִ\�qJ��z,�p�ۆ��Z�+%�#Y�l�Mp�st��;C���%���%�l����GRωhLo�B.�t����(���X�M-C���ng6~jū������-��u2j ,���d�Os:f5��e���GӘ1����{U�KH��I����U�E�g�81'H�WW�;R��Bٹ�[`��@�M��"<[�˭;=��}���h>G��Ws�~ɂ�-u	W�&��j��ٓ�ك�gڢ#{�Q"��NhG��ـc��;�5[�U#>�^��P�PH�{�B)�Eϙ��nR��gK
����WA*��ϐ|�ª��]��H��l6t�?��t�6Q��N��#�卧�>|��f}�R(�FD��_�I��y��������.���?Z�Gs�}���aM�������:�N����W�a�O�m��ر�gf�9D;Y4�0�F�98n�)��P�T���^����/̡̇z3�m����L�'�0��B9�3���
+����~w��BQ��g�������jr�%6L�k=��[O#j40������R���{�D�M����B��R>(ڈ�{g�Oi���2���{�v#.7�&���J@�D&`ֳU2�$�Y}4Y�h���I�}d_���8f�z���yV� J�b�%YA7q��M�A��?r?�C�]�8'���s�c��2��dK��­*�r�)ng�Px�Sw]���J�0䖓&��ޔ�ȋ1���1��d������㾫���V�nM�6��C�x�4F*_��X	j���&�։�i��Dz�}�ޱ5.��c��_������դc��`��$��n�EM1��A�@��[p�ي���xh�8j�����#�,��k~)�В}i�w"U�����ܓ�Ȑq���f�7�O�	�W��p�q[�
_��&�;z�/��z��9���$YXh�Ϻr�u����|9�DHT�L�����6��g����Ndͦ�^	E�N\���q�/��[�����0\��ɸE�,�9�U��l�H[��J� ��cG���O}��y�7�6?kL��Z�2%P�P�z9�83S
Y��Ŗ���������vf���j'd�`������2L{t�B��.9f��'Z!�
-}�qj��=����u��=�a�-\��<r�TW�q�U�'w)����P&��߇EO�E�Y�}b���-�V��t��]ᘇ:� r�t�T�v������8pe*�m�����X,��Qy�q�T�� ���������Uqig9�3�L+Ȥ۴�|�x���:��_�U��H��WV{���~2�9��XH�F���.7�zb����b���D�eÇ[_����^#��=�6!0����L�RT�j��?��aj��p<���V�T�Dk�-�Z��0��{lʝ��g
ƊSv���)1�M�oS:�m���0�7UΣ���j�2�pT��օ�5�N<����X$�$%.n8 �`V��4��[0&���� ����\K=�p��w��%@ٕ��m2�������/��;"3�q��A�#�Kxܽō,�4%_�4�&^��� �W���"�j&�!;,-�����΢��{���-ZQ8��`8k��%=�X�]���S����Ht'w0')@�bsv@�]���r�Q9SUo�|�B�.1�6tY�ڜ��VQZ�l(O��* Yh~Y�)0n�A#O��|��e�*(J�����11���Fh��{%�(w�:��ʻ�`y�'w��%�V���b&1�$X�ay	\&c��~V��B҃��/�6%�p��V�A��a˵�d�[��Ȝ
�N;�/I��j/�ũ�$�� r���2���t��:i�(�6�ˬ�r�f��8( ���5°ن���Xpį�p~M,5�x���5�2�����}����&A��*��v3-JZ<�򁡱���;u��Ĳ�� f{"��|E�	�Ȕ�@�u3}�8H�h�8��Sh2w�C-�H^=J;�|�uیRA�	��#̮�3��{��~�ߤ���"[YB���x�ԧ�#ǧ9:$�p=m�O�}N�4,_�������kb��cg'��69� �2c����G���Um�YMl�ӢҚj�8zs&¡��Y	�����+V���&&W��5n1G�ܧ��~������	y�����nj�[�����Iq�a�,߁\U	��}O������f�L�A9��f���������O��+]4m�u��͋xRtG$	�8�����'�8O$�P)��w�/�A�*��g�Ky�������i ���BK�	QJ�B8l�!��2�{�Į���wy��d�� Sޖ3���		dU�MP^�X�x8�UQ˛��%�39zU�;E��v'�,�e���I�6|��~iNW�!	G�˾\��o5,���`�{>�L<���Z���H�:���T7P�z�	��K#~�: �?�g���,�����'W�7w�p�<���t�\Ǥ�ը�9<���	��y
�KA��ugw�RD�ᙧ�La*	����7z;�=3�{��ƣ	�Y��d"��A�ϯK�tн�x69�z���p�+���V6X��T�m)��}V�X2[@3N�7�4��Q��e�-�hG�^<1)M��S!�9>%�T��ˆ �;&�oy��iX5��6��潾��4�k�71�]b�F �ox�֨��!Xm�@?�B�d�_5'���*�'`|l���#��Nx
{\/)^c nu��mN���D��(�����>}(2�����|tc�A�h������_�iy�X��*%��Q��f'0W��Wκ� *p����N���hP�+��^R�^D�؆	�
{��GL4��O�ܚ	jg�1�@Hd��A��8^;x�3��Ă������ �a��"�q�\Y>ZՄ?��-�X+��XՊ���h�"����:�H���XY����5�s��|�S�E�-X8�M�4�Ұ����\T��	IN���~������hW���rF�O<�`]�5��GI�t�V$���ҹv�*=�N��l�^A�щ&R�'�W��8G,��&6�K��N�P{B�qw�Ú����o�0���S���C�h�ލ'�T��a+���R������@�e�Fx���xbxF��+��9�,̄�Db�u輱�ۖ���lgWܜg.l?_����	�k�y�B�Y	ݲ!u;X�Q�Y�B�=�RUU����������Ǐd��#��v�}��B+��7a���ý=h���]��GV�����$
ڇ���B`�-2?�4�f2un#l��ˣ������C�T��<C_���k���˼�=�@U��e�Ώΰ�����t�)�=]��\�R�~�4�$z�J���/���`М��%T>>��>�9VT=LW;��Ge]��%�>�Bp8(�g�(B�,�9a�Z�
/Z���Z���z(i(F��^m����`�yq>T��]3J�O�d��DϜ��&�t�m�ǉH��)�ó �:.���)�A8:rQ�a��l�Y�\n1����y��=�P��|2g7%&�	�z�J�Î�`e]��p���o3)�W:��Q�*�5�yۦ�]�1�������~ۗT��^ z�G!�(��.qJ���U׮!���?|�J����%Q��yM�(�8=*�����Z����s�u�T<��,�c� `C�����R��y��OhMY��͵�W��J��F�S���[��\&��&�ٷ(��^v�A��@�C�,�WCz���(r0IqWi�?�^���,��.��@5��Z���)C*�!I�a#5�"�*� �(��.���"(A�����v��6��?��M-��=�!1���@)�(1k�r/T<���8�F_�X�33&�+�-[����R�:S��aAL���q n�0�;���*��Հ�CL>EE|�m���ds��{�q E�q���X);�9#
	WT#�Ļ��B�	QJq5%�߳<8�v?�/�Ƒjx�
.N�lOidڽ���Z=��	�g?>k������Вݡ!^��&Z�G�V��b��3CB3P��	���,,�$^!��|�ΟO'U�j̳�b�r%2��dq	��-�w�hf���C����64��N�M�G|��1�?m��g�7xqa�*F�o%�r|�J�}�,��������(���� Y�tւ�~�����,F>�-?�����������������g�&a��b�[1;
�c3���\
��#l/�(_.�����������1�h����T��7���B�f����Ji����k ���d��F=-���l
���"���W��Z/C˻$�yp����8�G��?pP� ��N���QV��&q"�DB�_�b� ��ӕ�T��yK��d���l6��n4���5�p�mSf�7�m}m ��V���������DB�i^y����J�06�ʹ 4� +{FZB�#��XaKg�5~�9-,�}�d����H�a��|���K��w %D�wK� �o�G�1<���o>�M?����c�j���#��y�_*�X���l(�͝jrl���u���Z(5�ҳ��Bh^(��;���{Gk#����W�������4}q�E�񨅕�����z<�{�D��Zv���#B�
��M]tvr��!�̟.}��)��@";ftGδ(�h\܎p��
�����7�C�о��_�_rH�F����t�L�J	�˾��ԓ�L E�$�rMW��5�h�A$�߇f.O�:e|6`�D�W@h-Zb.F���j7|�))�B	TDpeb��Y48мC|���~a�����C���#�M�콰�u�ۭ���鉟$��%X��Ib� ��Fȫ�B�zz�~�zd?�2�W��9,�kp�l��o�e?;��߃:*ua�xMT��ŕ�#�{�&7�>x�Eψ& �Q�j9��j��;1�x�w,PE��� ��J`8�Ap�	�k�&�zdVs�r�A�>��kz="i��an��"����u���.��.��S��D@iX���^惝��MQ�>j� ���}Ȯ���o�4.H.��J
0`����ƣ�#>���5�ɠ:]�$
�Rg���'�J/e�o �JQM��Zڀ��z�ѰO�SBn�H��9\���5�����t�P�+pe�tr7{ԃ':yu�?/dK��M�(0J�j�D���&b$a�l���*z���ߘ�Jp�8򙽸�#.b�&�g���ڱ0��;h��c`Ee��GsD���߻'¸��&X.dD�L`V������~���C�n��]Pb.�U�)�"���"�X{w
(G^
�Z`Q`�{�?��P�"sڧ�~{U���

 ��&c*��\o���*�
���ygBד�|.���=ge��\&(I -_|����6�3ՏL17GYp:,{ ^VK��2�� ��GN��A��S�_6jj�`8DR9�/���pU �tۓ;�t�x��d�<��P���y�����s���ȅ��4v��ź��T"�Epj�V�z�%So�
��2b��)�u���G�5&��I���T!=3���A*�f"(��q�A��.�)Z9�&(8�+��,ϭh����1���S�=5�� �ۂe�+k��P�o�7. ����y��45ˮ��D��`��j�j�`@�'�M���T����Nѳ���ZqLL���''�m XX�&�:�nPШ��=Gw��F����(BH��ҧ��t�
ݓJ�F��t�7�Ë�dzʓ��/�?�t�K�߬�:���J%?��b5�)`/�p-)`�s�����5�@�КF���0�ڛ����`򡪲o��!��>࢛���FD���n�&5�����鐻�[B���v6ndVw��a��Ev��ƪ�Hq@����Ĭ����7�o�䯓4�n�W�Xs)z� �G/`.�:�S�-L�؄aj[�PUc!4�İ'�mN��3�h?�:�4��-gˋ�I�x��˅(}��5!��������$G��K�BD�̥���hT��
�6ɜ��I�^�8��yus{����5�̀s]�r��WQ`)���8����Sh��
�~Z�>�A�?��׈4�X����5��$���q.o�:A��y�;�K��<wR��4�L\Ř�p{���G\���`y�������%ʆĠl[�*��&��΍d��&��dͿ$N�I�Z�N���"O����B`�������H��PvC\ ��yQA�op�	��+m�[��),���`��5�N�)��.o❎/:��s)������|�x��C��CK����� �;�l�>�)��}��qѹ�@@�n_J<T�����e��"�/��ǧ��� :d;�Zu�~�laX�F'�>%��'��*Y��Х�`����RI��hc�E2�Z�
.�΀RN]�8��5�lD5�M���{��i�7�tflqGE�
��.�9�����<�7���;�l+�����"�-�'�NI�����ӬO�X~l��X� ���%�_ �0�z9Yk�+rǉ�I�C�����D����/�S �����ET�o3{��K��]�G�L�4�¹�d�p����*=T����zW�^�����Q�
<���s��hE˃�qN�z�	r?pvG,��~�y��[��ZF���6L��`ksJ�y�:=2r����ٍ�s�z�n����e|�>c�]I��4f�f�^��
�-��1˕"K�R�"Ƞ��t�Yﵠ�o)!�x���'�����"�ڊ����ų
RE?J6����v�A�`��E�ê����Ĵuh�љז�v��<����%�ރ^����ߞu��7��0�Z���fR��qꯪ�����!���)�5�����߸�\`L��rN��+u���f/�d�-��+��F�*F����P������a�G�!ʪul#r���V����L*�� �OLU:�@0�;ٓ�IR���U��e�O�l������m_j]�1`�õ��).���w(���Y��s"��1nhrڐdz��g;j�j�K0�Z�i���>�I�����ĺM�F��=�-�.�k�vj��2/��?�@g�iF<�G3Een�g�dy�>���0������1���;���o\��ٟ(���Mq9I��}9W������No��͇C=z�q��	e|�b�!�`6W��::=�M"���5��v�ڇ�S�0�򦴽F�4�0*LUS�\[p:,]pDۼ��e{hHK����V{��J�BÖ����9q�\����<L���S��[}���{��<ud�ߔW�D_Kc��z��`K�"h�Z��2��B�0�1���C"�48����k�����R��츒
c�&y�W�POqja����P��8����i���\[�;i�|��h
8��N�F��1Ȉ<\��i��D�ͯ��}��gY�����j�:rS��(WO_�T�lO+&�s�@ĲCw����Ŋ��L:������}Bk�����鬨o@a��G�<��w�S�#ֿ����G;Q"����o��֭����T;
��"/ymK� �[���~Zю��L�u�����Nza��(����e��y��f�IbUS�_��:�g��"��{`��0̿��&|q=��?G����9N7��!@?��������V�ޭ�V����E �,;�S^��y����NPE���=N\Ri&����Z�W7B�����auD����B��|/�.�+_OF<bT�;n5�`���4�QICT��Q�p���!���r܍TU���wSF�)�Q�����kR��ѕd*��`wݵ�X������IO�/I�F��p��z�����r��h�\�p�W� ����ֈ�6�Uh=�� 3�i��mX��WH��*ګP���=7�v����/�T�X.�t�أ{[��ݱ���3O�`*[W��ZH^~2�0�m�=2T(��<"��H��{����$3�N�aM�|��4�>5/E����sy���O�R��fϝ$YD������-��n�?�<���ER3Z��|���z�Ҟj��J�#���r/&�-z�%_��S����jd�B���m?3Y(�������	9�Ғ73�c=�ޔ��/�Y*�b{j�'��?/��ln_���b�e�����f�4��7�;jb�'�Whmny[�4pPl+3�"|�q�������T��}�A�,�	`��
���z6�q����L�s��{�gKrz�=�Z7���q5,��m���g�p�I�� E;��X���b�x�#�j�����=��s���I�u���L���}�����PZ�\�u"�V%���>�8y0S�v���&�blw|I�_UPX|w'���Ѱ�K��0�ao�o�I����q�#��V����%n��0��E�]b;m����H�{MQag��Ou�ִI��?��5 R�P�����<���k:_6��?�n�Ѓ�Vߴ68ӞF0����ގ�	�O��ΜsL�:O.���D�*M�Y�-�(�e����4>\k��!���|E�u+���r�*\@>Rp��"����`]��דi���8<�ꭩj?���H=���M�F��M��Nj9�w2{2)vo٧$��ȧ�sY+��B��*�{�=�7a:�2h�����Q��4"S�6�C�z�j2l��;u[�<�o/V� �t�8�O2vH�;�w6mU!���,�EDx�"k��W(�#,��S�۸'Z�"Dxx5mwE=���	k�#���SirY��Y��H��t*��] v�� �:�i�����m�H:�N��V�{0i*����0Ĭh������+^���ݲ��g�aR��Q��rP�7ȏ��l��
d2���LF�B%PY�y*B��H}%�%�>�2i*�nc��W�C�	P��T�n��ỔR1B�Cu��P
�i[荃����Kt�jŷ<)�N�E�ɯ1��X�=W�	�K�Z���BƤB��7�t�P3q��Y��|�)����)j#㡩����\S��n�Hk姦P�++�9����fV��=)�
�v�p��A�R6��i-��{�Y�"P�	�9��#U�ǋ읛�j���Y�+~E׭q�&j�.Ҡ���8� �&���.;�A��h��ݕ���o���)����9��t�~24n'�(��,��1�BM��BF<�Ot��w�ظު/:�}�]��ʎ�y�h�R��ї�H�)l�MVt��gi<L����A�����'3i1�2d�9���������xu�b�x��pqB��O���uZ���«�gWV��
�v�cD���z�X5�\ZVolg�DlA4�*XB��飽N��I1�,V���[�-���Q����$\J,��,ld_��-S~���f-M�y�Jw3炎�i~���ǅ%מ�	�E!W���϶O�+��,������{�<n$�v��6�e�� �b�k+%���n��*��{�Vه���k"��nKZxe��	d.��.���Q��u_����h �j{\>�%��8��Z��O�n�K4_APo�BAհ��b_��M(��|�&�<� �~)�:;�����1�7І�,�+C�M�)�-I'�[��`���5��o~�Pa�x��PFi�<�C�^B�XR�������0X�������d<�|�W\���K0�\S-8_�xU|��jsr=�$Q��2�J4v���ڎ��WY��c��
(� ��Z���i�Ynq Q���x��^ �͸\�OQ��]���I:�V}c;U�-ҵ�`�����C�B�v��j���3�~Kol񯲀z_��&��lSFP�zDޙK����莘�K�_*7L�����3� �2��(T�N�[�?�����-9�(��>v�3�&��B(�w������[Cjt]M		l���|x_��_:X��F�p>d�D�;�t�Vjju}D�˨)}�w����5ę�#���~R�@���!��&�o�I��0v�LOD[��w��`j�ҹ��8�0�[����}�0�Nx�v,���UN+���-MC��A}���|9 3˴��Fτ�9'�)���S������eN[�CZIh�>ׄI!()�����I��>D�d[�M����La�C�Pg+�c��U�h�=ZOx\D��������7*��e\
���L8�m>��� %h�J��DKp�G�ԔN� *\���5Y�wg�:���CB�=���ӝj�_����gq���d�t�XaI��_�GD�Y~�f/z{%�Fz���>�W�?�Rr%_�P3�^S�`���I�P�t�U_>��ck�(;��!���?��$����_��sj��Ŀ�*�B]�2��+I�K
��StC՚Wsy���~����݃�r)����X��x� ����g��H�H�rX��3£ ��pf��"�9��tD]�~u�	��1'�9�}�phˎ�q���.�m%��o�p��4i���)HM��+p<�^�)�����K��Nq'N8��c?aPW�b�� ��:R�$@I��L:A�}I�(�$t��/��i�8���y�K9&qH�v�T�٘p%pz���6"/�~`_'A�6�y�/S�sc�`��>�lL�*��N՝�L�WZ%=e)�0s_pCm����=��[��"d��+c�������03���$G���2,'�����Nq�ε��n�R��Du��}����9M]T�)A|k�)�&��@�ݽ^%����卝�_�sb��[���L�w6���l}�r�U<��f�`ȯ:J�@�D[�m�=GF�N�V��s܀|s;�R<�,�F,�*Y-vU�}d�&��O�[���U�-%��)C�{�,G;���-$TǑ�V�+B|���Ml��m<�w�4#�D�޻���.�vCN��{��ug��Y�1xo����L��2��W�[���a\$o��q{� �� �n(\�R�I�Ԛt��O��j�XH�/���ǟFC� �r\�K T�m0+�V�?k'(��%0pU� N	�Hf~��t�bU�*G�Zg�\>�R^}ۖgp4����T�.�D*$dqA]�8�AM*��!ę�����)�i�Y��S�O����k��v@Mpj�>�1�M�?I�G	Ҵ�4rm{��Mr�o�&qq�^���w��)��9�?�ji �l�"��6���V8ޫ+z���6P\B���<���̌�ȵ��Ǉ��i;�(-!�8���Kk��:�ޙ�\�M'%��s/O3���������`X��b�Ѐ��U.�	z��U�C>��i[���}�	S6M��I��b�D�ժ���$s��*h}&��Mb���]C}#FH����AEo�OF�c�����$]T_����{�^�S���m��0V�	wB-?�n�v��/��`lt�\�ɿ��6|';$]�^K���J�-�t�%&�k�M�Z�6}/	�3gN�])$O�+���vÇ >�8�_t�HG�R 꼁�d�yde�h�rP�p�"����㭨|�/->������,��V�~!�Id~��;ܛz�j	�=C�����_�(]��D	Хğ[N����T$�4-�H� �A�C�*c<RƋ=���{�6���o��l8k'���z;F�!��3.T�r�[[�� �&��8�5��	^�FL���$k{���O��<A�N����&�*���O۷C8��>y�_�pM�YF�M����)ո j���o���z
�¢�l�Л���>��P-�C���=H��N۞�����yN�p�����f���-�ծ�O�f' �4�����K^-C)Fw��w���h�Cr����P !:�`S�e!G>��-�����(�zF�J"�?1s�w�E�`�?�*�}#w3�ә����vC6�ʇ��:% _�n�s���؎\��f&*���^�H�Q޺�\��?DG��8�% 9_Ԭ���"b~`q�� �/�>o��gx��\ne6�Hc ����z�m]G��h)�ߌ�q�>�iQw�y�yȅ����L�B�N&�j�>� �>V��IR=0B�l���5=H�7��eo�ȹ�lkȟ�K��KH���z����Oِo���Mc%��b�CvCF�޹:�jW#2��as�U��P{m*J����\֚7r#��EOh(G�8�m+�E���~!���:q�!�ʳ\H?~��=]U���D�/�� �#F��i�OI�2��%t�NӦ_�� ��+yS�?�V̀���>eBiF�<?�q�u���������B:)ؕA"��V��h�׀��gEH�}��o+(
��� ��Z�X.
�����X�js�e�|RB$PŮ��l
A-~��ۥ�vM�	���9tPYUH�T%'��ȨA���"���7���࿤WD�|v�5��T�>w��oc������q�����}׎�q�!fnQ�x�2�Uh?�T���I�n���������`��#���v��!��l Y]�%y<�`ݕm�_��C���7ɇ׷28��9����R�Vq�����W?MM��g���	6P��	c�pB�O<rn��w��-��:���T9�F��p琄~�	��ո�O鋴/K�&3�N ����K�nx��:}���B�^�R}�����).���$h�#L���m�&���x�6�����p�E�(l���&�2<}�ua����eI	�N��lXl���!޸o59��F(݅�bǢz����+we��J^9�����C�B�sU����ȝNx��/����[^Ar��Hې<W1�l��z����E�&����8��1¿���V�J��M��]˯w׽��K�I�r�g�	�����9�]��u�q�p��I�=�� &ʝ�!�0�F]^e�Z��lB��q���*D{�+�@��P�ة�+r�����"��3��)���N�'1$�͇���� ��4*(uΞá%=���ҾW��f���"�\2m5T��W{��=O�p�n�����9�B��31�����C�P�B����D�k��Μ��U��B���CgMQ�T�w��5��B��6�{�LL�.2?7	X��?�W�����|L�_�����S9�+�˜�P��_~��"o��.n�n�@�k�^�Ob�c��N�.�C4'����%��m�|'r�_�w�}��IC�ۘs�,��Ej��:��Q��22����P��3�>���w�w�q�ON��Ji;\�%2����͍��|�hx=O�=ð�6�*\��j�t��@�n� �N*d��er��R��-�g�G���:�ǫj/M�k�D�V?�I��ԍ�T�V���b�&vx����Ŷ���"���P�L�l -U�,l���0��gO[�	ܑP6Z��L,HD]k��X�`uyc��1�]Ն�"�Jt�-	Y�` f��r;�;�!����Π��WD��g�*(P����������\G�Ryl�,�~���3�avK�J�!<�z�a?x��a�\t�PC�!�j�Z�8`%5/3��ux+^�fgTҊz+�T�c���L��j��X]Q
��B<X/�J�c�@��K��5�m@��)j��fbH��9k��[�t��q�j�=9�'Fh�8D���z��)yQѰ��
IPJ1+��-�m���s�p�ٗ $
����t����穛�����>�u̔^�R=��'n����|m�<| �����#�W;~>S����*�C�1�z��xA��E��3:�8��(��ђ����t5=�i���&Ѻ2I�ӄ��`2�%'f�ܪP"G�h�MӁ���pi����|R$l;؁��j��tHM��b�˚�L�뤼]�y<��=%�Z�vp�?����2�U�x*���UJgv��^�}��I�i��}^�v���m
s<�ފ��q��iz>z����J@�?��;���Q�Am@ė�A
����N?2^��@���d��:�e<33��Gm>��	��b}B
�{����ؘ8��=�JJ.�T������_YQTn�;��jB� �]��+b�I+R�U(hs���-�O֕;��Iў��?��^
����8h?�.Pj���=]���L��- 5�T�$��+^��Lo����<��P���C,=���:����0/�&�1�����d�$�]�-M��i6�5�*Op)2�%��*� ʈ ��ܬ�'?�Ʊ��*�;+�H�  ��Lߌ�-z>����Z:6����n_L�K�{��<�
����o*�@�&慂�o9�h*%��qJ��� 6V�	���]>Mg6k��W�,t�nd�DUugN)�M%+�Gį�C���z�����H�G ��m��"��_=�@�8��md�@>e���j{�!DO��'6]�ȕ�9o%�(���|���І��gw��Q�-f�j0Rlw*bޒ6:#��������=ˠ�k��i�{�/�3̚�gx�rk�	�����>�8��OD���9�\W?�'��8fF�ҭ.#u����XfJP�v�f����LK�r.
!�
�ӑ�����+��-�D݊hN������:�y��C�2!x��	�F�j��\Ј�t����A�&�$f�\
vJU�XzZ�ׄrh��(�v����Rj�߀?��C��\��Ԯ��m�krXb-�O0�N���iwQ�H#����X�r�#�G�j7Y��cǄ����M�e�����<ѵ{��"j��=}� ���'�0*Bҍ�@=�&�����K��e��C���p���e���b�������-<	���̛1t8��%d� ���ӷ�",�����I\K�H!�v�uP�3��	}|��"?�7���K�H��Q+�Tr72�� ����9�2.�w���C4�������1%�sa.�wv��G����YT{U
�&��{ÇWŲ��l�z�)m��_�]7�kg@#q>�����4���0����3�P÷h��j�"��$j�QX�$r�,کO�y�SjļĭH�q?������R�>�}��� �k��X:��K ��b�M�����
,i��؄���'QM�/�*HI��*��@U�M�����EZ %a�ֶ�Ř}lj开�%K��<Atf�Ћpx5���챸[`+e��v�I�⳵n�%/K���mE�������\�{���u��}�m���f�$���R��O��G|�k靆k��D��9�Ȕ �`�C���!L<yy�k����g�`=������b��D�zI��iRl���Ib�"=���@��������� hߊejv�کp��������@�����X��7w0q���s�B�G�R�~�C����FәA�����{�Kd��]Z�gp= h�\5wPxw����fեQ�n�!����qDb��΋�.�L�w�n����)��/�
�l!=�U�1����S��3t�����ъ����0O5�xӖ�"��[Lu0z��OSr����wsäQ���@�xh�z���ʈuЌ�fj��*l��d'��:9����f7�i<D��w'��֩�ȕ�\0<��NN��%���	��ĸ���U<O��d�PĿF:�G�w��疽v���&[|��<�%9�U({�+џ��_9�%BVt����V�u�.���Y/|�m�ł�V��=��.�?LRN�i:�o�{���x��5mN�*�<q ���1����r
:+�Y�sJ��N�q�_�47���J���N(i�d��T`Xe������\9T��b�X'�!�Y��9L�!����3R�r9�Q����v��dď�GJG��^�}�~�9׌r��{!����$Guz�iD� ���A��\%a�9�"�	�-/��������a����-�͙�j��1U%����D��
�o V��s�&Rd�:�F|�J��;�+7��  ܏���/�%[@����ǜ3K��V.�d[���-j���7�ݻ�.ꚬ�UГ���_Y�9�V�/�&8 ����ʱ�b���@��3��pmy��w�(,D_k��=;4[��ׅҶV'��Y&���m�*r �a�:]��jv�&~�����0���P7�\�d-<ב�o1�㧝7-5��`9@4�%���r	������:�wّ&Z@4���d�Y��Of&�q�8�<�Ib�h�snq"�{������[d�,��S�ʼt���)�����=U���/������z���og�D<��1���|�~~�hu�-9L3k*H�[%q����E�^�������: !Ő2����r��
\F�E��~�_�:5�5l�,=�.R�H��:$��r�"��'҂b��}Blb�s���%�������o �A@��ﰆ�Y�~}�K�	���"����M�����xFqn�w>�,I��+�2Ou�H�l0��O*��˶��3ϥ��th~�#��}��Yꕫ_f�奠����%nIP9$�js�Y��Qf�H���1d�s��I�:��Ee�?e����F��Sa]��U�@�u܇�H��Z��LP+�w��^|m�_���(b���^ޒ.����R�+kؔbPƍߴ<�h]���>���}	ܗ��7���]?�TF�����m>׺�Q�s��f�!��m�i����ʗ�"J]���ET�w���$�"v��O���C�khG}�Y���S\��Ř��R�u�/Zv�l]���R5T'�۬�Ɇ�F��q����WԒ����"^Q��{������=��=~�]��ab�X�5�E2q�K|��v8uEa��2����U��y �M��/������2�0~� @7��n�Х4���wL\S�f���sn�=�+�����o�P��E����!sX[�X������B�)�vѶ�yd�K?���H��+G�+���C��d������h˞�QW�\���o��و7���|��K�7�p���v�-����.b&_�u~�_�g~�DVG��)��O��5�q�=/&�K�odY`��%[k5�M2�9�G	�i��lr#����o����Y)�����g�T�/q��u&?���𙿴�]��b�H�����oӇ.�X�)ʉ:�g���JI��KR�'�z���j��2[x���\)2��
q7�rc��}.��䜹b치9� #��],�"����)vҶ�(�.4���u��!l\��h�[i�B�Ӧq���(�T~�������Jr��h�7� ���D��t���������յc�U8(w��˕�CU5��y;[��-k�5S2?O��Y��m�3���	}�	�woja�~*��ƚ�ƛ3*�mP���f�c�ls<ְ�U\��t���fz�e Z5����Tg\�R2s߿ԝ�I�E�������Ĉn	4� ���/@ңĽ��W#�\a�55�7іE��͕�Y
d���}��z��w'7�_bI�-���L�Xb����lm�v���ua�]�bUs]+q��ƿh��jpƁm��,;��@b1g[<G9W��ZV��*P`��iC��6�ƛ��^��j T0���`�Xo׻ȫ"���Zd��V��aK)���烊l$�q����x2�4?�L�H�aV]��n����T_0a�,�w�]h��<����N�yא�7A�Iۈ���i�m5����0Ո,p� ;�����#�5p�q0�?'�8,�m�'4�l�F&��������V���Cr��'!�{X�C�"�7�]ꣅt u�CP�����/�B4�7�$;������������Ä�
ˣ�*��99,�$��h��n��ǃǫ�r�b�Wun��%y�6�r<����侔KX��]�ڌ�UŠBſ%W<פٚ���qs�����.w���d����EӦt6�>+�M �*gD��_�� k`qv�K��%>1�A}�����%�/�p��z�D�9�p����c�ޠ�U��`E�� ��#v�|�:�=M"L��7>��p��GL�텺'2ҍ"B3�T�z�����T�Ώ��ڋc�����Nik������o��_|�Y����a��B��LK�ꚣ��Q������܈�ų�(Yv�"/y�{�FX��P�@"�o>:y�H+�~}�#֐�LP(hl�%H8%O(�	 {��=���_|�=_��:��U��; ����1T�ot�N�Կl,ĳ@s�L4�nqM��]�� 7�Z�r`��������{Q�$���T�w"u�pxjs��a�_O�OX�,=������� �����K�hR�ɖ�C�cJ��5�����3�@a�4����~Ӧe��1��h�v�[����]®�b*�nr/Y�d��x���������K������b�$n��������Q߫o�Ռ\�sd�G��|C�7��u֏Jz��' u�
qK���"�HQ�D��\�����OzU��
#]��L�n!6|�L��w���h�EG
F,�;���C��%���?&���%<AB�8֝���e�dl�uZ��9oP�`b�2�ݚ����e��|�� �Q���%�o�#������59��V"0������=
l�ŀ�r4&�cd^�_���:�������9�=���d���뵽�6|O�E����*,�2��zN_�9�g�A� Y���bfK�e�@-�����d�H/C]���U��<���8Q/���c{���=6(q �������;��Q���p��]��/s���H61�+��;���vδ ��Qk���e��Z��J\�=���Í��Rr��={`/I���S�93v�&�=V+A�����dR	���(�|"CX��XY
A��Ϳ�ڂ��TN}���L�L�L���IxE�yN��ۡ�p���i؉f��D�u��mS�bӔ�z��c4�5"�M$�w��sN���5�<g�E���A��d����vx�~�Xe��<�+j'�FW�aR]��j�v��?̡XC%�����7��M$L!�wS�� 	5:��;Xң_���]��`�z���DHj[%�1�y�^����3Z������uo�_���=�=�sZ:�Kc�� ��Z�Q��V�H@zQw�Ӈ}��Pf?�VZ^�b���r7�/;�vq?�`^�.Ե���FJ����⭄o%�D�)8���}/C}w	���H8���-�� Cf6�'�Y�AV�L  �=�@��A`����me$3��1�Z�l;�)
jT��%�k��ϟ#QP5,l���h�p���x�~Ҹ�۾e�婕�)����42D���*Ŝ���ɨO�&-����4]��.8Q�C��ǝT�v�}A���Q^���3�őP�=L؞i:��9���/W�7��=#�U���&�9��n�����\�YE���3� ���s�@S��.H��k�������&�HG���&��B�X֐zȫq��Fp>�O��P���ct�>����BU��xkb��2�����-A��se٨�G4v p��İ�,��L������i�\�Kh�I�m����۶�ȣ��|�5~:���D<p�3�F��b��#��S�&S$|���=,���\�C2n@ɶQ�&��O`�Y�0�'�[:a!&W{�/}�e�+�9?|��m�i�G����3^j37"�9J�TH�Xt[�{�&����DZ8,|�ś�d$��h��Hx�����ad�� c����y}Z`re��Ն�����g��D���խA�a�	a�.���b
ٷl�eS��N<u�����	��<ڙu׫
T���ފ5 ]�Re�}j�,��	m����w��A����
�	~K4OT�J�S��a,ܡ*�Ft���!��|k?������f��y� ��{��O)�7��~=��v���<1�;���})�l�Y��l�J.\D9)6vT��gm�b�}��%j����	��VvPr���S�L(<����+�/��L�,eP��*���|�6?�<��\�(P��g��f졻��y��q/�fƷ&f��{ �O�v�yt��߼+� ���)��yEa~7��D����%�%��2s��mP��l!��S\�6�v��JwL�.�d�Hr�SQ%�B����ڠ���nT-�E�1�P\Ł�c\�;�	�Ow]�,c��U˜�ݿM�9�� �H�<���W�fħi���Ĕ>GM�C�g��(,��"�;6�����-濧'����Ԣ� V���Gܔ�}��+jK]�B`��,�'uk��@@��MA�n�:�12s��h%aď�T�5BD}������*'��{e�@���^�g��Owض�<Zљd|��r2�֊P�v?n2,�5,�2�6��,V�ȉ��O�W�=|�zD�u���c��S�wq�w&���wh˻�U�!�N��C5�Yb���Y�~&���ReV8m��GU�!H�a�y��_�U]�B�����n����a�HE\Q*���q��_�Q�>���6D�3 �3;�D�e�%���!GN����Z�Gg���ǵ�~���$!"��p���Ե�Q%�Fؕ��/�δ�I�F)j������#�vߊ�$��.Y�CȮ��M���*�(t� ��sd��Hs�Yk��o�G�l��[��kX�<s#N�EC�����G�&�J/twXT�s�J*��)|���$��u6ڽUN-����q��)eN9^��,�B9���j7<k'(�YA�j�e���v�_N���ܒ����B.��=�9S���N&L�%aMF�>}R�����ǫM�be?����?e'�����V�a��y��K��Q*듢�g3� ��>�ie<�a�E[~ٟ�#�@�w�q��c�gPΘ�R�_��QZ��ER3N%JG�_�o���s�'t�A8�}�	�r���sC���y��;̄����'u{�|� �����p��HnQ� 伙� �V��+��>bH�D�;����zZD�����3�<�~N�P}	�*W�fS_�a97����(\���G�8)N�ͼ�B>�UD��m���[*�)gd��ס\^�A{�.Y�:&LR���	�'�̆���Q�`��g�q���c{�����r��1&`|�������d�Hv��bw��?TA�:���N�N�i��۵Z�:Pe���'����`'_c&�9W��\T��Z��l�ƛ��O{���^^̈́o�؄�5�ݩ�C �jk6p��
���	�M\�9�g�%$"�n���U'�Wj3�Q�U[��x�D�����:��}����2^�g�0vSOֺ�����w��QW5�<�Vv҄����<蝣E���Nf/�v$� 
@��+]z��?�Y�lS�[�ןm�K��ĠtηRA������o�v,�_-�rms ʩ����I{nQ���ˮҁ块(�wl�`3�Wt@���9e&j��Gh�<iː�(C����W�3-��c�Z'�S�F/�v��+�N��W��)묍�'E��&�X��Րd��L�7Q|��)Z�D9F��fhٻ0����WO6������:����J�o�RZDأy��Z��2g�lv��|Q/X���6�sFiW�#f\�j��4(�h�|�ϮQȠC��,�6�0�(������n��*�U�p�&�f��,nȚ���N��g���徘�z��u.�ې��
\����D�HC�:�>s:�^~K�@��r�#f������A�������q=)���ǐ��n�Pi�#����4��i��`T�4��AQ����VI�{��Bʅ�#-�o���4�2���;�#�S���� }����V�2�
�K��Bۻ��m4Q�ci��"g�z
�>�l�D�l���#�&���40i�3o���*��U/�ƶ���xI�u�=���%ρ/h�Vq��n��Y��Ӥ���	v��`�d����ya��N��</�9�����=
�Y2(�^�,�|FY��vf�L�c���	Q � �Xw�@L�\��s8<k����W�t�At�2^����ꍼ���~+fN�ghy��&8�k�Fv L�}��n�:b���\�}��xf���8fO7��'C�٘u�ڠ��<emC_���M��4?%�~���0I
���?>�:h����#����<!��o��6Q�p�liC�@L )�Uo3.�<�n͟�HÔ�����%���3*.�Z��b��Ӛ���?z�n��nĚT�]x�C<#���N��p�jۭ�JЂω��Bb0vU9B�:�c��Y'5�g���;';�esP^�x0g�.ս���v�8�l��g'�ckd�XC��R�%1-=܇��1�3�Qy�l�Lrgzt���EJ6@iz��wN}�4S���e��B[��n�'���㦜���&y��"l��yW����VT��=,��<��9x�v���5>�ǈ�vv�s��d0ʕLV�=��I�ҿ.�m���v�QG����nk"L)Y�ֱ���i���`T�9if	��i�0<�+[�BիEI�8��;=��Hl�Kj��{m	M�Yv�u���;��mB�<x9��x�6�C��^c�,�}���6���;^R�,�-rބ���'��+���qI�?=�j�F�%`gQ4���t���&���jwrR�^|�@��)����V���d~7S��)oy�q��>Ap⣜Hpx�h�LG,���k�e6�e ���t,u�C]���Zz���3v
oxʔ�0�����RB�؁	��D0MEqj�MR�I�C�������G�����'���#�XW��V� r�&ϙ0�	��1.Ƞ�>���G�_�7K�Cu�/u�@}�_��BxC���U����^���\G����x�<��Q���N�ԧb���Ļ��P��ё����S�It��ı�ni��0�?��΍�����Y&���Q���fDn�������,�SX�[2c/��F�k�%�E�?u  �����dϻ��b��FqϱV�:y���G7E�{�6Mk��Fn��B��s@�CZ���2�n���+�𚖦���vJI��ȥ��)��-E&�2ΗB�h0���T�c�3�ˡ���CϧmY���3�0�\c����N��\}�ʻu�E�309_�v����?.�#F>���h֨i��j�I:y'����Yq�	�]���`�!ū9�3f+uaj��ʼ��Ϣ�,��Wڀ�؟�aFD��c<�m�E��z�J��$�^B��)�i�'����k����q���?�iqR_��"H���5��]������//�ZΥb�!�^�ȽJ���V3�� ˫�8s����N��yX�:յ����_� WW��F|�-�~|XN���U�8��5R<�����m�u�(�!���f�k��2Q��2xVǛE����g�SsVR���J_���z�ԩ�}���2(MF���^7b�$��MizAj����vH�B~A���%�Fn��dʼ�#̺^*��q��΍�s51#�G�u�Q� Ey�=���Żx-�X��`@x���"@v��:��X�,pR��Њ@|J�w@���7�UD�?ڶ#e���=��`��r��}�\/5o�-��6�ڿV<q�`}�?�c������g����%��0F�C�˓xD����!H
���#�����leI�
d���$DKh'c/�z����f;�>N8%Ҟџ�c���� x����O�Y��<p�>\�*~fsL��M�y�#�D���M!K��a�o�1G3�5m.O�e�6o�&黩��wzmc���Q��D*����8����h3�(t�C0��il?�qV���s� 2�3��d��k<�`�fDO����|ߒ4=uY���e�q�"e���3TX?�vh.��p������z�)t
YK�[��3��׻v ��'����1����BE'$�J N/�v�3�B���UMe�������-�b2C� �G�oa�J���J(��r(=���g���k1���/�J�匘4�M��!p�F?���*N~E�iU;7(��o�ε��w�8Ż�U<P�vpJ�GhbL{��t�.�Uz�2�A"���b[�e�"�MD���׷k�4Q^�/z�!�m�@z�2�|���hx���Ǣ/&���b@%���=��6�	юf�Z�r�e�LJgw���hm}j�]|o	�dZ-��Y�R>_I�`��r�ƅtf���a�c<8��&��-�Ji�#]�c��M2�_�G�`!����e6M�s�.�phv�*����<	�=�0C�3R,S��h+S��|�Q�̭�J+�N�VqkfȾSMP����X6�R�%�"����Ƹĵ)�M̷�A��z2�"ϥ����f�7I"�
a��*�]Iy��+\�x4��*��|
Fn��o����}��Jۑ_s�m?Mvf�*�s�΀˴��:%����
��8�(94���
>��%�V�f$��`e��C�8�Yj�;�$0�� �\h��L��<]���޶-�' A+�X�5���U҆Y��X`'VV5���9��{9�"�s�0����D���p�DY9@/gh��;��!� N�/FU(��:�7�D�1��K�M�{7n��d���A5DU�����\���?��ǳҙ1���%���0BL��?:���p���5�o�b�j�x�+���<Y:��h�qc��aĜ��R���̢�����^)Cn8�5Ϲ��t ?ۧ�*1q�AϠ����K�>��z�c����b�qj��GS2�l��82Iy���K����0�����I�C�А>�i� ���ۖ�	��k���A���֟* *F�W5�UU!C^6�4�C�?c�_4y	�6�_Qi����~����ڈ6�q�\���ǈ
�B�SĪԘ��Az��woj
x�@��e7�G{�P&1�`��D��@�ߝ8������x'����tͶ�a�kFO���e	HxNa�.S�,����Gxe��7�ES��̊���	������]�����VO�F�����n+� '0��M�h\<��i�J�~@Β��6��Q�2���@�Ǽ�݂�O�d3��K&-;+��:�	?&L�!��6�<S��i����,K�k��@v�4�?�D����`����7�23���ƿ!C���_��
�ߊP����g���]GCg����}Ǥ�y��d���v�,�XP`$A�\�O
�U��Ͼ�y=
�%���[:��i��9u�G�-�������kP����X�c���Dƿ��󀮣��
�ԑ6ښ/��+�&j��>�Ԓ~S�k��Z&�2鴒J�Mpϔ$���l�zvR�-�|?� �?�9��v�(D�Oi�������/��5�g�u7;��� e�9P&{P!KR��#P�����"y���´��9pZGю&&����!��`c��y�����K����� c����pIowtHJ��:����M+�
�+�G&{z�0⍎����;�*~�ݾ8�k��O����I��4�{��>韯�Od�N0-�4Yo����'� `*=�Iu=�����j�����z�(y�$r�i��2)W�ȓ��n6���i�T�
*���������� "�e|�"��}����cf��Y����Cb��S�A�G	tzs�V�O��%ĠB��׸�p���Ed��Qhq;k��Wa>�g���]���F���r��6W�Z_���	Z��{���� /�����4Q�rn��^d���ᢹ��3V���H���+8�BT�ɏ���1f�.�I��6���1�AJz:�ݐ�2�v�����TS��0����C��*�R�/]��X7�i(G/R3~����"w��z�t���������&�wH	����f���K�M%�6��~�{�d����[ɘ���	[�� Gc���Iv�j������Z���������(��A;���vt�!&��꫞{���[����nGʲỌ�H%P�g��e��z����r^���Lă.t��i����ꙁ��&�����"5t5\�9YaI9�s0�(����yI��?C+����Wl4�R�����WG'�^�r>��YJI�DӘHЩĢ�IWv_���t��pY9��v�ea��b;��@d���<���.]��XZ5�͓�c���k�K�Sz�$ƿ��R&�f�X
b_&��'"�uDD8� \��V�=Ga���X��ѾtKH���A΀j#�����w��>|�U����t�����djv���+��L媤��孚`kya��!a7Z�G+3�|�#2�o��M��O��u�i�/t�/�?�-����͈��֟��@�
�d�v���ˣ�kC�ie���Z�1�9���)jX9vX��:���ģ ��n��o�ғ��}`C����$���=-�Q�B7c���5S�<sH�VÄ�7��Z4{D�Eb>���f��޳Ay{ܓc���F�[��Q_�-P�'_v���Ѷ6�
֣2��8��I�J�?0;�;�~n�r��~�9;�u�_h�dx�8�k�:¤����;\��0C6a�/!���R$qE�Z�;⓱�(2:�F(K�\�]<����!���_\�q�Y��Iϊ��T�s�U�������,�:��'2�;D���^���\�ӏ��Ƀ�L��kmkT,�~��kS��g�R��Pv
BMf8���H/
��H���;K9��'	�)�G��^ij�gg����m��q�p��)�1��uK�%�Lb����v�5T�y�f��6ı��!�_~h�8��<?:?2z�Q���F,�������6�3W�r1�"�6��?6Wu��5�2�(:Q#�s���k���Cďkꭞ�f�*[�j+٦���,�)�jx�K_sO":����|I�W��g��>,�赶��x``�����ņk��!�n��-QV�HB����蠕�������cJ����v������h{1E�o��2�\$�͢/8��r?z�)����w^���ef�0�h��X���+��2N�ԥ[{h�w��8��Sn	�i*[�p`zoPz{x0�`��3MhW?B�5�R/�P��a�9��,��T�2�㚱V}](9Oԡ(�E
����	~��K�i��76n�����1�?�S�c4ɑ�p���ck�З���x�C���m�Ň ku�������,M�^ZGb�̎�U��e�f���pՖ'��LKN۩F^m�W	w�ý�}��6;���׃��� R�7�U�"tXvO41���`t5H6��9}5�>4���4�@l��2U�*@_��Db�D F@ϳ!dM�S�e�%��2LZ}���}'���`/H�T�sH,Qm�Z��z�����R�f�g`�����T�������'�ؔd\�������1�.�YIݽ臜b�NZ��<�[>͌����K�X5��@��p5'6"^p��J<+Ybi<y�3F�����7�14��t�
��F�d�}K���n�7�%�~В�h^�>oEZRA )�!"W�1/��@a�jVʣ�k���z�T�%�F���gOuQ/�{����B@�"��L��ɑ�TO�	�����0��}�xHy^�g)dd�{�2L9a44VM�M�,V���L"�&X4��b-�NY`�T���Q���F�{_
YY��`�j܂T��A�zc�O(�	c{s4���Ȗ���ArH���SC}N���h%��h�b�m"�(A�"/�B����4�|� �$=�K�՜-oU�B�Gk��!|�|�J�l�y���N�(��g1�2x�
��w��ؠ�d�K	��f��l�T�A�'\����"���u%ؠd��s�Q������$��A�V��;e�G�����t+���[QiZt>�f����Sf��r�Q�_�d�<5��0i��lٝ����һ;���3�i)�ʹ]���ѣ��مh�R/mY�1� 7��j>����T)״	�8p�?�A%�YA;yrr�-�	 P���2��������&*����n���jl״��/�[�� O�@�y�)�'�<)޾���M�8s� �Pu���[�K�IUt'����ˆ"��O��d5�PL��A��
el�j�+�#�Q>�5]^� ����4����#�����K�䔲MH�1�FґevE�������1#|}�pemd���>[�g�H��
�S��/r��-�T���s�C�&
�����4<|v��r��������v�=Eŉs�̨��ɕ�ʣq��*Ø�s.D�L�/{�)%�~�D�������,z�`5��©x'5C{a��n��4 �#�x38�K���ݛͦ�8�8Fs݈(u*�@���ԫ�JR��Ar"D���@c����U��r��&yl��spo,>@��F��"{�$�'&��xp4�qf���O��5`��9�F�|�S/�	�|����?���d^{�<�(��Da����"��3FC�>����S]�N�V�1�����b����jl�F�\�S~K_��g�`ҧLYCf������\�G� ���;�K��[��"��"e� �UҰ'��"G!U����U.9	:񲚋�Фv��FSi�B"���o��zk�����K�_m	}}7wP{���)�ɬ8��L��R���#�yl�(Y�Uڏ������a���[C�HÔC@IG��w�ŉ�O8I�LB�M|3G+�$I5��t���g9���)�c"1���ez�6��dO��"L����"X(CL���Ē7����^}���xL43���'?�{Y�����E;��A�)�k~�9��;$��>5��w)Fk����=+i�fc~L���I)��������Ɩx%}�JO�jq��-�".ꪱI�h�6��L.�����&d���qYX��`;#ۚ����T�O�Jڋ��o�Ԧ��Y����/M�����j����	�X?6 �4��1j�2Y�K�����ʸW�cƲ���ґ���.���NU2��'r"q�� h2[��^6$�i�>e�/�z(�f�4<������H���TY'�g/Δ��3�q��W��L,e��h��'��W?�D�zx�����3�:�g���?/�4'������ڢ�*4�"dk=�3�%:�����v�{�������D��u�Y54���<�cސB�e�(�so�Q� ��pI�Y�����dܝYC�+�n	��<;W�����H$P����x�C�g7 �;�A�����)�Q���)b���� 	a�blu�C�3��5[�O�$�u��n���3�ꃮ�it�J�޾fY��]p��4t�r#�+�&=��M�C�W^�T}�W-��9�X��A���,Q�!�[�6�JOl��Z�H%��M}Z�Xԭk��b�ӑ
BnzC�dZx}a�j�J�#��̓m.N?A<O�(�_i��黸�XP���2����7�NN/
�d�.�20�����8�?bQ-	��y#����@:o����/;N���{]x/mUͶ�j.>)��)�FLG�{.#��)I�(.��"5Ȝ�����ݵ��`�l�$6[#�e!T�V4e����j�2	���cw����	���F��7���q�p�H�+΍�}i��j�(���V�a|�(��d���I����|�a������ۃ��:�\�Du*�ː�W<u�0��bv;�`G/�����h������W,8m�Ѱ2E���,��������� ����bߖqB�d@���r��f��#O-ek��,s�����Vs�����c^.L'3�Ďr���"S\`�R�e~�~ Ӷp�����	�b<�i�`8�����m��<�c�6#��8���5@��sB����a�X�,��Ժ��4�e���l���F��I��}��I�ai	��:�9�҇���;�4�W+q��Z&�3A��mZb�"RSTWL/����y���%�������%R:�J���q�|3�œW�*;ϼ�3�P��4�l�B5�y|R&��W~������� S=
��vڲ��?��:��_~)p��'&���(G�s�aoh7a��@�,��*B�<��l�)�����iW���v�F��*c�*Q��/�ª��=�a�@���J ��[�?��:NDy�f���yTcx��S=D���,�#��pO/f�aO�����,g�A��A�K�3�����q`�lM�F�4mA?��G왆��Ӳ��6P;~0mN�|�<Eg��;�(��m\�8�,$�T��v���aJ�d͘�إG=� ���n�HH)"�U1��E��*@�ձ�%�KS5\�f`�z���$oi|�@�j�37E�efk�>�6^ǩPZ�>��TQ/P�	�U5k|���*t'pz#Q�����2V�*���&�����nj[�������+o.9=��gKQgַWJ�A��5�?ҏ�/�>�SGT&��Z:�3�Z6����,�k���#\�_�G� ��4���L������W��