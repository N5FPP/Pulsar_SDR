��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|p�n�Uˎ��|�-��P�W�l�#�nv� 0�΀�<���8ʕ��^��h���v���H� 
�>��,����v#���Vo�g7�fh���b���g���[Nx����+�Ĝg>�(�A=� d�<�؇�;����N˅��鿌�a�&`��_w=0I�����ϥ�?���F��UjM�[�:�W\�w�èR�'�N��m�����-5��~���,��J�W�E�����vXщ�I��j��TQ"����^�V�-^0!�F�Ɲ����)k��Rk�KY�r]���/���t���MˁQxR��b�%��+~�f��T#��>�6@UZ��&=J5_8�� ��F�qa
��~�1��AƐ�}�J�閽^Ui�y!��w ��c�]��nX*t�p��!!h�ݟ]_���)������:ni�L�I���5]U�gw�[��gT�P4��x	P��0T0΃RRi�>�U��e u
/��w�"R�O�h�fq�����j��}��������zA�V��D�Ⱥ���)��҉�V���
�T��dT���S��������%J� D�,�a�Ӯ��F�)�g�$�FP�ij�+q������S�U����nz�JI�ࡘ8MGc)1�z�H����?s��dY�E�������xp��_T�>9&�\i��Yb�Az�2Z��T�Ʊ���qea���u���4��5h�=�o�@�C�껡���\-����-��(�	�X\""�8�=��=H��˃���:�Ok
��E���l���4dbc�	{��?G(���cU8����W��>�������+���'nPH��g�),͜�ڨv�y4���2h���#Bu�1sՉ�3�1�b:�]	G���Zv<<�4�����Bٵ�X�=ޒ���\�)}'�X�ϋ��.k���Kl괩��������}yd����J+d
^�Ժ7�fF�CM��rـ��d^�4�.4��� -�,e��2¥�N_��=a��c�>�f^��('��4���ڡ���rѐam�G��߆�v:��o}Jp�'W���(S�"�$��`��![QC�4�C�!(�l��ې'�$i�W\����$I����i���	���:B�.>"�P�-���,~|�h%
~��FS4����c��h�+_i���z��a�|�	u�5�F�yTj|B#,-a�N�IcJ�?��3|���Iȵ@-'r<i<|0��n�=Z<����b��-I���~�%��[���\0$Ek����]�Z���{��-+ȶ";��?��Q ;n� BC�p�$�;ĵ�A�e��e4��s�ɾ�-����hۢ�Gyz�f%�S�Ts�^*�˸^�V�tB�Y'qx6�C3w����&Wٶ`s
�=Eл.YZ�l���X*�{��lF*�X���j�ʗ�=ǲ�xs��"�g���u�\w؉��
�D��{�X#xg8|XQ�a�a��b�b��-k�MIi�ҋ��v%�OCt/��֩�52۴��XR����!C�H��\�4�> �ʎ )5�\���+��9�ݴ�K��e��� �L"�H��:Q�T�;
</v�1A���?5��Μ6����q0s&F�#K�=�<�^r:Y�ݖ#f�Jd�ѰI� ;���hw�^56^��,�d7�¬g�oi�f�[��������%�~�/�@��p��w��`Dۧ%5�=;��Q%�jf2�|���V`��/�1x�L�qp�h\��K�D�r�_Hj�Ӿ�U��5��9�:�!���k���լ�>\F��IJ�|B�K�o��� ��}�Y=Q��n܄��(��y�d�9�,>,��)*�|%�_W��!p�����LL�
k��7i�1W�sQK����=Fayte�C<w�F�3+$���'���_J�3@
k�M��u��R[5H�����+��'��%�0��6|��3"����x���k�K�����U�KM\��n�;�R�X�U?���{��4�}��Dд���v�$#���+��]���y(4�$z��=���V'���D쨴2�@�9p}�Q�T����E5ͫP�
��{$w��6(9��㺲R�#y&r# *�MUJi��>�u��@C�F�uP���19)�s�ʖyɒ۰*��l���A�ݎ��t|����3O�kK�KYkCi`	s#�����n��ҍl7:�F*{�I���4��	��\j�����i(�м�,�x�L�1I��vN�m��>��oϸ�T�8�œi�ۥS�x�������>0y��saĚBc�/C�#g�[�nȽ�2#	ZFm�w����Y>G|ŀ�oG��S<\�M�|�e/���1��k* �LG���� ,~�����[˧tTyw�"Mx/cC�>� �3
��u�5�`Ҍ�:x3F�,.o�c��c�Ծw����/��c oԩat�5�B'�4.S)$��v���u�	Ӟ�uTYV�t���.�+�Zz�;������<�g-~X�?�o�E"=����ŤYq�,��WFQ[j�9�
���Z(}���t��݅vo��L��լ�J#�s�Ϣ��p:y�?�)TS��f�9���\rp~N+ά���ɆkO�SQ����H`}�}Ql�̱��h{��[���ˢ�)�o�����9�{���'�t��_Y��m���<*���d'Of7l���Լ�I�d|�(Cě�U$�fz��3��|�����MX�lP÷��a����&�
}� #+z������
�v�����d�es����績�$�ٿ �m=����Y��{؞�������ۧ1����rv���WJ�H\1��Hk��4�)��YWJ
NQ�[�͂q�� ��>�U����G����CD�k~e�t���?*�FqX	s��9/00Xn�쐞+ﺞ����L�\ބ�[���e��+qD�� �Z�c���w+������
i��|�Xr�rE�YE��p��q027Aj�2^���X?t�7�+��n���W�Q������SᨅDC2��Q��8�����7*fԤ����qf[��oN�An/��9�n��Wk���l���3�?cho���~��߆���[>��t���O�c��g�. 䤏ǘBX���&IϷ���9�G��:O;vN�	#N�Pa�l�����D��Z��a��~N2��t��o�=4Ж��%4|����BA;�\�G�4����Ov�)��~3c���&������,̃�  ���EE�C�4xs*�^@��8_�]�<𽋅�g	���&/�%ǀj�fC7��字�8hl)�гR窢-���eI����q�k'�8��F�#�l�=�?!����>ԁ�X��&V�S7�&��!��³���R���@"���mHq�}�pՆ!7�����H�(���� �fH��,]f�c�B�vR��Ğ���?m�^u��.��7 ���3�֔L�����~<2���9N�jn�6q�ә�^*����S���N ���~
`6P�{DX|�&�����"7J
2-%:����n>�\/����A=���xe>�Z��q�v�y�v�V��9t� ��b4�y�	_�.��6�����T'^�ڛ����ɸ�u�C�pP���,O��u�}���N� ��
�/�p�|eEʇ_ i�R�o��:_ys��^��Ά4ԧ��;V^L��uB-�������
ۇ��X5$���7�02�no�:qI����$3}�O�6k��3GY��[iCAM����:|����U��F�Z�h���@p�;.E�A5uxr���b#��s+g���S��>Pa%�%�x�.8Τ@^>��S���#��ߧw#��T���xscf�o*P	��$���~[�ʸHoe-Ԍ.�r�.Q�L�� !;�]'� ����Ӫ�B���d��u�̖���ww-6I±�Q��b�ꦌbuS&�)��Z��q�x�xB[ĕ�R�fބK$�4�s��q��pU�~W\+��'��
��ڭE:,���85k{{/�o�@\j鷑��aSί�����a�:����#�GR��2?�̓ ����Mb�F�@������H��} �ź�5F���0�mY#SlK�����Lp���Xɋ���"^o�u�'�&�{��`ZE�))Uߦ�5�M�9+���'�̬�1M��Z�k3bGiH��=[ \�W�Zt�IkU��X���+���\M]r��+g
C:¨ͤ�V�S��M�`ߣ2w4\w\���=�r�k_�^�#�)��#�#�3��� Z4���� q�i�~��,�^T$���jY�`^	�D�M�D�	�	�����w��zb%L��|@����[3��z��;WR��c�K��t���_��6V�"n��hC�K�p��*����B�q�k�Rƒ?���(��p,������W|$�j��,��e�=�oi��u�6���@��̿���`�������l?G�V���3�`�������#^P�ո-b���T6r�`]�?���U���|Ҙe��i-�-au�2���]�O�q@�lW�	�٘��'
;\�:o�R���5�F�p��������Ze�c�t�D���O���<����{陨I�^��L醴}@LT'������N^5/(oD�2�178�l��k�1n}
�=n�__�	��bU����Vԗ����9�K�]L�-��̀�����Qǟ��M�W�;($M��"<dP��H�S�}8{���Q�+��������v��؞fT܋���,y�������������Lҧ�1�Bb�0�0��O��S�Lr���ZkS�ܟLUT��_�8z�n�W\�Ne��٫�'ҍ�L������D!�5z��ç<�c�@q�s���I4����@�Z�)_
��v=�xݜ��mڣD�{�M;m[�Q ��T�m�)�.���*Nea��ʃ����~�o��&nt�rAu�|ˡ�Kn�<�.6��*�*���ѻ~�8�7t��bd!��7��/Ǥ��A#���ε��0]V�ޕ�E0�YXN��q�9VO���H�B�[,Os�:���}�>�W��$�)5���@t�C�i����9���#��yz����~MX����޻�Ὗ�����þFoX|f�Ӌ��.anl��҂���B��.�n��[�V x�:c1�%`-�Q� �KwNn�w�<8{�$o�l�3ᠿ=�����"��>2�����i�ns��,��1�̆��%#G��J��3@wvK;�﯌��Xb�{��K������"�4��^��]��x6���*3,����5�4ЛӪ��KL�Eg;~�h�J|�9C�6y�Tι�4��k{A�\���L��`M��4�!,�}�,b#��@b�h���w䂻F:T�Z�x��,�oUl��_��o��ʷ��� �Gǀ`i(��y�5��8m�!C`�}�A뇕k�0�U��I!�w��8�H��Ie��X���Ōf�.R$}�� ��	�	<�?.bv�Ϧs<ޢ3�
D�S�����Gz�|p�C�G2b9����Ls-��a�7��(��i���'��M���,Û�^�i�U���X˶�+L����i�[��ۃ�_s
�W��M�ݞ9 �yc���n��}��;5�K#��P�n!&(�F䐣�R�|�ۦEKq����c��ԋ�T<t,�HPn�
b l��Ez���`L�b�݊�p�|[���z@!��5��T���ԑ�Fp��� @e�@��G��z[F�T'��^O��+ZH(�I��:��ͅ���h�7uĵ�e��8}�-���E�X/�ǖ�d$��T�@�n7��۴�l p�@���<���	b��ߍ��ٱi90_I�}+cm�3��R�$�gvn+��N��d��o lS��������j*/�ۡ��;�I��T�*&�x$^bn&�?d@��BJ���o�ry!�>W��,F��sC�@�/�F��]�:�5L:�_+ �d�3�fG-H�[��u���^�iG�5-���4�>b��u�S�^24n��?\���6�4С��u	'TM��0��xk�2r[{�!�$܆y�X���/M2T��4����|�ݷ�ԧ��-O��	����G)@��q�X�3�/`��� �	����2f���VY�[�IQ���:��v�U3����H��f;-��(�=�$�݉Vvg�[�3��ǰsZ�.������%��F�X)	�z�0e<�8�(C�/�T�Q	Th�o|_F�m"��E��؍�>R
��;%	s|n?]�V�cC��[�AX/|ȳ�e������Y:���`���ȁ����� ����f�t����e��	Y�q�N6.y�;:�y�Y>�@�c�ʱA5�-�=ृi�d]��S#��둱W��-(]�	?}�)\:ֶ���K�%�ds.NE�gٙ�4"�gM��	�����V[��g0"��fZ��[ b-��N{^v�e�x�A-@׸�TI�PZ�|S~�(%���b�Y��.�������Y����gKȚܟ�GUi<" @X�P�7�C�j>;���w�B�$�`���pG�%�������	VN��kuy*c�S�����b��tm]�;,��F�ӔM�?m��-&�H9��E>��$ڈ��/ƀޑ��1�X]/+bw<��x*���I�s���I���r����L���W�y:e>͸yL-8�u���Q뙜mo��߷����w��gl_����'�[�iuސt��"�9����*�Q�$I��!%�ɀ��� ��\�`�zRLb�)�eܠ�䑖M����!=�>J-�H��8�64$?�����1m7v��)b�0���T�ȝ$W e����-o���tfꂨ�����a��1���^��
L��ykBx�^l�6J Q
�I�zĖH튅=��:w�He�!�$ydAOџ����@X����l�E+��K�Ԯ�h`�߮�f�UH�����k�s��Gn�K�w-=.e�lDs�N�
��]rMA"�Ԍ�y�6(Vڨ�٪s{^��'P��e�2/���mO�;�ɽRb,��6�5Bӹ]�Z�
̱��8�*�5�͚��x����H޾�g`�ck&���=kD6Q��BT]�M��h[�oK�Zv��y������wM�)�9�����\�a�J��=�`�/���d�]�ܰ�;�<Ի������Zt�����&���m�&��S\!%a
���-��tlER�?�@_����2K�4�U���v��&;�'��Ҭ~="SO�E�ߌ��qIi�)���t��,<�7�CY��h�����#��RV%.�Ec^��֬0,��J3�'�6�򨐫2OW	Lwws8������'���1t(5�f�~�6�T��i���~^O�^��[�o{hLJa|��'�!�>�������^ƶ��?(	�L��v��@@w�X&���߸��ϙ"�{V��;�1�@�+��l]^PÝ�)a��W�͌��I��~�g����N�4��A�4/��<�lɓ�r�~�m�P������J�0�3�V&��#"����J���2�ì��o^;�m���⚊w�-Ҽ�D��9az��׊ao��^�k�jE��k!���]��إ�-����"k����!�ZL5��T��uMT9K�T$���bM(/_�!Ϝ:��54T�Ʃ�O%�K�>��r��]��bH_v��N�z���i�R�-'zai��~"�Lu	�).lY?�t����x�����t7���υ��,�!8d� Vq���P-�.�Nz��XO�6�A&^U뤸�Zr��ي��=���(K}�]�Iؤ�B Rw��LWB,�sh�6ov�Nx��SΒ��S���{O��L��5p��z�ǝĮх_�{oGc���WpsLq�&�_���{7�4jr~EAejĩ������{K0�~J����|p;#��#�����)��m�Hd:������Q9yD�Q�F�O�ؠ!�M,�4�lS8^�V.���+K��SuBƗjz�[��eAN�jJjHe.\*m�I2Y���0v�`L��b����SF����M��
ĝ�\����hR$b�j��WΖ������g�z���T� �)�MkJy6NQ�XT��������m6�j�f�hҼ����L����{�[Y~�#��ٝ~E��+�bh�5y��cV���*m���r9��ү�[ ����
,CsP�6G��;3� +�����I�������*�Y�� ?Ʊ}kug	��q�h�����U�x�hQ��J�Z%ujqcdO8��ԇ�p���g�Ǉ ���q�H��f<�[�sX��U��D�ە7ߘ��r?��ϫ�-w��.�i��&�3Iͪ�@}	cਾS��9��\mmU�m���ρ�|����䱨��^�5�G�Q����7�&��Ƥp�J�AIT��0̉Wq�/}�<���4q�T����P~*6N�~Y���k]n����f�����J�6�v�s�c��2W ���ƭk]�+8rߕk��ƾZ�١4��3�g~���t�у��	BE��c�z�b`�M�?غ���`��ޮ���]�q=�L�ImK+��fLm���<r���'Q;� 5�y�Y�Ѣ]����7��!��|llD���]q=;@j��q����?z]{^\���S��ln��-l䕏;/iJ�X�A{}�X\	��уy���y�3bSR�}��������몲�9# 0�(���'�X+��6w�_�^i&A��8��c,ퟨ�!����A����\ي�a�xe��dwR�Q0�Ztӌ��B��u��X7�p���x����~ML�J�	O���Z(�h�L����^�[8>@t�[����f9J|�p}��2�إMe�� ��ޙ���r���}���э��Io3�:C�X�N~� ��<�$K�&�N.Yɢ�!l���`�d�)7Z�yصܶ��r��bܵ	w[8')BA��v�y���R;�?�)��z�ݷ�ĊhXn���93`�Z�c�+ak��a}���[?��*ōk���H�� ��D���9)I��V'�}��~o�h�o��n��2_>������~ o����JW@I�a@9z *�7 �����i}�%�lbkl��#T66U�}D���L��"�X��{�Z��&Ŏ��Y� 0��2��am2�m��Ӵ�������9�����_b�D@'Z�ؔ_���X����	�H������{~}� I�� ˏ�f�n/e�����iښ����ֽZA�)Z��g_j*0�آ�A!u)\����;�!��ڝ
��>��ޓ�Z��%�4r,��X)�J���n�^7��0��Lٲi�Q��jm=.�i���bw
��Y����|���U��w�@�}Q�֦�,�b�M���n�?��'�މ$ �VH��P�O�,�[n�tF	
v��} �x�z��aOny��WH~��*~�IS��I?H��U��Q�M��r�wԧ�w��K��	�2ႜ"� �W�Y�7;��A /bT{�iE��5��e t���7��e�V���VG�Q!6�;����i���]�
ѷ�CH�1[����O����z��W��-����O����5��ab2��x�z�� ���M����%�\�e�^�F�A�=aa7�Zq�Zr��S&h֔v��W��;!��]�����UZǺ���s*:<�`�o�l�4S�I��������;��x�F��Oo������mQN�]}�{�R���� �}����f�)��#�j�K�����Ƨ�$"^��wՖ;�$|����ʂbp��^��F��~U���>i;2v�2;'z���\�\|�L��nf����dBL&�O��;�nFw���A|L��G�H�ø3���Eo�[��hK�<����Ŧ@��v�������s�� ��[a2B�{>����+��S��1(1M��2e��<rv��C�P��Xܰ╽�0�tq��]mc�rz�s)��w��g��j�C�y�������g���p��]���u�0��>@2��!62no�Պ��/Ц�E���4{�u5�����gk���X��_�6�?r��gI4�L��bO�5sZQ���}���=�<:a�r����;������=b���&�!�n�}��<$�.W�͝ �3\����I���#ov��g�v\j[���V0��`lJBڭúw<]N�$%���#l(O��XB~�,����z�����4@&Z��"v�Az�0��X���/�i�Ո4I ���΃���F�D{i���D��Y@>G��U��*u�'Rb�yV�BVPY���͑Y�fL?�{ȮZ�6�LR�͡��5��h)���[˲ю�Զ�,��S�y��Y���Bӥ/$�L�ĖR�v~kr{T"y��%�}�;��e\m���t*�~fX���4F\+9gJ��Ϝ呑w�*�M���6��7ߦC������9W>!�ǩ0:UN����M�|�}�1���2 ',K�����bc<�cPJ�;?�RS�wݲ�,���s�7-{/�dJ�_R��"�d��z_ڔĄd�l,�]�S�pb�,+�]a���Ƶ9��X;���H�tSg�I����X�aB�d���o/�v �Z�!'��j����C�8�+����b��G뮫��m36��!�ĹɂV?olٳ�h�0@�b�u�V���L���G��@4#g.��se@��\�s���
�c��k��R�3An�%�C X��~xd:^6��s��_���	�Ôٓ$ٍ�y?i������8�`a+2fõF���P:��&�;��{U��T?l ���DƼ�Q`1��/~nZa���_�4���.+u-C�L�T�Tw_�Z�>�̦RYʮd�f|�-o��I��� ����*����~��"�TA�6�}������y�'A�&�^��H�c�D*uE�φ�c��6���՞vZI���@X2�߄3BDTa����{`��Er����vF��;|%�J F��!���wDͨ6���ۊَt�)�Z����|��93��Ёx9�<�:4�������!#�[�#ȫ����$΂b4	ᗈ.*�Ŭ�E������cm�C�I/Ǩ6����-����c9�g:.�@��>�"������H��"��V*%%(�8I	B��H�g,RS�g>���X��uc	;��Ǭ�8��Z�2T�x@��/�j��?���[g���c{f;�SK�P�E}d�o�ՙϒҹzU���rhjT܆���ҙ����]�B�?)����6�w�$�����\���EM�q~kM43�]~.}��K��Д�JZ��*�#���:�oBQ�0��dy )�τ64��O��FX��D�~ap<IP��v�6	�~V���À> p��gP& ���a��,;���R��:�Dx�z�;��%�����G�R�����2�r-�"�	����A怓��&b(E_�Xf�+�	��+�F�` �����\�N�i���g{�{+���m�MX�)��`~�b_+GMz�wn-˼\[nhw�).�5�/�����/^�)(י�Z���zy���M��I#��y���g�2k�ɂ�dOXU$I�Ϫ--c�r� B�> �x�t:⋝�=.���E�w1����.��(&�C���t��R�#M��~6�3A�:aW��~����G.v��������o0�o3qg�L=�ҍe��x��+܄��Y�?:��|a2=6�ͯ��T��ҡ'Y';��TxP��-���AOM��!x0�� q�V�HCG�pAKo�W�/���_˝�i�G�ym��I����(?v_Q-$?ιk?�e�{��L��*����#��wYp���y��QI�����is����%�jp��L�I;�͞�2\�@�o��, �ݸ��7�n���v�ρ���TڌF�P��Gl+|�W충mւ�c������S���(��mg�ve�8o��nb�)�E#��GƉ�pZ�,�-(��чK*^05��S�9eI��D�'?v�o\E��`�].������ez58�)}���Lj3���`g�R�mp.$6(`�}�N�e3t|P���-:�HDbӒO�w'�E��)�}e��������~Ad��=�~����8&��Ŷ�*��0�?�'�U���|T0j���|��V�,��]'bS���end�@4��h,�w!/z�Oud8����ݾu��r����W:8�%�#i���T�K��еz٦W��>��c�(V"\�9�hS���n;#v@���H7&V�:�~��s����o�<����{����"FT�����d؏�ӽ-�;�<�5���m&H�^j�w�`na����ĳ��$�h�9�. �`�W�
��9�7Ws8�?��Ű��V_�*�@����d�����6tib����B����Vgx����%5R�/�o��>F�A��a��B��>���
�v{�^-1|���c��F��O~:s[�a�@����lC�K��lC��pwN��҄���EX��#%��RYe�^�N�!J��6
E&��q\&�7#�mx�����Жb�7�'4��Mj���W��˶���'2��K�N�Y�K�X��q�0���-Їu>����[Ʈ{�y�TEu7-�4{�����[��]t�ƀb:���0E5�뼩8¼�m�c:��}q�!>,$B/�}~�ְ���|_��{�O|D��ۓ�:���o�@��<����clx��Z�y�7!g_	K�L-��[�H��e����� F)�Tɧ\\�#2��J�JKwk�%�?sn&�f*�HN��#��e������0E8�:�&ۏ�0��!�R W���6 =�*5\`���K�����آq�Ǡ�-�;)��)��A���90���	���"�O��!I�����;��w��'Ʋ)���bS��%0�]���ze�CXik��ю���D� �ٺ^~y>�OQD�h]w�M��m^�0�~�����}ҫ�@΁[�B��}��}���k�6T-��F�A&�D������@k}�8)<'/��4g��?�T��F�'��UﭧX����U����@���$Qs���	I��u<c.�+bs֗��p}Ƈ�륃p����ԧqw�|g��&u`�/�c3Db�I�R2���4��k�vÝ?�8�9�J��&��L���|�w��!�7P�毹���8B����腙�ZuW���;3�U�=��i[�.ο}/�d��cdT�5�浌� Sk:w�?�H$t�T�4[����U&����z�GO�z��OFA[����
�.>�~y���W�n2;�KT��vn@�g��H��b�R�H_���)�2�sx���J>�R4\���΢64U��L�}���Mf>���b�aeL�wl,�����!�y>���D5��x����wP��T��:,1m�S<1��T-�T�^�4�<��t�]���I�4�-�2<Oݼuu;��QoJ$�@d<`�,ԯ�,<~�xi���@Id#�ڣ��<z��%;=ߕ.i�I�tY-�8��h�T?a��%��Tf+�a;m�5R�#d�5a���u�<�"�o���M?�7]'zD���}��P�L�'��B��f��6Ɉe�~X6ԝ�ϸ�~�EFe^����[6G��LO&j2v=+����˒��=�G?r0��S���f��WkL�x�<ι!;���f{*���3-rO�2�^/�C�:O�L0Վ�WT9t�%��Ќ]� �F�CgW�3�a���L٬�N�ߚ)�-��|����4>#U��q~J�x~#C~�ߚ�	����5�A������l6�=s#8�x�:FLY��?�w�v��Ҳa��*;i�I͋N������M;��Y��ԠG�s[H�j��á� ��[���uQ�2US��3��	���Y	��c0�S�P�'pO�gZ�����~ūp�զ�)��?)Ct:�G���������2�'�Lo�:,�zM���L��{��2�^OH��z�O��\%<)D{��ok�����`+-��:�)��M��s��P�2$��yYc/h�O�w�\���VE��w�ji5ї�l��J�Qo]�|�b��_]���VQm���.V߿��v{4)#����1�}x�B��1'�G�2����8��JG�o�)�ZN��� Ыu���
~K��l�����d^�d^�1&��N����_���r�*�穨bU4�ǃxԣM1�l#�[�[R��ϡ�LM���{�\�7/����Š���Ps���T���D�{9���]x� ��}����1T�}��� |v��uUݽU��z�
�q���(�Ge�Š��Vk�%wZ�)%��>�ȰչƋ��q�5���8�P�eUѣ��G�����C��'�:������j�S���7�)�Ѫ+ХC�|�?��~�دwҮ��"eo�/��xm��i�A��$�P�,�h�a����;
??O���
�:฼���#ΐV
e�߭��.�X*R���O��ش��/{�U�<	������{`���ۺ->Y���-�����7�6X�Q��=�a��ĉ��^I�A��Q��J�>N}q��CL��"_K�#����b�Ns�%˨<R� J����־���E���(,�%�U(����$�̢A�b�3j�_��~���h5E�?���p��kѰ{��C���-@�~e�W�=%6���(~��3�?X_���I��x�7c\/��%��=��qۤk�?������D�3Ó;t*��_Oy�;l6�*��%� O
��7����U��A��lӺ��ڼ$;�>��ߠ�;O�rmHFwh�d_�>3���s�e!N'�_*'�"�wz����@O*�,�]�baH��^$٭X>б��P>�I��ܗe��HZ�L��I�m����������^[����f��C��W+��������s�_22��vB@�I�e�t�0=��=O�w���D$1P�R��o�t�&WNa�C2�2�z�
g,5�p��x� ̡��k��X���c�ha��k_yt�W�"U�f��Av�WH�n��}����J֢�盧���pSg��`�.��P�v]Я譚�U�f���<�?Hc�u�7���)��^*j�:��Ω|��#y|���=r��M�i�Q����R4�?)է�b	�	�g��ؗ�g��8�M�b��W��͜]��'�p��IW���jL g�3ڨ���R����RNS{9���X;�u���n��R�쪙�����k��=�%��f*8w�,�<����;��c���=y{P��� Mv0k�E)h���/�X�:.lb�x}t�@UIC@�7,l$5i�,_4�c,v`(���MD�L5��@E�f�X�j ��J7�=���"�B���	��>���!�<��[Q׃�%�j<�i����X�2Ċ��tT���*t�Wch��Y���ߞ�L���^�jTh���+d���]'�+>-G԰$���쇯q�N�Q֦'2�������8<�J��HMk�2�x��I��0�.�Y-�{�sY�e���WN;Qb:P��"�2�~��q�P�;{ �ܖ�F�4V��"ƞ���/�:�i��}�W�u�ю ����/�S�+��U�S�X���9tz5L���"崻������s/B���bJ��� 9�����c;@��)�J��3d!�������{��v��=j7�]�3��z��	+o�\j��dt��>5i^� ��9y���U�3
o��kڅh�o3�<�M�{!��N��-��!���l�'��0ghF潴Z��4��L��_*���.|��kD��~c̳Y�ӽ�����\]�������/���+]hx2��ӡ(�A�<�wɜd\�~�cx���i���SP��9װ������)��U�CK��Φر|�����p/�JN����y��I�C�ZI�܂��uӷ3�]b'�զuq��*m� ^Slt$%Y	h���7�8�.��:�}�8��k��QH�{N8G-���ܫ�m��Ȍ��Cw��}zp��� RZ��Y��p�\�P(r&pg%^�e�:�'�0�$�_ǒ�����{w�vcd�˚$yFh/�ͦ�<�-��ƿ��v�z�,��f�Uݸ��x-۰�Q+���@�k`á,`-�{q����Hg�c"*L�g��[�;��N���Y�h��G(����,J��<9פ����'~�w��	ˍ����� g����,rH&Q�%6��
�����ѽ�@���ty@�St�������{��G�C���H��2���s��\��������75��LUbd���g�Mӻ����;�_p�U��f��~�9ga�N�����Pgnw�}��!!Ak�Pމ��/�Z�/FS'4��
&-˘�ie9�u�=�Hsr�4d�/��X:��@!���% ����g�4��2-�-�
�_ȹFߣ�Y�>w���V6����.��g����+{�
Jl>�����m���`���;| /N�*���-�y�<Np�Uy҉�@�m)��&�Wf;�?�q]6Qq��S��b���q��I/�*�IUն�x�V����I�/�T���6�۸�c�3�8G������y15M���8��~CUZr��9�iM�|�t��©06�U�ߐi���0�F��,�����߁1�����lWxc��u��vb@��˂�ݷ^���̽�!�R���L����~��eAr��G��9��Ϸ�;0:�=#�o�&��=� \�	�y,��-���`���Z}��v�0�[@`�ၴ�:��J�sBv��� �7�
H��sJ���>�C��� m[կ��;ئ��d�,�^�>�",l'�S�n�/�I��щ0	!!���H����+%ã���/h���VYj�Py�{A�l及Ʉ��z�j�|7"�u3'|�t�A'z���'�
7@̭*!���%��˼�ÞK&2|(v�b���C���+b�|6��ٝ�̴c~B��2�I��W2D�ґ�����h>z�J����~{�j�G��G�+�Q+�����_� s�I��[�Ug�f�U<ˆ@��6ԯf����-_��<=ns(b�Y�����:�&��!=�m1�����0��"�L$b(;�3��ih��2��3܌��������v ���GVꕎ�#��(�!XM���j7�Z6sM�ӇQ�l7y˻�kƥ���q�$X��#3\"���Fn'RԵ�)��S�WI�� w� �$8�a���|LS���=3̍+�I)f�OϿ��"	�ӭ�ϵ����D�����]B*{m�3�|��*=P��}�x��һo�[������[�-Ѷy����m�7��v��-?�~L^�K�J���*���ښq�Q�nD�W�b��<,��c�3P��z�-��c�aS4�](���4ǒ�<�Hl�f9û��j�U`�1S=*�ݴ��ܝ�EyZ#��ư��n�3g_��3�1�m��W�ani´�,��ݕ�ՠ��2�OvZCY����:����2m89X�,�f���@k�����i�2�p�r�S^� tLIhe!�4v85��#2|r-����3��L?�@#�FW� ��u6q~�a1�b�Ρ�:�E:��,�nQ�R�a?�>Bh	�&��m��s ��BriP��躾��;_~i�]�湞f���;z�i�^�LO��j ����\J���C�K�;ߚ����(�Ig���ũNNY}�J�Ф��;_�o��z��a��΂<�ri���d�ʰC�|�!G��5������X��Y<�����֡���Tdcg���(gmgߠ�#
Q�7t&guA�l�X�$J<H�hA�X�uvh�0���$��%�&��kũ���l�[�M��-[�l������������y\d��Y80�C�W�y(mݨΥ�M;�;f=Rv*Dȁ���'D�+�*R�N_�J�¥2�^p\�8���ʹ(A�Aa�X��BJ���koa
͠. �k�X 1�%]���V�ߑ�&Ҏ����������%i>w �[�ph�m=|
5"�I�+�ĕ<T�λ�'�T�T��!1�!3��,#D�v������/�ql�ziY�v��K|���_}��P$�p,��o��`+������{���x��j\.�)[+̟�Թ�|C��	$j���HZ�WXT��B�{i��~�ŕ�����5��~�Z�iĸ�����:
ۙ^�B�%��8Uk�Q4�d��:��OO�'=��f�����*�k ���۵���&�2ߡ�����Ja&��p���t���b��F�(W��U��W��-����TO�)` ���Pa1�]
0�?VͽZ��w仼*_�1
$<���l|I������T�P��	�(���,}�#�����H�h{Q�΍$c���ar�i�+K�G���Ki��L���A��30 �I�}����aDk�S /�Dg_��5+�,lf����Z����1ƽNc^�bf���P\ET��k,"�R��sY�#�^By���&��
����:�9G��ڜl<�5���W²����xH�G��9�ru�EqL���V�*:��͐8y��[jԴ�����6A���5L�k�RT� �n�L�d�����I�3����'.�.<�$�+3d��͊����q>�^7�40�{�&�C��= q?�vq���WHَ��w'�om�s�����=[B��cs�A�x���_o#��X��!�����&Ɏ{.��!�Yz���ЏW����|Kl^M����P�h{�<��7X>�
��ï�K)m�H�1���i�E����D�MUf��Ġ��W�Ê��Z�� <��r��M�,F� �o���ᐽܛ�2��BjL��u�\��Վ�^�y]���:�K�X�o9VE������B���N&\�����m�`�Ԅ�3a�j��瑥��h� Y:�}ȭU��k�U�j�pUwqH��0�B��(���C��Q.%�R���3�����B�� {'�'��sh����J���o�8��i�*�r=~��j2$���^�Q���T�JK�����Py�|D�+���36ΫC�kMe�ٺx��S�qg�|��������)�|�pe=JH�L�fA��O�W�BSl�㪐��r*�#��8"q`.��O!�H��
>��3Ϭ�(T4=��p��<�*}a�)7c��U�Ɨ�bG��9����X���K�p[l#����^��3�'���bvȍ]����B�:�}x�q�btY�pe��3����N֌F=ii��r\��>�.>:�3�}�ò�H4�-h���ȘɌ9�D���5�Z��J�Ֆ�{2�38��3�V2�~��]���n�x8_��9�!���9S���q:�l:H�筓"�_.;�]ѓ��U��@$���"�	�@� �(�p�ѧPH��t��U).P��>�Gf�Q�p�K�.��d���R��áw�����#\�����dO�rK�\�H�j��J�M�%�?`9�@�j^/`hE�e��Q9A��6V3H�޹�R�m��L�������ɮ�-u9�����PP�:I�J��/0Ğm5רm��#Ǚ�O[����=�5'��c��F0���y��Ɔi<F�-~x�
�="E��a�*R<0�#ş���c��\�,�e��I���/z8��k��.1�o��zoA�rC�e�N�|H|�p�4s=�Ȅf�?����fJ/xI�LW�2��M�|ꝏnz5�J��]���[;��o�b}%�4��57V�(Z�,�V&�����L4e�S���'4ё�_D��i�Od�w�˾��O����9tG���:�����Mj���k�k�e;K�[�B�q2]��������Fq�m����ᵅ����i�$L�bD�%������Z�%Xț'GM�AR2�%QgJG�$�(��ʹ_>�yBr �E�� �,�Y���b�����A[ �2�9�q�j�KVN`��-��h����Y�.	��J-m�����L.��`\���bc�熾rwM'���|c%�\�$��1v��5��'Zpqֿ�ר`��L@^B�!���5�����X�"��
���%��=HBV7�t��T���զ���0W"�K�o;�@�q��7��W�V�����*����2�F��T���}��4��3����M^#��k�o#ܿ1�\kn�a�
�ȱ��@3~��B�jsgGy�٬3�xy��t#��L��s�[�����pS�� V�'p�x���A׻�2S���0O82���A)��U��m���%z[vxM�i���N��].i~�d�����n*����}���+� jk��D9&�;G#x��%i��d	OQf'��Ɵw�9�=+�Rxx.;~޳m���Eo�k~�^�7�����|>��[je;P��J��|ca�2��la��^Ay��2:��N�֠wx��J��u�Si��c�m�#-{��)#��k%����E�W�����)0����/�7M^@#�!Ǿ�� !����H[���aRb��`o2[{�p;D��=����ii"E�p�$�r	#L��%�ǰ|=�V�f�.��m��P��Lh��@{E'r&r(Z���7)�
Pǁvɯ��xr�e��ZeX,� ��<�0#���Xr5�5�u2@�:�zR%[��>����`Y����_�pD�r��mP����g����`ҿ��ܰ���*N�$�X#*RU}���g��?:�0
������X]��j��n����hU��QUS���ܡ?��!w� �=<��æV����Wvq�*cW�X|���Le� �����q� [���OE����?������`���"�b���%֏E\L5���`7�},$/���|Ӫ?�	 �jȪ_������j����:=fd���S��gNX^�Қ��22�f�$_؎�<|c��ym�M'�3T�+�E��̩�w��n�H[�y2���������7W#��&���P�O�LGm�� �ƾǏ<��<D�`� #
5,��e��Ewzo�@��,P��m��f�}i�7§#^?������b��:���=7���{��(�B��
C,_�� 37����7gS-B�ށO��͹�"j�&" �6(z����X5��Wl�+���?�5�t�L �V>U�e�������P,�QB�KJ�c%#�כTƻ�������nU�<x>�PA'6U B%^1���P�@ڷ���+���z)��0�Ԍ�6(�*4ҭ��'kVۢ�p����;��M���A�g#M��^�Ҫ�Jq�R��:i���x��h�������r���WA ��3V�@d�V,�$��f����ꞭgPl�I�����ǎm�=k�g���oZ{�R���tO٦���As'M&��� �����ݺB��5�S�	�Z!Jdm�P�WJ���;V��|�׀������ϼ¬�Dҵ�9�L$Gb�L�u��U��]������GR�j��0o��X��r��-s��W)�R:|�8Ҝ4;q�co��NBLK�'v�ۚMnZ,T���-�a	�;�f#MN#2�J��O��b��E��pv� ��[�Ի�&պ"M(iE�}����k"���ska�G-��h-���SH_
�����1��*ͥ��DY#��S��*q�B%�<�ꯆ�&��E`F&�BL��L�~��1Kt�+̎&��%&O;;$�L{���q��9�-d/I>�!����]̦�P�^��,���LmY�lD8�	$%ې����]�"t�r�;�C}[;փA���*���c�ȗ��V;�Xa���?Ѷ�RL��-ÃJaf}�����������G�i��2}�Y@��o+�����w3�Z~QЁJ��f�ډW�����F1B���cP`AM����������%�u��;�+?{�3����מ,(���?���/%v�ݸ�x��p����Un��89�zO!��8�A��1��)���	3&/5=�}l-U��*��T��׼'Z�V�U\���
!�a��D��!ÎKgp�aV���;[e�M+�����[����,��17��,��C�e2o÷@͆­���m���Y����(��5����>��ڮS0�!Į)")��$�N`h�oX� ��ܤ��'�$n�	�8� ���-�T�u��(zܑ"�-Y���?�1x��e+2�C��5�Q@����Ryx�x5��Y�_*)��#�*��!���Y�=�(-��ǁ�l؁�-k�_~��>�<h;����W�*^�"eX��٤��Q^Nm�����(Y���R�|�y�=���Q��&J����
 жT�n�d3I�a�ih�1Y�V��1 I�v靕w���jz*1�qF7�\8�e�H��"d6�LT>W*�E�[����v����6�/͉����V�1��O��GFzg����� ��<��:j������ڃ
���r�/vmqh���3���m���f���\���'��k)ԉ��ԃ�JAo�����#LE������2h0�6�iC�w �jt,@�D�y]��66�����c�-��Ag1�<��������m*~M|P����9,5G/��+�`r�d��Y��O�Kh �� lrM<$b���%��^ќ��#��k�Z��5�[� B`����!��{�m�Fw
��~�"�V�R8���i ��)z?`A+3�42��\,ԫ���sPc�A����|��;���Z��d�ڇ��t׋���@��O����_ںo�R�-�$�8�Pr�H��s��{p�	A�z�����|)�ŀ]'��bJ>�>��t��Z �W��p��˫*64����.�Uy�W�W�Wz���>e�Ȼ�YV �
$�*�P-�[�ǟU@��5;V=2�ƶ�N@�	�G�9߭��8�!���݃������˫Cy�w�,8���mK��׉l�����ք1�E|6F�sPz�M��4䮷�m��l��u8��7TS\X�X������)��c�~_R/�����Q-��V@��C���0H�k����Ti�a�Q9�=`i$Z�h?G�wj�)4���l{��\��br���(����q�������ra��]9Q�Onq7� -n�[��	D�)Л�j�(ޥI����/�[����5��M3&��\<��z��^y��d+�|��fT���
�ǷK^���4�{�(�)����z��p�T.A����&��B�Tj�/�?�W���u�ҡ�Ǫ�c��Ã�����6�����0�N &b�1�~[�f=�KH-�G�<�����=Q|����'=U�:n5z��&݋�����F.%5H��m��Oa�,@�^,��bRFk\�S�ng���uI�,9�.���=�aHJ4pq���AX%0������vz �r<�[Uq��٣-�|2TC� M����D7-�&�"��c귰��7>dG�n��ᣜ�z����uOqt���?���ܲb�g�����B�W���G�������G4��\�B�E|߭fA�.��s