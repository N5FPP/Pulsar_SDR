��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY����ﻅЊ���v�-��5���Hb��$Cp���j$w�AN�ΉQ������.�m� bn�X��'�Tq(�<��3�%�E�C]6�Ü�@� v4��$��n�F�0�B(�y'0�'�0z� U�zXe1�: �횅w,�ܷ�F�U�s�AT`��?�[`,�;��R�=���yI�D-êLP�E�/K5^9�.v�eu��	��®�	KV���)�y���(Psζ��U̝2�.�� Nu%	*�e�"��,��`3��6/�4j�]�Xs�%e�P�.�I�ݵ���uE5��GPd�S�+ӑ4�R%$�jD-X����R��8�p{��kMӗ5z��6q�a�م�c��i�=a�WXep�o�q�49[�s�}Od��8U_feN~���y�#�~fEZgf>սާ��R���[�V��p�ox������)���!>������W�`�������coD�er3f�bv�?E�?=��ӯ�=Kh &y�b皨�h�9~Ue�J"q�	�ҏl�\A�qԻ�L�'�I����'��Qʣ��x�ϵ4HLh���*��0Z��x1m�"r�{�	G�A,Qa��&�u.��p���@�c��A�?�Rjy����{�EH��%d�v�ZI�UɊ�RxN��r�h2�X��L���}�$�n��l�D<�BA�d��%UZ�~��$~=�j��1Rl��\��l`��L�ڷ$�,��%M��kFV��������Y��=��o�r{��C<���!�(u�.�3�;,�vh�(CDi1Ed���&��u
G#����(:��-���:���p�ߛ�������OǦ�@%���`Q'%�`������J"�+~�DH;��ɰ�Ƌ��/Wg��MD/B�kP:o!o}��ܙ��6�96�������*���@�LNhŚ%Ƃ֤�hQ����J/0�^�N��X��;	��W�bz-p3f�	�ʁu˪E�e���W揜N�]�OhFmQ�7~m�ʻ>#T������@u�F��w�����)hÓ�^���b�8��E,PY��J�|��[�k��`�R�ù�ӵg�����*�N����-�0�R-�śv����!D=ro�S�>۬]N2%J���Fj�-.�Q)��\+�>{!c�|*��t�)��:2�MW=�ҿ�hE�rTLn��z�b�=�AVZ�c/6�w�����@�M���
=R�rm?$*7�,eU�� �cN�!}��4�[u�;s�iz&��2�
C:�6��Izt����E�tba
:�g��J�"Bw�J�BE��!�"c-!O��&��'!t�M@I����F�q����Q�y$=U;�d�7yrS�N���B!�n��sW\Pe��Iy�c�?���.m�bݔ�C4�, �����T��5+l��%�G%���0M�:�
3Ω�2�[�vι�5�r�����j��praV!���(6�����˝�+�"g���/ިYO:�yi��UB�7�L�edlm�#��/�㖮�h0��ь�9h~�����.m��hĥ�@�U��:3<w����92���0_鍑P�r3t����ء{��N���h�9S��n� ���+����X'Y��rr1��7�Ę�c�������-l,�#����u��/��Z��'VW2�����V��,�~���M��F��+��N0vĊ��룾80�O�\��u�}H������Y�%�b�8ƣۅ8(*��<�_�E�e���Z�:p��3�ճu�/���3���y��Q���qb�m������Nb	���(et���Ap�!=%5Z��y	t�}���?Ko�1���b�a�i�FX����0���j:��oq��0S�r���߭�Gkp3��L-7w�H�~T�n��0cc���a��+7{�I���T>G�4̦+�@M�#'Z�7d�XM��vG�x�����X��5��.,{ ��x�<p�]'=�t�k�8�C�dk��R�h�Ɯ��鉊�5��m�3\�\~�%�����)>�dE�}��~Z�ȥ.�c��3�#Y]�|���Y����D&n�e��:�0/V���o��)7�*�&pYN�Wi���}��\��%�
 ���W�~�k�"��xv)8�&5�f�6um�����9jY>����`�������֒۷A d7�j8��2������ o�]�SkH���A�x�j�<9�ձ��T�X�Lrj��85���S(˻�G�5��� Vn��¹C�s�A�g
�.�v�D�_e:�cj�t���	�T�0�<f�@O�X�N��Ly6/9+!ڈQW,����&^00n�8FD�+��5��t��!^s��֘'��"������y!�6�+1����z��^�u(��ҕ���B&c
��?�^�|��a���I��hEͤ���k)R���^=O9�S���q?'�V^޹Wݪ�T�����j��;J�B$��p�{p��R��H^��W���q��3��B�?_���O�}��rY�'���Q�MyA���������sHw�q�wfQu�.n%d#���M����13uTLr*-`
¥��w֚�����_��Y��k�����Yj�!f	�,1ݻ���~ԓ��|��9��d�o$�5��~O���x�H	�7��/������-�G�D���]��D4e5�7�'���'P��*��w����(�_W��,�����p�$	\�eǵ'^#�ڙ��|��3�V�7Q%s�u
��,xءƚc��Wh�N!
�Ԍ+���VT0�D��Iԅ���)���.kx�k�W���[���fp.tho)�3�FG�]:�K۱PrxE��4F��F�l  �2�Q���]sn�� J�PZʮM���;O&�Mm<-R�t������Ƞ�u�d�#����M��	6��r�ѰR2�ՙAdNRh�q��#:+읟t~z#A�x�Z�J�t��ڑ��F�Y�?L�ȶ�#�.��F��XE?*O�����+�H�a[���\I�g����]��Q�^�4?<��4��ɒQ� ������M0�	L�<u�T�ϗy�d�S��Wm�`��&�������;h*�
���+�x?8g��>F�K!u���'k��9Y�Cps��c�Vn�]���,ӏ���������X��?tE^�� ����1�!4rk��K��s����"��	���]�N�ʢ�����s6Ϥ��~5e���z�:��ň�D6���-u޽Q�ڏ��H �렣�l�>��j�fS�p�@}�����1��XGP*���p�-!�~/5E�/^c�ᑚ]�苮��v]H(z2��A���bf�\h�L8�%���W��k^��x�8֬o��oͷ�=$[�,j]'��5�$��f�;��@��<hS�?�d�Y��y��8����%���x�#�:�*F��P#e��'�ym�{b��k��l��[�d�(�5�V���5|	�ހ(PD��r��S���[6��R>��)�#�k�������F�����Ӻˆ���5��4�����݆��&�k]�9NNM3�'�LX���@xK�??W̃�l�\�����_A�Ϭ(o���V�L�
�!�J]`�ƽ�� �ZW5���q�T�'��^8H˶�B�#%����8�Z2��rE
f���W��j��PIEk����|�CFa�ױ��{%=�p�q�h^j���p�ޕK�x\�t���}@rf��v�`��@�`y�)�W��.&z �C�8��e��C���y��4خ��ū�T��Y��悴�CA��o�����t]�;+'�T	'M��H�����F�e�/��Ą����P+�����
gL"e��}�����7/�U���RiuV��C��c	��4���#�.M�㹗e���J!a�6���#4=o6�陝G�f�@��r��䲚������1� �5ݶ�$��3n�W����ϓ �>T���g��	}�#��qS̆w7��M����o��7��jY����	X�����)���Y'��1���X{���]OR"Kv�i~~��X�ԣ��p�1V���J�Ԭ��nDLћ�����9�b��\����;3+<=�+*�v��K��pD�;l�����������*�&R�[�;�����\e]N�"�v ��t^���Z�KF�K�C�Z�g�ɼL|fuW4��竚[���NE�f�>�����������ވ���TKķ���"��N!�c�М�v��*d���}�isH����V�!{��))*&�l%��8��e�X#0�$�~�Y�y�!^�{�,5[w�LOhm|�,��8���X矛�u��E̟�gwԞ��jS����@1�6g`�̻:.�)ޅ�T҇� �~��|cuT�]���S���L=�5��̦�|)c���'��w5a�/�r�Ɋ|B�?�ce���]�z$��p�l�S�ڀA��̿z��N_��h�:�?����A���I+�`��\'c=�I=J{x�4fWg�]�sԮ����H�8Iħ��]e2��g>�,L��hb�CI{eal�š�9~ұ�FQ���Y��KU6�_�_��Y��[|?\��xmԜ�c�S���ȗ�<�TΊ��3� ���w��sB����]ɜ�m��f�����(�k�k`.�z'���\6s�:g{���+�ǍV��<�c��c�N. �����rj�L�(����b�2 R^�9I}ө��WG�ŧ�5^I������c-�Vإ���|kݓ�o�� �ޒ�s�S���1�T��gu�&r/�$l�wY8D��nm��m�6��h�����`b��O�&�_n�㶳�au�{/ \+�m4�"��m�
��o=��f7�_9W4��'0��#��j3�7t	���ן�@l�J�y7�4{;a� ��C��5�`{��i&�E�kQk�a��Iޅcey���ذ��5 P�ܪ��AB�z���ץ�בK�Ưf��* 5��w�}�wA��˝NL�O:뼕��\i��A��>̀��$�犉+^��j�E�K���©��;��o�]��*f ��-���{i��R�u�j�l�x�3���E����'�mǩN��[ނr��y��j3]�t������e�4<S���`��ͱ����?Cy�4���z(�vd�J�=?c�8���ǖ�/مrA&z��~`p��"��K�D��/��৊e�or�TWF���f6��PnVu�'�y�h�����@�f'gRT%g�HW��Ox��
��>��=�N"�^���i�K�/������}��3�nLEfr���,���"��!6��jV�[s�P�����2k��p�_��u��oE-O�[����")��\���/��\!1�͵\̤�m�l�b���,(��E��{x7@��j���o��N�(ҫ�%��"��-��Tq�u\n�-j�q��O�j/�SZ�����&���%�F�rn({�[ї�s?�,�_,���s�X�^)V
��s���vv��ݬ�"����s��C5��9�-,�6Į��L򴉳�J�����ů�jv�P̏��dB�(;HŎ,�n �$Tq;#��g}ŝ��5)��͋YE&�,� H�QO@g��4-�I���3B?���8��h�����B�t���<���۩+i���jFrna#w�y���IX]/T`ԟK��PPZ�m|w����a"gCyVe3�����z\��*	���t?`��W����?x�g�[ɋ$|������U��E�Ϫ�a��˚������b���,�mf����y��^�]�OxS��M{3�.n�n�&;Vo���uPQ�=s�K�Fc�{�����pl��:�e�(�ں�ٔ�qR���E���r~X���vxk�!����x���[�G�c|c�R8����̔u�!�����]On��᭖�#���a^#:}O�B+#�9�����Ox�]w̪pQ�s�� uxޤ7EV<6��<N��^�<P�{�oH���LU*U��JV~PhA��8%%�l��enry>,U�g[gV�rƂ��D(�NQ/�]���
�VI�he���.���m��p��d�����N�=`FU�}z�F��A[� g�_è	%�d@B];�|�uR�Ѐ{�p��#�"�p(Xf�8��f��1�_���V1�����F���#�;[Yq2��ˍ�ў��Lq�y���#�,{B�d��#���iI7QϚx��,��.e�yٽ���G�-;R!��.#r��	V��7�S�8OFLe;�|������Qm�t��O	鱦���v��#q�RdRi�!��~(�/�O�3�p΃�����;1+�L̻�q���@v��W���&Hk$�(_�s[.��y��ekRb�h�/1��׍,���Jk�ܧ����kx��N<�DЩt볧�!���@&g�����[��Y� �����}��-5y ٟ�G9�hus?��T�豔�n���cF���J����x�� A�bB�Qt4�ƺe�Ւ������}�Tla6a��a���=t:��Q!Q��pJ'?�<��X.w�u?D��`:nԾ��t���.���˻F0pl�
yp�<3�%�ͫ�F ��6�D���a���ts���fJ	�6����"�=�y�uN�]_�^=���z&�{1�&��\@;� e�G(`��t�I�}��{��E��{��x*XS�<�d��oǩC�����E���Yӓ�Iq�y�2�N���pȏ䤴A$̭W?;T�����R�Bv2�E����#�����H]�G����\|=�i�=�n��8U�%ݯR�Z�E�Xz�Y �Qw����I:(���߼X�~ּ�\VL[	ra.-͉tL�x��s~� �g�
q���ۉ�ar�-�c�/��I?�tf�7[Y@�^�N�	�ˀ��_��Lj�e?v"�����C��/*���/;�������V�ZG~%,G�ר�a�	:�P�J��5=U��9P���"�MU�Hs�=-u��/���/g��uc�z��]��g� 
�Z��EE,�#�/Y��<�6��|�;��ӭ�{�}6�#��a-da�D9&d�|�ҋ.�%�x,g(�6�uq8�E�]"�� �{�L��G��j��G�0
;�s�t�jQ&�a,&c��[C7t��	�i�{�`�u�woQN�S�b���9�w'B�CE��^�.c�6x;��rث^V���`��$� �U�`�?ӥ�,,�in���^�`���7���f�k���)�����ʉ=���ip��%�*�IbM:C'�����g�p�2�� D�ržB'!L0ś[bS��r�����^Gj�O~;�v�=\�N�]4iN2��=Z5+�L8gG$����Q���;���s��3��K�7F!��Bh�W6�?�'QD�u0m/����r��	� ����> >_b�d�jed6���1���O �p�=�D�EM}O��/	t��F��D�����Z������u���ܼ=dE��+%]_��CE|Bc�b\�tc���0�X�O�;�؀#�F�j;L����L1$P�M1�й1g�b�1h�.�n���Z.�q�S��y�R�u��~����%��)�ϵ��y�-�f���~�8H)$�� h���h�ں�=K,�������
z���U�֭���vp�!r9��V�z@]�&旝=DP� ��� ���k�s`efY5k���_�W����e�����_�Z��ӄ+ٜ3���"�e6�Џ	.��Ys���T�e�U-��y�2.�|��R5���{¸����$��H�`�\���k����[tW��r�R���8E��b�
�
-��Mi�E�5zޅ�⯟���,��Ѥ�S�L9����82�˗tW;��ѯ���"c
	{(�ò6������,�s(tb�i��N�Ib�[{�]�8s&0�
I�pEC�L�S�)"�K��"~k�;������� Kt���mx&$��
���A�����9�G�N��uhoulk�D��3���y,պ m6���|�[	�^��K�I�#T���#Q2�``�(�u��r���eV�r'y�+�ݲA���Y�FZ�M�'i\���p����,CUpk��3s�}U��m�Q/�&�Tk���H����
܆��1
uH��­��3�U3��0�!���g�,�������ZC{��b���MN��w!?H�c҉�?�֟q�-�ڋ�8bY%g�t��|��v]˹Q2?�ؾ�{f����3�Ǩ�
��W�,B^h<���@��	�?�`#��E:�縙c�&��A��)�A'}�;F��8S<¦�rN�]��2�$�P�L�78�6��"Iػ�>�{}��ӳ*�R�T�6��d�E���c1mk���6J]�.��0�6��"^d�W�k�=ж�2�Ϫ7-�Y�������C9MD�6Z�}���g����I�O�_ם<3�~�;\�e�S�����};ED����%#�ה���#�В"�3p�v�)�l	��Њy䧓9S]7P�G��R���3b:��+T��`칒,�ŢN��7mX�^�l�UI�{m��=:�r�;����)�r��r/�����c�����/��d�a@�MR��yy+A�ޅ��u���Am3w+�ŠhbB�x��ύU�O����.��{Ì���������z�w�-�%#v�Y�pO��Tr�F��x���	l�O���W��K�%��b�o�v�[�OԂ]�P���A��;k�����������yI�+�B�O&�b/�X�j�Wu��h���
h�:2$�{�<����
d[���l���.�|_֤l���z��`�{���.��X��2@ɲ~�ڀ�8�ȳ�k�K�9^*���;EN`��b�D��ft�ʻ���ഞ��Br%��녖㠮œEXzJ��O�?7�)��Oݞp��z��y�M��-�b����Z����ϛ��C6�u�Xt� ��[s�~ȋ�UZ�G�[���ޏ���k�=x�2��𥳼�uF��O�1R������;�ؼ-w��T�y�Qa�2r%��)d z?����9k6�\�,�r����?���v�!��*@�VBt
��r�l�_�ۻ�}���B|��$�p36a-	�_$�Z-}�C���n�A�0���D,8�L>_��H��Epd�)
zR���S�X��=��(1v�̜9=��W	t��1:ůz!e��𴤁{_�������RSFT}U��N���~����3�A�.M��þk���-���2]Ԃ� �rY��P��^���0�%�8&T�$V�$A�Y���i�^TRS)ޫ�V��(�����Q�'1��@eQ���b9M!�ƛ�r\N�ȸ{�<g�
£8Y������`[�K'M2���i����=�ˠ�we���Z�q��4�$.|�F܁eR�d��x��Б*��h,�_ЫDv>j)�	�H�zq݊�\ؘD��w����C�J��[�g� t�h��z4���|h����w|HՒ�Rc�ٕ�>�C!�e��(܂�R�-"�;Vߞ10g�+l�yx��eG�������^|�<\����؊#:��tɍ� }��;�]�����l�I��6uq`�-Nި&�B��	~�g�[ ~Ad������M �+"�8���
<��+�%���b9�[��{S{!��s}�|�Y���3l����]vp�x��W�bv���ȅ���$�ဇQ���љ� 	��u�˔s�C�6����cf���1���N	G��6
��5}u|��pU��\C;m�]ւLu-[��[�Ho]��h�HJ6$������g	���wЄ8����:3J���y��K�����κ�IDka���*�(R�U��ň�Ư�9��gz'�0[=HoZLQ[�G�aS^�9 s�P#����-���y/��'�|g��~2�\�����,�T]�T�j� Z4ut��.
]0�cC��j7�$/7����	c}�L���9�m�W�g�௿��W�#`%��[ �_�o(|�6�k��?i�]�ad�'�}o��U��ӢK�V�ri�Q���`~~s0(��8�M��5�Wp}K�J���N�s���9��`5%������݄���d��9B@��!��������m�b�z"�d�<)g3�6��!��4^������S���U<���_�����7�CܻE�q�?��;PJ�6��udXؘ���5I�[�y��.�|��;%$``�K\��F�*�~�#��=G���c<;"��JEqY����T��h7 k���e�Ѓ-B���&�Eǌ���h���[��_�ln(�g��	���@��������(�������>�7���6݊�~����0,��Ṟf����	��9�M�|^"ݾ X"�V���}��*$U�a�A���.!�5Iض����չ]���,�p��,��5�\�"d��M��~8v��-f�a>��0�=�?�;���u����%�[�	C����{�'w����]�ٯeYP�� 5�fE���O��9n���M��?��X�.pA�|h5����a#*���}��=.�(C�)�f Q�J�z�!�j��ۃ�rW���CV̓��3AV�^yIjTY-+&R�~��šf�ݫ�����V�ǵ(2%<A�X<�R���k�V���)�b�l ���N���t����屡Јw����̗nH��S�0�Z�a�}�Em����h��4[��ŌXr��S�?�i�|y���ٍ �R*C���{ix�b>-Y��e3�AgN6H�}��6����T-Q3���^�P�|�0�戴,�E]R/����	PjD���$bIh��@E�V�+��y��-�h|~�?\�RmNmR�8$yB��CD����5B�9�%��3�J3��$s��L0���ml�v��˨2�hA��?�ȩ�;u��n�/�Z)�6��%�4�<�?�w�2c�gM�����;©�8�� Ga���q����Γ���/	^���8;d�;��m��3t������/4SS�h�?����8����Jr�Sq��u�s�l�In�W���;0�?o���Y1��cW+�*$�NO�Y�����68����k��'~VV����~�)t���������&�q� ��d�ZȰ����ێw��F���B*Ԁ=T�w�d�ɀ���!�>�T"�l�n�Iu�������x��t���h��l5^e��vSs�Û}U�A����IFr�?�G�H���,�':<�V`�>�nƫ����U�7�*ޞZ?[o�4zR���そ�i�XRו����]����m�ʮ��A�g~�)��'���C�p�!��%#��0�aC��k*D~>�.M�2��-�rW6�T-�7�wG�@˨��P	�O��@80�T��]m�����(7c\�5PUV�1�Zի�j���5���P�N:vƕC�1��#�		�ifj2q��!e��@V}�e�Q��f���T޺Z������c&{T��6{1\ބ}�]�������)�&��6��o�6��8:��eR�A}�$�zp}�X�lV����݁�=u�.���@�~[�������fDy���!d��
Z�n���g��
�/O|���������IA|a��1͸Zc��x���n�_����[PJ�� �S2�L 퇋:�x�mS��^���o��)�R�À_F�'M�lu	�[;����J�)�k�	�),�ňּ���h��AîyDMb�@���)yT�rrJ���uz����*Pw����j��q��sjv�g�Qg���o1[g�&�UY��F�ɂz�I3�g�Kk��cm{c�jǙ���ɀ��B߀o"#Y��j�H�>1���E�D�掩H��Kwm�y���z���t�9��Ҕ��jO��\P���?.񠙵����,3�Tg$��~p�>�~6�A3N�0{�;.����uG�]�G��$C}sb�9�Յ����ϓ�n�O^x���t�}4�����8�㎎��c����3��7joFM�5��h,��j>��-h�ܣ�`b��Y�B�������}�jeA	ǌ���g�ZB'?�1[;^�`:5�r܁��3�:�)� 5}a�g����)��Ҙ��3�P҃����s�.���փ�����%����Z���V�s������dVYz����@R}�����\ �~[��������`��״�
ϝ���1�PL�0�h��F ��Gި��n�xҫ�$+E��w�m���]&`�J���Ś����	�3L;CQ���7����a��T�]x��GD7�e�맍R���?�)�l�@|�ʅ�]
���A�w�d�g d��+V��t"�݂�RВ� �?�"������'��,�����8�C�a˿��;.�����^�o:�q���"T�P5Tutmϳ�R���b툖t�QyG" ��:BA� ��y?�S��p��ݙC�t��?M�@�!�$Ss����P����@ćt
[��;A������,b�d�k�c�X������|���d�O���3�z3�<;ҽ@^�+��� `[��\� k��oO��ԟ��4o����? �p�d��)P@�o��ǥ�[Uo��+�<m�9�f@����r�"�"��U�rm�tA��.<����X�x�J����}�k�R��#|N��@��`�~1=���X��"�e��Ɯ(��z�gP9xh�U��'E��g!�Ǎ'�^���6A#��A�>?�[����O�D1�}Tlt�2GHo�j^u�[��:���,��0�c/���m\���%��!�|k�I�;_:r+.�N;e�a:y=�6���M�94�7q��WV�~>�m�"u<����|��6�-���9����f4��~�ը ��������}���o����T�
�����ⴇ����0t���R%�>	�j0l��Ζ	���h Е�[$���ب��.��/�+��������\޻�s��;�$E��Y<��= >ڞ`GoBԴ���S�u��G���^���F֥���//��Cը("�DW q\�&G�(R8�7�q��E���Mٓ
�y���+&+e���ƃE�K���u/�=hxy���b���L&���'�j����	�K�Y���S����@�q�B�uؑI��lS*#ȮvOc�_R�<0��U����"�()i�����Z%D,��d��
or�gf���@>�<¤����L�� �ǥ�H2����vvh���,h�,}Y@m���1[쎿=�
�<\tj]Z	V19��C�W�܅f�l�z�3{w��*��Dyt�O�# k�2��o����*[%z$�S=2P�X���o]����W8�O��H�&>�^`��U���d�U��6�� aa��D�@|��i��G#��0���e�p\uOl�ǳt[9S���<�Fe����q�At�T&<�V)�*-�g����޷�v^���@���� 0����U��s	��j���	�a��3�����o���B����¬��+D��.�ӳuy��H+|<1T�(и¦2U�H̕�H��;��l�L5���*� #>pDH�j�?	~t/Y�4��.��lK	�2�!lK�������Ƹ*����`�9��[�m�Ó�͛*���欏:A[G/�Up^� L��,��N���"��t��e��Ok�H��9�ic�Lɞ��P~%�Y����3��Ͼx�եx�1$0^�Pz�dXsX�\�Hm�|�o��(��V�
ּ� �MW q��ߜ��8������g%�AUw�ע��n���'()p�?$i�A'׍���HIϖ6��x��)�'"��_eb���q�R���Y+�%��a�kZDY�ۍ�v�lA��4KO}�j��v��c'���h�Ŝ���?���>j��a�m	Pә借�����?�G�^�?���s_�ӿc�"a�J�UCW\��	VCr8]#M��i�1Wm�)(gװ8	}
[ғ,�����ซ_5�Ts���da$�'̞���R�����wR�����\�X$R;�S�p�q�nF�J�O3��[3|m��z�$M�}�p#���PH%3�c�k�Ы���(�<�=�0��@���[J^A��%�a�B;޷���մJpԯB�y�#�8���{�l����S�:e�}W0P���b����N>���: ��s
[���'��lY,�U�_v���~j�q�d��\S�9I���O�b�"fRc9ݶ����]}�t4�\�%��-!nzjP�������K�/�Bݤ���A���� �]5�	E�E��,��e�t<>��7+��PF��U4�������Gf�4]A*x!�~����UA�B/4������|�4��ރ�S]�k��7M��)x%��H��]1D e8J�p��j& �����,��)�uG&p�nˏ<*q��O�ô��g~_$E�d��{�BV�N;rR�"�7�e��L{�g�-i�w@Y����Rlx���fN�FbS�f,��b^A����E%��:�_�]P�r��hC������#�����M�����?[~��n�j_���{U~?��m�4��G4 '/X!��Y�Y������Ο�Pr���RhL��j�JH�e3қ3�}����߷�6gz�I<�T�k��jAU֋-��'��f�3����/��Y�߃m�ɩ:1��
��S*�����e�t��Ko���/-���o%5T�7�bB�iLv�moE��b������<a��fhXyU����٧��e�����.~[t�����Fe$�o�$�IIN4��Pf�$��}ߘ~�	�<�<�׿�;ѕ��L�D9a�@h��撑�e�	���<�M3"�h���f�4Z���;c�e�{�H'����T�*>�֞�3�����W��ӿ���&��Y$Xwu.����{U0�E���\~6?"��)+~E+�WHտ�l�j2�rs_����jDw*�퀇�X?���/�E��zՑ�]H����-`3j�ɇ����#ͅ�Ѡ��84mƚ�7�� ��+���ǠD���8޸��/Kh��������C&�!"�>JjV�΅ْ��.���yN�g�0�V[�,-��!���bdC�̊I�h�Y�G����6��b��o$ِ�Q�����y��v0����#s�����%� �F�ҋ�o����xL��Jt��.�����N�ܫ��i�O�U�/<��	�ǅ���$H7�����6F4�n;G���#��;sRGR��3�<�~fK#�j�L��2@��RUJ=P��=[��4�9�e�tLa��Z[�b2!%�ad�; ��*������ha�<$��Y^��Y�z��W�Xgcy����k����ە]2s+g����V���A��X��uX�P-2"�h��)��:I�Ar��z@��1�Q�����̯�����!��=}�l��9/3��g��ݾQ:AN��^$�5��s��s4��U�so>��
�%�ѿl��I�`"2�*�v�,*�%��@�E*�CtÝL�R�kuz�ڶ�?I��+t��Y�
�O*U��_�8�?S���!��Q��ߜ"9[L�sn�5�xe�v�u�k>�~y(j�s�e��:�S�ެ���֎��M��l�&[��ё���)>�1���0�v�gxh�}/���/�?���5C�*3.oL��W1��jM�h�c�ԧ���)��.ګe����W�L�~ %6Qc�$ݶؙ�L�	�����T���E���r���D����-x��.&�[����"�Y���N�tD	�Y��;[0�l��ӂ�5N���11m��ɚ���@�P����Ho��d(��̯!蓒a��������I����߽sۖ��ʲ]s;#�������y{���y�H�zK¯��]Snz���B�^���Xp��nB��Je�>@ �+�%��֎�� �㭚�qd���!��[��R0��|�,	9�B�:Z�5ސ� �T:MM_4o"o��'m�c44 ?�C:�9���Ȳ?i�U�w�p�4l�E:����2��t�nN�4c��|�A���qF�o>3�΂�,]�d_��Dr{c<�z*�K�]�C� �7��/�)3��p���oڛxjŭ�s�y0.6�
��	��p�@mhy!�Ě�D�C�7����NX���#�Z0)�-@�h��e"A!ڊiz������i��ؑ�Z;�A���B���9�KM�b?$T5�,�c{X�H��ܰ��KM+�����������L�%�*�c��Q!sC0f�ǟx������+�I<�l��8��"�6v�Gr�q��Nځ~OF��9^��\ �,x 1F���֠?b���d����vD"bdsB	a�w�xijo׋~�}���e�!g�T#ъ���EB�iG�G����~�(�=�N�*{7dF>I�p��+��{�Ŷ�r�J�JJaz��f�G_��< [ai��#FI��]���\�u����˼��w���it݂�[��+�1^L���.�G�bd\��DbhI�.�s�˶&��!��3d�y:�P�Φ�n����1da3��y��:=T1x�,�䩪�#T�ѓ��F� �W�'	,q�������'>ę�R�?,������'!s�=}g�=(������Bcq=$�J�{���Zd��ƅ���^DC)B����!¼E�1ǻK�A�v��A��,
	b2Y�fwE�p�B�CGm��l�
p��r$�x����4�����S�>��
�#ot�Q��'I�tg���(+�H�r�Gb�].�Pkީ۩��	�l���r��H�q~A۠��N~����#ՔI�H#��XY�<���\)P���є��/lo⃓�'c�vY�v���q$������-[�B+�����:��N)N9O)�L"�ZM�d��9�5� ��e\�$.�CfIfr6/F���$�8e��#R˛3����o��������w�i)ג��pP��r�'[�G��p
V���N�C�7Yqn��k#�L�I�=(@KF�
��-зA]Xn�����;���� 
�U:��8
�z������#4\]6���r|8�Xmb
(�\�L���MV�̖^��+�Fj�� Eݜ�D���83$��G;)@Z�i01nO)L�H���˻>����s��3��gg�����н��>�Y�z�=b-�M6!���W&�L�b�$���R�W��Z$,Ϫ޾}�$0��Z�c��`�b*a�LY��z
R�X�������-Ûz�KE� CH�e� ��� 'R(�e��d]�&N��Dx���5���]z֕'qD�H�M�CҲ}��ͦ��P��j���>T.<�'�ݦ��5��0m���P��I�V#P�P�%#�J�ݎ>A��bJo��І����	N<A`ַuW��n�j�Rn��QHؠ�[��unn��Y���.HsX;���[�������/�n)��~	К?l�(G׮�����7�_��D�7�2�ɳ(�b�^Ii���� Q8�p��R�˽7ğ�m�м��۹��f4��.cC��)���.��h4�Ꜷ�tb�Q�t��ˣʹ3߱�]+f��:�K���"��CK��z�y[��%ٿ�Npxl2)C~K�Y�+��yp�j���l�a���&i.����4�%���.��̵�!���t�V$�G�o�lk��fs�hFA۶-�u���T���9�su��{�Pz0�
~H=���\���YN\�70s�oH���g�w�#���
Wߠ�f������}����.�5��΢-���6����Ň���f0�KS�1�QV �c^<�<��g2�l�h=��/J3<����`�ƴN��Č%���u�����*��r���K|��VuON��@6'�Ý4�q�6�K��u:v7�I���8�L{��F_�X�~��E2�g��g\L��ʇ�h��na��8���Tb�z$ I�ح-=�n�F|����o��L��."�t@��C&T0|�EG�zu �5�������<��Ŧ�S����I9�y�naT� o��/�o�-��@�\&G�v���I5~i��
��]2� �� Eh.S�To�Hq��8����pMAR��4�@+z��H�D��<��	�m}*�ԥ����ß���<��w��oB�&����⎥\�9S�s���J�@��(���nl�m�z�Ԟ��,{&��f��{���V��{��ЙY�%�ux��O"���t�� 3	$j�0�	̞Jh�V$>��U}nG'2�#C���}8.�w�Ҡ���9���C@�R=yD1;)z��M^�����ew_�|�֩�;*P�g����R������j�"�N�ς�j�af�l��ĭ�Cb�~���}�d� Xnd$N�ؙ���u#�Փ�KCa��$��f8�
S����scvA�3�®�^���J(e�	@�ֱ��1�n�]=x6��،aO�Ϳ�&U%�D�;��	Nx
	����P�FXX����P;/�.Il���h_Nco�~W'(Իo�݉R�fEsm�%αj�F�Sw �99��^e׻�s�`e�ݖˊ�:��v��ݫ]���x�u{h|)'��J������n��ۛʯm.۹FhpO�t�*qw���Ϟ9#ѻ�P"���'<�ҔC(~�({4x:��gohx>u"��+�m9��v�;�����j&�|��F�^�����pa��T���z��������-�Ml�RU��� %�8���R9$
�mlҔnO�vn��q?ݘ(C-3g&�6�y�fa�)}è^`����$�st�#8t��9f���FR���@$ˊ��=�k��=zvP{*�%S�3�`�C�F�2R�T@��h��3-��&8�"sR�@M�ZYԾxy�9%�g ����������٭�P�eŠQ<]&�݊ql�uf!��@����U˺�b��Ȑ�A�Q��7!�T&�� ��hZ��hɢX�{|�R���K$��>�r�Z��&��!�v���7��T�#b�����[��wUDp���~.R��߭s��ʊ�8���mJ��g$L���V����Ӎ�]?�� F�8Ї?� �,6Μ3Ғ��f�I)�pL�b�sCb!�~T�i�2+>���,��k�-�2�D�R$		x}�~
E�+[z3��Ѧ�}��Ө#6)m��������b: "O��0��{S��7��F�?e�
����ts�s
��aOLt���!��,���6�����"�$�g�땙��KCS{���	���! lo�C"'�m���B�'�Ñ��������h^�?p�~�A��B�^ϟȨ�lu�y�Upu�'[�><q-8B'upJ���-'H��r8�ܰȾ�K%@����)�i- �����zܖ�k��Ê1p�W�.!XQ��tR�V�VW�b��W������WŞ׮�� E���`mM��H-���G���&�x6_j�`�u/+9��BnBe��B��Qj����k����y��MƖ���~���Ցh]�\������I�Sq�P��sb��꛺0�����T=&��]��zF~o���;��66[w'�{A
0��L��ޔ�t�꧜�9�:��T�u��z�����Z��/���D7�����I���6��O�J�4�j���{OJ���	_�{�Y���cn��²�W���Ex5�J��>b����^,�b{�s�1�&.�럓�35P��]ϯ���؍Z�;w�s(n>�@$��Մ|)x#�<nS��7fE�vw# �'��
t6�lz�����}�y��Z�����x��Ho�	e$��'��l�ǅ.�ڃd���1X/�q�o;�1��U���lh�6���+��1�e1��o����M��#H��&0�5���ư�ia�fb����- ��]�S4�r��_؋ȸh���
i�"T�X�`�e�<4���a�(���G�0��3U
��
�;�QB�w�u�k�ecM����rb6�Նg\��ȝaܮ��'r#�r�NfSZ�j
����S	ZC�֯o)��2ˁN�-��8^�ݢ� �n��J���N�a��T�bƽ7�!�V��5<�[��F�>:%��>�w��M8������As��Ro_�F�ח���^�����!=�������Ng�:�ܙ���C��í��J.�e3d:f����O�o�S��ۜ@j�O0yK-9�rH@:B��u���O�2�bݲ��K:�N�m��R��^�ќ�)AK�G���@GQ�2��Q��11Τj7N�pӘ��CH��U�7��
���9�_}!��B�L1Lef�����:#%n��Q��&ۉ������,�P�3�k��J�C�̍�O���Ҝe:q��x��k������Y���8����üݽ�6j��:��I�=�.e��H��J7��aR%��Y���+4�N��1�澯��C��4P�k1ӳT	�'�dsV�g}҅���]R��O���1HTr��qgGk���ϻ2�� ����fc�����r���4Q2W������[uVwA���kN-���>*r�����y=�A�,�����#��\`h�\�*�O�`�\]�5��E���6��!�5	�g2��(�r�ޟ�Бx�����0����u"J�L��Yv�,�A�Uz|��ӂ�ﻺ�B��)�f�eK�A~TzB�`%E��GԊw�<�~�����Z���ީc���m�d�'A���@�e�r�uoow�����Q/�zt�:��뜷f�Xю�f�`���J�^�2-�!o�5NRd�qݏ���X���n�mOд���S��i��a�;��Ю��N>�N�l==������5%D���>���>w�[��4�ʭW`����O��z�����W��K"���}BTs 𚫴YP�'sN�ȵ����X�1I��TM8��L��Ȕ>J97LME+fU�e6��D�.Y5�x�E���7� ִMU8!����a1dml>�e�?�tlƞ���p�.�;�*�w"P��Y���Z{2,U{��tw&Z��Q1U�dS���#��[��t�����:(ڶ���;>���.�
6\��G,�n�kݙ�;_��<��t�������R�ശG���:,B�X�����W�����y�G�a�T���lK᧭�͗X�1{*/�����_�4(��)C�Ga3`+4�@}��X68�NfXx6�\:��U�s���ݶC8X��NW@�u����z��L>��5�3?&��%�ف����ӄL���p-�B<����w<��4qhB���e���c�њT �bn�'���Xt��̂#?;^�<�`�P���E��[ VLSS���rK~0_��cA��X&�$>^<,I�~�C,U��n /#I�e������	cϟ0r��H������,3ΰ�/-|rL�vʂP�l�<q�����4tr'T�@[|�"����W���?�~�q!O��Irj3�2\����;La�]����.���g�Z�H�]m;�c�1Ir�S��t,~�ir��ۊׄ���X���y-���ćxon�}�t� c���5�蛹��d=C�]7 �V�[���REH���88�5~���tsΒH�5����i�`P)�z���Q#�R���$v<�"��:Z;Ȁ{(��25S&c�ݧ��iӈ��#�SR�SG0�S�
�)�2�p�U�te��4	aRǩ��4xΪ���evv�v5LAێD8�Ֆ]/�*�X�Ú���_��"�ie�p���6�(P��&��K֞����+"tC�Ql߭��yPYv�ػ������KE0F:�(H�z��
XT�d��yH\JS�!G&E���Tz��$�C|~P _4Q������"5ꋒ7[*ǔ�[�=�лj�F	�H\��a�w�k
��ڟ��S/ތ�V�D�8Y<�ǆ����ڑ!l��U幊�f��
������m�0L.�CV�{��X���*< �RO�����ۢ��ڧ
����W\���	o�,���+������,o=�Vg:	�i�ּ�Y�c��@QD�K�TD���V7~/�UK��T)�O�����4���QN.K���]Kx!)X��d܊�T�	}l�Hwc��kOy���7jk�j	ʒ�H�D���r���7�~Q��O�.��<��a(�Iݝy�h�%i��C���S�.�c��g�- �i��fjZ�IU���b
>��+�=#���J�T���/P_gl���e��u
\+�O�	�Ɔ۶|���hP�IoH�b�1��$M���0`<�!h��D-պˊ:4�;Ѓw��@�����2Qm�����;H�d1�Sf+��5�O��X���V�� �N����X�ڊS�ɝTq�Q��B��탯�#]��Ц��ܼ�A�/�ILE8T7g�=L �L��tC�����SF�1��c���y��*��i8�ԙRfZue�B90�#P�����Y�����>2K�ozʺ;CV��`�ܻ�fbLO��'7]�u�zjL��H���t�?�b�9�t����٤:���U�E���on�F��(�`T2Mݗ��g��tt5B%_0���*��@	6�/
��.��:ѱ7�}�$l���&�'���9�<r���<-�A�gOzf�u}A�F-�(���0�њ����I�FC�!"4p�Ǆ�`���D�w���]�l��^�p�pc�����~�ĩe�V��OO��7B����g_��EɓZ��W���ٸ���!: ��w�#�X-�������nA%��nU��wk=�0���>��ifp!&���X���P�dch�������Ie�xyT�\��}P����:..p8�g9ub�nZz�vV���p�4#i�'��8�p��ZK{�J�gHݘ�������X�}P���?d��ݿ�L7Ot�+̹�d���T�(U�k�wfЩ,�><	xP����Y�sA�YQ�eN����Z�wn�I:Yw������b}p��Ko� P#C#��~G��� ��0^?cK��?u+���� �N�ͮ�&�eIԌ~{���6.�ğy�Wi�'a��)�Y" ���7�#��2������x)����z��f��,u{<��%X�H�R���v�����q�t��B�m��yY�GS��Qi�<����'8[
<6�.�*������P0͚����\#<�Y���ZN����x]9$vg#�y_�R�����".��P�C��.�.�YP�*��j�%ʟ�P8���M;Y�]���[�(��\{Qc�k���E/q&���9P��{�)�Uri"e|A )��굼!��&!���з��[Ů�~v�aғ�-��,&E����Ro�1�,���*�����gѩ��/L`N����*�.A���B��;B|���^M(��
�Vp�(��Yd�g�Z߶��ʂ��ޡ%0�(�#}� iʵI?oi�g����a�lXv�r5G�v�`{��۫�Q�b�3��� �C��|��� �y�"�q�C���v;���{c���Q� �J2�l���ʂ�0��:ӳ�Ҁ$*W�p^�Oe=��	�g���l��R[��55�7�ME=1�����#�KOQ��� `O��h�fSfS�;���tYS�/]�F��r�"�f���|�������0	� �s,=x�k�[��}f��ˇ�@��X?c��
�j��r�d<�˛�J���F9ᓦ܊�є�!B!������u��G���E������`��oV���R¹��_�
|����-�EKx<y"b��A�zKC`LZS�>�n[2�'�+F��[�Vh-�z(M�L�Ʉm��ۏNC�$��p�N�����ߍ�~�~S2Hh��A���yu=�R[��}qg�f�5�=(���#�����q��v�V�b��L�����`�I���exu�T_�$Uŭ$'s����}-M�!Or{����Nָ!ɠ�]S7��H �>�ֱ H��ܣ�O��et�<���VA���댥����K�X�O{�ڪB�a��f��Y��h�}�����G�/�ﭬixDA{�
�_��6<��{d�4Δk���nHV��e}�RO|0ۑ����o	U�	�< 6� .�S����Ő�n�r��H�0�0����Q{r-2�(˛gt�j�V�Ɓ@fsD=Ң�!�f((�y��vե)wk�f�����t��_�	��=���ѠJ ̈́[�������,�Cf�����"R^ԔR_!Z~
��������%���ũ(C����I��{B8�@NX��8�yZy�nF��"O��)��W>�C��͞u��GJ��	���G�t�ul�)����Z7!��~D����z!!X}��x&����"�H��@˰[��X2|���6[rg]<s �V��|wn���s���8�p� ,��\z2i�pic-��L��8��L�J��<v��d����wR�Y?����4&���]�ud�BK�]I�*��M�`��sbV�^w���#���#�'n>o�"-أy�jݦ�رn�z�#�����+�Iǰqe9���������13<��w�T�Z՝�$3A��Ѥ�[��)i0���ёj�YJkTO�_�O��#4�,�]��#h��+��ٱ�֡�-l����v��.k��:��a:��p�JΕw�1C�^����΂h]��n�8�#q�����*z���CV����B�ɶc�@6Q�/A�ǩ��W��=���M~T<WϺ|����- Zƌ�}�cJ��h(Ɯ�����`{/�q����&�GT�������p�Mo2��vĆ�|��Cdu�T$��k�u6�\R�@�%W�R���I��*���C�4
)����7����n��V�$8�
)y�X���ʴ���/E��1.�T:H��WUF-7�U��OW��a�DM
 鈅��r:+m���D�v��V�"���< K�K|L��]�F�op[3[�}�X��S�$_�e�����!<A�v����(Es����B����ᦾ���;���s��E�*����V`
���Y�t?}�a#3/ߚ�2:�qMf� Q�k\��O��|Z��u����hօ�ۊ1*�\���x�O�Cyg���C˦�I/�ʂ�gg�v�?��v ���X�����0D�x�*/f�9,��B7	 Y�C�8��
��Z?,-�pSU�3P�N�
R�|Z����bM[%��6���1UuG�����q�er�(��?B��J5�X��(ǥ���n)��B�H5O�CI+8L���4���X�����FVX���s$;�ժP�����U�+�l��g22�W;l�}��x2����+�:�uQq�.k����M0���&��ϱw�}-��e���˖�YT�NI���Jhx��!M�Ą[s�{�{C�!����݄�}/5���rP�T���0�$�#dG��>;���ŏl�7��zݥ��]9��Sb'���Z:�G3��ˀ'"�"�P�A�ӰB��z�,������D�@�+r���ł�R�+R�]�b�U��9"?&܀������À��Wܦ�,�?=֘���( Lr [r�%Y4�Zj���S����P"������%��J��H#rMd_�;�x�f�9 ����m�3ު?˟�K� ��\��.� =������ii\�e�<0�aX"��6��"sd�˯!Kh����K5�I)�b^�k�+J��;3Yv�Rt�:ju.�x�W�Fv]Q'+�����S��E����Yi��	2�sO:G�����t0�E #�C�+�X�leX����[��TQGipT*X�&����;^�$�qZ�>L�o_���J�p���x�A��V��+���p�x9�5K&8��f�d��!����xK�ذ����0���Oo3�QC����ޓ�Ԛ�h�ʣq�	��#�U�lOMC�HN_߲��Xw�9/��=�*�2	]���D�	�މ�|Ј���/V5���6���A�	�G�z?��e-�#={�Kba��e5QI�6��7S��W�ѻ��֝�
F�$�J����1.L�rC�@��nA�-2?��^ٔ Wd<�?h��XJׯψ�SwM"�G�u(���	�{�kgt�z�pr��{�U��r���'�o/�p#���*��sW��f5�?s�\����dx�v=�enM�gա�P0�e��WN�����˷�c��S"s��wk)x��vq��Gfr�inD�3I�x�';?���wY��������C�x$��&78@��)�1P�g��������f���9c�0�d���66����ꜚ�W�M��ܡ��$�MK���������������P�JlwZӰv��'#�(\�ںP\"`bs��5g0���J�l���kY4	�a.E~x*	� ��.��xS�إcL�뺕��g�$��D��\�p���1!����e�	U�O���S~���aE<����菕������/��?��0@�t�e��'N%0/�����O�߮�8��-Zo�lbqQ��R�O�����QM~e��K��C�0��u�_���aC�N'�]b��F9P�53~l��k��}�)uX��[���1e�^��{6>�2��.SY"ˢ���OŴ��שxkV|�E�ឲD�b4/F�YiR�}Z�p�6�~���0��n�tR��k���I���1����8pz��cg�e�M_�U���K�l�io�ZS�xq�ڈ OFP8�#ܰ=�1��j��w�)�`2�;]b���%z�6�{C��I�e��A�T�e�xڰnȅ�����?ΛE�j�\���aN�s3Yhm;qF���Ϩ� ��g���̅�#c��[�"O}A��Xq!n4��u��-;�Q@��;%���`�4��1�����U �P�>Sb���m��ӺN�la�^`�R�����f�������9�z��ں�<G��%@mr犀c�T�Y�ب�NpEfo�j���]��t�
�X]��^~8(y$o1�a�X���x�CT3V^��#�����[����u�e
-���m�� ��~2V�����?�� 5!W91p��4��'<��`����1���)�ԟɩ���B�xP�e����/F���oа�z!KgKhA�O�Y�Y�C�2��F6}���wA�:7���`ff#ǵ����N����-F�gܵ�>�jOU~)����ݬ�O�T�f��o���$���hy`ӷ��E|a���V��"?�:���l��Œ�&��6Jml����G��G��X�C�:p�e����Ńr�e�6�(�����a:c�:��A�g�|~����nUL�$ȞX��hS�^���<��%'��&y����<u?%�Y�
[R�������ϻ��;�$ծ�N@�h�8f�2~ ���5��!���l�F����)��ukg!�L�0�a�@�|��)}v��3��.[�rF�RR��� ��ϩ���iM>�Hy΍R4��敐C��Td@�f�0#���D	�8��w��`V_��?A`J�SVC��4�I�!� HCN>R�m�΄#/�Vc]?���VRF=R�C���v�f��h��5���G����j�Ӆ�����}4�娤���P���c��`�dN�v��p��@��)�6�]����R!�qVp"�04H���ߟ�|:�DSQLs�|��K�'����)9�1�{�F/S��wMl VV	��+A�bw���6;��#��D0`�ȥ\�j�! a.�S�j٦�ň���;�&���%�Egl|(��V��u��8^7�2|��KGR�����u�ˈ��j��]�q����l�&�7�7�B��i� ܩ�~ �jGl��0�Ŀ2�}#���~�oK��)1�ᬦ��ܵ���?Qb��٫������H�&��G� �f@!L�g���XM�E�w����� ")"�n�ָD�|�u�f�f�Y���<�DY�^�5�:�5�'<���P,�놢{�q��:2���^C��l�3��r�fy�v��	��rƾ��� �0����]��u�anb=��+@��`5u�%����Y���%G��-Bם,5�y�0n:����
cFw��F6�G<+�~R>�?��ɕ;"���*$����rJ/#�@�"���Q%E�ài�2T�1�t�C���3���zu��P�I�B�	t�?���Cٮ}�L�
D�<�U���bo���q�_[��(�cmY�nw��(���vG��p��ߔaGZ\_��A�Ɣ}*x;ώ���5���;r��ئ�{d����ǽ�VX���lm���D<����D��3�7��Q�ǽ΀7�rp��oer��0!N�m�$�VpN���KA��L�lC�I&h1�|&�Ƥ�^�X`�F{U�*Zq!�ռC.(�I�t�ؠ�x���j�t�Ჳ�Bb$b(J���4X_Ч+Fj}�`R�9�d�'�e�#J�N�����OX��2!�xH�X��<��)�7��>�*�Y��-�Y��_e���-�H[MD(^�b���.JWM7:q~ڥ���U��ctT��S��$;���M����֒0MI��/��xJ�m��}�����¸��tlӜ{�d��(eQ0T�p��6��"V\M +��9��X\� ��)o��w�U�$Z�>��@J�A ���Lu��1B2����>���.w��jt���`J&�$��YYI��U��x�]/�	Z�ž����K��<�p�3m�C	'�ʵq���ߊ�}�Q�tϲ��U�p�Ro#����z��u��V�s�RW�4������2!8�Mj!-�\�΄��~�[) ���cx�3}�-O�g��2�����^���Х���qϣG`u�XYu;e��y�G�`�Y|o��Ea��h� �5����B~��]��� ov{F.d�ޜ��"k�Ӂ^9����;�c;���e_��
��a�O���)v2'd����1\{�t2Ib����(y���}D�����-�8�����ݝ5�B��yD�x�b�t�iB�l�MUh��T�X��W�L3
S�3Z�-��޳�VJ4�]wF���T�?{�Tҫ��I�����Tw
2Y�{:89�}�f���C<^jS�^�2qOs�.���e�\e�xfl�P��>v�zQ��`p=���yr��Y�߶ s��RB����JC��B���5^:ڼ��W�n�p��	;GW�.�0��w�0S,؉}�3��DJw���)q3W�u��8��;Wfn�U�F �Ɵ:#���y "�^(�9_���@�U��}QA%=�:vxI1���`j{L�]�b6�\�u��li n�Sh("E?t��Ͽ�өV�(Ӏk�$/O �'�c�e5f�N�6gHɅ��;t�es���H���TQ�x)�ܹr�ڬ�V窕:I/�������ƳhG�|�4VW����z[q�=�~4K�)G|)Z��\�^c�UpZ7�?�z�IV�[ڰGȫ���Iy��<���S�q��' �S(�)���[�w�';� _�G����S����l!ֹg)��hI��ڗi1��+�š`p&�"�rp��[Jwi͏� LO���<�P�X�X~�IJ�u��QWH����Q{��i�������ڣ�$�H+�`��")W���wՔ�|\�,Y�f<�U(����_��֐_�Vby��T�>� �L�����mW렍��;ţ��!�H���_��l��_ug9���&�a��x�d�dŐb�w��R5�8
� ���?���\�)Rl:�{�cs&�󡇳=�˸[d��;�df��=��4.��]���>�p�ס+���÷�g���q�8dZu1����~�]�<��
N7!����S��������l�n�}��2�w�ךTj�|�[���3�C#`���=)���2=~F�p�b�����4��OS��7��Qs��T����4-�fC�M�H��y�NX�S�"�V˿����a�+ˢER]iĄ�&;�s�G����^�Ԉ�0��ev���i����f�H?s���z��F6h���n.�
�� C����j�=P�X�8�b�2IO�^lW3��?K\���0��Ѵ���)K��z�:dg�O����0��R[j�}���S�1	����:����@�4���t��_������u������]z��V(���#�������pgn<�g��A�rK�J�IeDk����]���J���2±����ʚ�E7���%�2���R�\O�^F���'m� o��4 �'#\v#��2�}q��y�%�1����'�#��m����Y%Gt�;�{x�Yу�
Kp���/��:b��S��_���Z�������$EvنD����-/����롑X�0Z��#.:�_��!�n*����Ъ�L��V�wT'r,-L1�;��v����x<=�]�>uK�)
䠃��FX`�Nj�Y��8%P c���,�N9� �+	`W�$Ž<9;���n��a��K���w���[�ߔs�|�y$���B1�f�槰���H!�Tz-��݁���*1̝��>��K��L dH/��a�,��$G���NO�f�*�⣇���3�N�l�M����,�$�=�L,���9k w+U5���@jgO��0ד3�,�E����������4�rS��Ò����A_����I9���g�5����@��g���Q67[���t��Lb,��6��&�n�T���'Y�˴�@�k�U�b�Ui�1Y=Ip��Fx�A8i�V<5
ߕ�Gd��-��Ϊڞ�-�V\�M�����O<��<C�A�C.���t�A���i/B�1	'[��vC���4to@�4���C�A"dw_"W01�,�|�DO����Ҭ�/?a��|��P �/f٥����I2�\��oQ�%D��^��0 y��A��-�k���T����>G����#�ri9�:#�f��r19�Aav� �N���:������/����,�(:�!U˹�ǭ���W�X+�Hn�� O�H��P�xY��1:��*��N��OBVu3M0�4�p!%���������j�9�� p��N��I&�'Qf�r.C�iZG3���D��$��j��^U�8N��f�_Aζ=b9d/��vޏ�IH}���_�YH�U΢�||
��ĈI�d��^uCLG��#�B��=�\��4$�O���b.��a{����u@�v[��}��������6�&�uP/��	Cc�'+oˀk9�fV&�Ă��~���cZ�_�3+^h�PV��ZAx%��]�mˆ2�;5h��� �K[	/�#?�����������';+�9��;��8'@��x�§��QE�_)��&��Y�JH���ƥ(��K���5�w7���x'�����Qc��$�e!4�����1�9�P<�J$C1bEЗa��ၽ������1�W�����1Lg��z?>4M�s���¯�=4�O���(6��\ʲO�$�N�,�HĴ1!�8���x�<l2U��d�c�!!$أ��l���Ϝ�4lk��e�l�����#���)���1��e����1���%h���}�\�����+��Y��\�@��k�)�s5��#j$�F��f�� �s�)h�ӽ�P4���v�_�vG���Kr� ;�t��hQطg!z��za���j�����������m��I}�K���e"��,븰��}���ph����D�<��!����C�q��,SO�����Z	`�����/�$�+�^1�{Ex�� Ds�9�UA4�FH�>�s��p<ґV�_�yY&�(Ğv���jxQ!I�F�܆���
��@R����5[*�����9�/�`[���+�;h�
�ߎ��<�t�f�G� �W��^��t�Z�	l��G�^ ����#�~���V���8�Y�CEi@����5�S������m�$���{D��T�B�s�s2�]�1�tIW��U�>�VL�q��ۂ�]�������f����3"�t�4�뜰�d��S��z�Ǘ��9򒎜Oo�r�����%�8v19,�.�B���2�������":Ǳ��t��9����8 �LG����C�rΦy߯��^��)߬�J��:N]�"l�����d�ع-�csP�z�{	�Z��6Aal�AMi��*+��,�ĹS"o��+?�q�����x�n��Ry��'c�a���\W�X��~=_�יpZf��x�u���1D�;� 1�qj�b�((��:Mv�lz���ߊ�0��\�~x+ߵ�F�:���q7���ٛ#$|���lJ�v%X8%Ð'�32���W�*�� uk��{�06��� dh��z�h����?	�g����&}P�)�w�>�J�NA����r�羇:c�'_���W�z��b)h;Xw� ��2F��E0�'6�l�@襙��L�]8�T�<�������Lt��/�����F�����uN �	á�`�mw[�OpO�w|U����I�!�N+��Ơz50&c���H
 ۸3} �J����)u��hsy�X��83d�$���c@� ɐ���ߕYr(Fx����L��e^ܡZD:��f����Zyj���� �L2vK�q��������YxWĶOJ[���;IJ���k.X.�a���M`���\��n�<��"���!�;��~�(������v:�x���MA���Se�=A+,Y/�ٞa�|a֋~܉G�7PΔ0|���Q��QV[yU6���AlwP,.���ܭ_�>	 ��� d�I������@�'/�r")���	9�v~��*�,/Dn����0j��o�p��ƾ�{_V�'��a�U�O�K�c;�.@P�y��'�W� �t�L��H��=����M��4j�r��`���rgAG��_��4��Y`���Θ�Py�DT�����Q�R���]�7�P�����[�(�Z�h�<&���6������?1����>&l�l��
:�Ja"
���i,�J�x����j�:e	���v �������o�i�~�RB�]&�W�˖^DPFT8Ӱ�9��ESN�ڷ�'Y��yO7؁�)Ŷ#�$O��g�$���z�[	9~�(���_u%������t��`3�qRq�7�2{�\z�O��\�KPL��X����Dok��а�H.;7o�u�ϧ��?Z��Z��8ߊS4[Q��7�tz�άl$8�L�x/�؍GGr���V���G��csp�z�����T��P��.�Y�PV�{O�U�4�q��er*C5�ZfvN���DSy9j�W :(>`q�A���	�|Z���dR�.�\�*,0�xM�,F|�O������{��*1`����Di��3�� �X��ǀ!��� ��dc���~�;>ԝ�hL�9��C�lMC��O�y�&�Ij+�-�ʒ۪�q㣻��dN������Zgp����&е�b?�ҫv�G_�z1V�!�Wkȧ5��ӵל��S�K�Y�0}N�]�A|�ExQ���n��	t�`p����Q���#,xF���E!�����n=���`�,=�=�p�s�]�_����8l�.#��m�*���<mJ =�/�a���X$�Tw��~�?Bv~�0ՠ�bA���~B,sh�����ؽa�9t8�?�d��B��s���b@6��2�e^���S�j�p�����׳aH
�Z�k�C��*l�Ċ2ſK���}�e`�u�p�~k�;V�MGМ$%���JT���=����'�q
�Y�ß%�N��2����U�ԅkm�5g}�J?�a��6�E{z��J ���⡢�3a(m�0	1T��-0s����	չ:XN1�����J���8��D�s^��	*6��\�.��?��D�.:�X��}�5��.��3F4�H
+*�j��s�O�h��R6�U�f2/R��gr�91'IB���4�@	�_c��~�܉��F_�,�O�5�+��P�C�%d�w�Ty�ܼ�%�fV�uͳgl���p�[���	&���8�@G)Z'��l;���d��Bۻ<���`[v1-O8�:������[ܫB�q *�ʜJ�0�Ţ���/&(*�f%2t�S�S`h�fYA{ə҈��ɱ��ѝ����@ҍ��P�r 7����&}��b�g*yV���KA�pk�g�j#���"!�kY�W �~"ꊕiR��	%)���?oG���ܡ��+L�lE?|�7?�Ҳ��]3`���F�ع�|�<2�3kq�SPH�ĝ�@ޮs��X���� ��k��V�5�Ҭ�k"��(iZ�w|ͣ�_M�!�ċz\}�-�%q׭��N��[��.�p&��y��}�(�'��G�b�@���p���?;���c��`9ߥ}A�lf.�^:��;̓7FrM���7� ���I缔S�lǮU���4@Ӵn�1zKCa�1�I)\89ie��q�vJ��Iˌ*����t��fo��%G���f8��8B��� ��bZ���DE�Q���\��9�heW��{#���� ��{^�,�p�j��,��d٨�-8̛	ۮ���c�j��_�l�5����ۉ?Wl{�D)��9�Tܑ�Yx�,���cP�����;-�w XA�Z�y�/6�6ʘ�&F�C�ԟ�Q�c�߻y&�9F���cu������s��l�jk���2�	&,ST����m�@#O���`���rվ��G$�b|�S��	�fW�<�󓡭BqsC�l�i�l�`����.Qև~g��f�뫶�����h��7z�t�Ԁ�ҥa����=�����|��P2���g��ۧ%��G(ڧ�����3h@c�I>�J1 s��[L@N/���H��
{�����} ����~�'�=uӴ��ۇ�C%�ьѺ�� ���J��
Aqϸ7p$�V�fmN('�=��}��[C6�.�Um��j@�y�/�0`6/�i��&��)�h@���T�H�Ⱥj���G���`^�mM�6��k��U���Gr�P�*��ޱ=k��`4�<�<=�J����p�u%~��Y2~�aP��}�1뀶���Y �$ά�"�ɵ�4?VB �SE��ڧ�Y��g�a�6�G
�~�
Y�iů��O/b8�v�G�Q48��N�/�B���������i	�l�X�N({����
�懅Z��W,MK�_��&� � +�v!#J�P�u󍏦LK�d����(3�VT���R=ʃCŀ�� ��9oH-54jM�@�����3
��訽%i�.��� �7@K�*� ��qL�U��ѩ�X hP���CdӫUg���V��rK��`���O	�S�m��AJx�#�Cl�5��j�;V�#O��8�0JSMC���3W����>����J�h$���/E�ۤH��·ˑ3s�DW,E�y�q���6�����f�����d!���\�.:e�ܔWo�ݒ�!Q�f%42rҤ�|�q�=�_c� b�&&�ㆮ]8�C&IIݠ��ZV�2��KB]��/Ǖ,��#��N� �f]����BC5U��*'<p��@!��G�� ���ͮ�E�G�������+���S��?pk�5��fe�Z�����t5vtk#-�(\7��
�N|��Ae�p�l��?1�l����j��?�/���ùM������+�@G߽6t�����_� )�L��v�}���_G�e?� ���Y�
2(�S<��,V�wM�����t��x�Ўd�G��4�O��w���/>�:��1hF>=������w"!���3��Dv5gdNR�w�wh�B�rkz��[>�@R��Xc�,2�:�%Ls�*�b�'T�R���Z���5��h�t\�ҕ�L��D��j��F�	L�1�/�֠��r�S�!r�<i]��>�B2�9�$�Zd���ɽ�T_/�����@'x)�㔢�9�	���q�7���4$sYmy�TؽZa���#A�L���y��@�*�09Pi兘���ɐ�_5F*^�5���T^u�*b�?%�V�6Gly``+��烆���At��5���W���ѫ�O�
��c��q���_������S�����=ո���+a���S����!g_��lRʚ��Gv �cy�센_��g��dn[��En�"��qE{�wZ�F3N؁��7���)NF�=�����ꖆ�r��n�I�YΔx�}��-�Ձ���� �F��*?�=j��V�����z@P������H�6-\N|qX�t	�k��r)F*٪v�I���I6�jlZ&
�����F���=��n�/Ep���)�b��A茒�y�%S��7���f��I1���J*fl���A��G�PV�y�RZ��Ƽ�A��Ӿ] r��X�υ�_?�vAM�iKd·���W�3�jc�CN���-��_�c�uD���#���������%b�~��J�g��p���$Ǎhxx��f}Q9T�^�V�m����9����0�^#OǨ3+�pV�c��&~A�=Wy\������q��+LS7���~�������W��O����P*D��+ $Z�{��%�A5	�o�5�F�� �uN�Ӗ�U�Ź"��x��vUwg,�WBf9���ܛ�/�Վ��d>.�b�w��7$	��h�ϖ`�M�r>xB���)��<q�.irsX�O��ʹȘ�0��2n��u�El�@���D�&��<?�
Xў3�y�\R?�;z*So�<��\׍?|��=�ӜB�6�\�d��d�7)Ϣ�A� bV��걜-�C9�O-Gcq��mW�R�9 �;��:[�`Z��k������5��m��#(�"�ҧ:Ȃk<��@��`�����R�a_�|+����,n�^&|z(�%��i������R�'��5 />LKQ�ޘ�Xޤ-'�����æk��q?D���� �l�\s4����P9�^nz(�Xu���I�� ��g��#'��d���Գ$�G�]�x����GS LX	�E�5�M�@vUp<0\�e�'%����V^:D0ћ楣r���^����G&�;t������%$�b|P�;HϏ�� %xM �OT�ts��%���͹��ߺE�`��s����|c[�)���}4���iF��KY�s{(���U3��l��^�^�16B#�@�y��m�&}��!����!�!Dd*h��pj.
���>����� `�4;����q=�� �3[�]�u��(��{t��1���I=�:�bdH�م��]fT<u��pli���0*`q=m>eR��(��:���h�3u�I�@SF`���`�r���l"���k�! 2�hxh��!
��qs��	��X�j��ж�����`V����p������J��OYŎ8�ő�WF)�|��������`A��k1���3H���ܔ�$���wӽ}����`�c߂��蠕�yE��i�	�̏8���c:MT�PJ/�+�S#����Jc8�Q�`4�O�Y'�c�N$0W����D�$�I�^��aHtQ
�U]|�+�V�I��S�I�#^*rUi��:�WD�&�$y�@a�EP�~0����~?m��ds�����Y9*˔�k՜,�(r�9dCɗ�{�����@Ŷ��\G2�]W���3��<R����m�wх�Ό��R`�|]/?��s��B��K��J����"n����6�q���������y��zM�\��ťu���Mn�� �]٥���P7~�7��$��^|��ا��`1��a����'E��Cɘ����-p�j�<e4dR2��Yo�K���3����1���4.�Xt�臥l
K���
���֮ཕ�'JS�h�n��T��د,P�� �ss�Z$�1xK�q� 8n�H�π���<�Z���-�"��^F��6@-�%YH�}�q0���h�l��p1�8D���y�3��okψ�!�)�ɀ�`�1l!q�@'����y�=��_�J��$8����T�JVP��e�bwh3GiD���I���F��t��b}�
�7=<i�Y@{�o���J��gש����h����`sz�8�Z�V��-��|
P_��Ly�D���z3m��/�'tIπ��-�y�wHA� ��Ha#�[�*�� �ڏZ�=�c����=`�[�HL��np�����B�X����{!�z�O��0���#��\
��ōZ���>��Y@��w�T���.GT�!�H;�ڰ�4�<��/�a~3����7�O�v����Æ�V�
��J�v��I�s�L;���v?���C����֝�(D�{�X�������ܲ��s��v:��b�D��zM�K��+��:�U��5����2���|��	�xꨉiKhc�D%e��S4�tyl�FH
�.lS��M�#� $y-~�g6�EJ���~�f��$���/j;r2��)�:ZBϣ�h�ǐy�%��p�,�/��
�F�
.���KR�ѡ����3"�^���;���-焽��O{���3z���	Rw
Es�H�}�xl�6	˓N�Ra�H�"Y\��h�f��&^l�ێP7�s�O�`��y�� ��-�~�z/�37��<CW��Z&̱ݘ��r���	�����NPqb���Q���^�VlF��w��s��(��eI���!.���KeIc�w(H@K�x8ߐM�b��a�����e���s�w 㛢�OӮ�N��;��8��x���R�h��1��:&�/�*��H���o*�j8���1�7CE���*�V�>�]qv���Ï,��['�b��K��Ū��H�O_��u����f�3[mqI����j�W�EOzx��?EȬ����Ie8��E��_p��!ܡˡ����P�L����q �D`S�'a�Wt�ڰA� PY��u�	��jkv�ĵ�T�f�f�Fs"�6bf�7����N�H̃<��:i:L����6�4FĨ�j=petx�CF���E��V
�9l��=|�s#�W#[�E����G�����qf9�N��ݯ��h�
�6��r����,�-�qP���&�Ʃ٨�e$�p���@fM;[q���g��)�?,<��ד�r�9��>���d8�����T�J�*7���8ɛ�*��)c��� d/�ȋS2�a��}����R`�܏�34#J����^���#��99>��>&Y�4C�*��8�W�!�p�T5^^���3&VR{�����g@V�����5����f�]Cx证��v��������c�G�9ϖ!�BwJ��>��t6��M��UnQ��ڍ+�ʬ@c-��ђa�ǧz�������SH��t�`�~��R"�暙�R�3V�� ����k5��8�E3�� *�ʣ�����*1���<����^�6]�jk�EӡmW�O�����<�����Ë�颿I�8����7�:k��C�G�B�G��c����Gf����
�U����ey�0�)��G�d�7���$�[�����.6l 񎭕�b�5t���.����yS_���>鞓o�*-�|������1]!�k��;�_����b�/ *5�X��sW�l�z�#6�����B�z�O[CUd�~��/�J��I����5<��9�F�^s���:H�
4jA"��s�6�$���3ͳ�ģ�c������8f��ݢ�o4_����T
��^l�hTjQp~�i����w�F)�XN��9Y�W�����4,/�{3��=���#%�hy[��R}��8�_[; ��eMEc@J����T8��}� ��@νȼĠ�1�HX��׎�Z�u�>�c���9ΤR0�=���
6{��ƽY�mtY��UF4W*�)����$���(n�W��oD��/��lmAG��x�4�{�$�%�a��v�UQ��F�����#���ϭ�i��Ӌ+�AR���x�̸MS�gl��:i�ƩnV ijmm�P�|z�ˑ�Z)��e�y��3L7{yA@�vNx�BS߻�L#ͼB1��
m�0���ѝξ�܄mQ#,^ѫ��5�d-����u!�r�\�"��Rm��8p�� �.�ķ��n���ˤ<:a���MP*�6�v��FٽI��8�	�E�� K����uYto���L=��G�E�	�7�exQ�'z�[�)��=�k�\/Kկ`hݲkѽS�k�6�*�?a������U�Pگ�S�S-�+���+0.�Fz3�Nt��bΑ�� ~���d��J���F���8Iz5�O��x�Fs�!bY���AO�R�}[]����g�2[�r&>,�k�H8���_��gwN����eƓ��6��u�^6҃�8�=��
sd�@���g���$w�RX�2�N��[Z��+�0s�p~�`���c�� �u��I��I���z}��Ө��RظM�Wgs���a��5�_�S	�s����7�n�c����\���dW�����n�e�� �]�hݞ8wF �Y�ɰ)�jܠ\,1uR�]��ME�A��3M9T�00��EP���?��(J�U�	|�o��kȚCh�J��'!��_��+��D��� ���|%��3�9\��_�M��y����/��.�f�n�B3�v�ꗉ�st�f� oͥ�=��y������I����H,VL���qP� �Zg'i��$��r�3�ae�%��;E�┩�(�6ȃG&�6�pv ;dH/��>Ǝ3�����ӽ)*E�.b��"�R�6���Hl�����w��;�[����45!�ip��*+�D��Ef�?rC�+uz�籁��+�v'�Gh��>�l��7��TN�}���5���f���9�� �*���q#4}��"i��J5"��#e 7�C�����\a�{}QE%����5�za���1�>\;)��쩅p(�b����>�����'�(ʛ&iY��V�YT3|�yҪ?�/��K�t�&	�V;���u)�,{#(�}Eו	M�;�MB�W�
s׎���ā£.�4���xG��U�N{�U� ��㶩�t�Rز:�Ê�������)�Tb�������Z�(7��J.���m-;�%x�Y�|+2:����LՉ��_�T-��7U��^b<�(R,6N�����ݞ��UX$-�@`�o���uV��?h탬b�~��a�}$�>`��`9�~��گu�'�dai�>oJz�V��dC�F��`ו7��M�P3��K8AWq��
X���@����ƛGLl�_�a+С=^g�9}H(;�h�o�}���BYF�E�k����Vm��j�����rdt��%��JH����~��s�T6�e�!��j#j�Jt�1 8��m�
�)�NY��N�
հ�멎Ž!ǼW
���@D���	I�z��"�%{��I�r�S���{m�����{���~��J⻌���S�yj0H53��g���S���#����2�7�5Q^=7=�%�;X�3u��p�z�D�a�����W��t�!4t����T4��h቟B}a7�b�i�����*'%hD�I�׳�`�á#�|�X���EVH��
��h؅�~^�<¾��8��ж���][kh  ����!2<"�*ٖ�QU�KQ,���;����vQ[*#<N+2�-�e�To�2�X�A��e��v���,����L4�()����̉�a��ޙ�H'�[֜�s���@��F�x���+O�����G��\J����'m&XO����p;��/X�X��l�E�nɅ@n���Gbz����t�w����{�Ç�u	P�c�UoH �)�h���_��v_^���a�$l�] e�^�Ƶ�umh����D��^U���;'%Q�I���DˈK	�8����9kP�#J��9���Ю�"cf��yR�sl������� �����jP� �Z?�㟰c�F���;?^�8�@����;vƅ�?����7���I��׻�ni�2�Sm�{��5J��}ۤ`?�d�ל���5cO�F�S��ڪ�ٳD{�޾W�6=*� �SJMX{9��g�����9�_��{�9)g��bC�ce�$��=7څ �cs�Px�d1� KhG�|S��Rǖ�~��z��ގ����q�.�7����7��]���l�Q�E�)3u��B!�Pp=����Ǚ*j�<.�:ڼT�G�܄��1��Ⱦ����8Oc	1�/|W����L��o�^:Gp��t�"��TB�c���]3c�/iS^�<������"m��'�q�&�%v,�����J��Ţ/Cڲ=������
OQ�t%$�=��[�%/&�V6��W=G��$���#%p�#�Б�����S,�Y#.C3F�?J��l�6e�G�������f��ך�эƆ#�_e~.���i�p�E�'����5wT�5`:8
�લX@`��Q�L�w�mq����4�(ch�qC�9XWxt�7�~�1WM��R6���g�9K.��.Y �|�I�PjÕ"kq��>�pb�d ��0ky|�eۅ�{A���Ѻ�:�tG�Rq�f9� ��ܶ���Fs,4�l����{�óx�!m�f,)9}�%x��2������	�k�X=e☜%�8����Ԍ�0�o�m���T��!�}�'���{��=�(���46�^x����eQo���7���O�e�E0Z[���d�Q�����E����KѹR�p5L@�N	ƻ6���X��>L ��/��Ɯ�l���7��g�h�Ys���c�(0�#fr"�*�+�)#�e�j����vUj���q��c���V�9��� �.�Xs\г����
�FM]3z:k���w��x;�V���d�&����y�����#��@�w���x�x�V<�H�;���Zx�&r���?<~�����v�N~��dp�� �cdz�Mw����k�}�N���@�^x� �ĭ��-#��İ}D�ʺI���఼|�j��I�5Έ��a�����g�}�p�ȗ ,2S�a��[�*�=Bn�.��-Z���ݡ:��'�G(��˱P7G�7[��p&%Včt���O��g� N�-��A>�����jA������m��z��v:h�W�����CG�6U���ƃF=Ӡ��ic�ɕ��m爊M��*/�[�40�v`ʼ�S������DH֊��Z��T��Lt�<����4� ì���t��x3p���Eւ�>B<�q���)J���Ŋ�yYC!T��)ᕻ0��J�#�p� ic��Z�g��B���������,�5�-�������J��*��\U��k������E��i���q���#YU����I�t�������-Ǝ��)��ƇQ��-]|4���Y-~���aZq1ww��ՎjvwƑ,��^��9x�[G���2uK�1#ތ�-�m�{U����H��_Fik�Z����%��'K�h���'���ʨ�\Y�M��0&��7��p ��V�����k�\�� Uڧ�4��<�h~/f%�ʻf�a;o.R`("{V�j���*�Ц��<�����5��F�D��!Ńab�sG�uy�� c���0�Y�� �&ykTV�wǉ]��ۄvkl��2R�5:@�u�]ßdܭ���2�_zRm�I/�����^�Xz^��
�R����`��i�j�k��m:١M�iÔ���ҫ!�_Ʋ��Q�B-�>ɿ�0��������^�G`�8��}���ZTa��m$�6�����R;;��ܨ�=`���1�<v��/pllЇ,� 9d�yv�,}�E&!h^�"	g�mr�V�Sj�;��Ƹ4�<�b9����LN�U�2��Sp�CC۱%�H_�.�� y�5[4�2�)*81?<!���8s�����0C���?n��&S��IJE�๰V���!������J�mJ�V���e�3���b�ӯ:�;�O#tߕf�)M��8�
[I^B�2D�"�\��J(���q�����oF�=C&���h���.�$r�\B���і�c/��6]̎Ue�f>���= �.0*�Gѹg���E�^���N��`���uɔ!��6���"<d�!���u�����,TzQ ~Tu	¥dJ�k%+�}�$�Hd�Gi��{  #��dw ��SwLj���)Ϝ~�QO<F�=��Mki�w�ۉm����
�=V��$P�e��g
e�(�Dγ�:��im�鵮ohK�cQ�E�9M�Pe�r��6M���>�#����<1����E�?L��Θ
�GC�7=���K%�����Ǹ�RZ�~�zR��fǃ��f?�l���u�(o��BJ<>���/�=W�#���A�H+����F�LT��xO��R��.�,°OhMgg����GE{i��N���}�9��@BR�-0�}�����>�_�Zu��璱�#�$Ғ����&_�+}�l5�qv	��P2�Y����i�ݰ%�F���Q���I~VTj�[���b���0�,w?�����zw�Ju�g��ɤ-L֤S��3��}��yG��tS��-F.Z��-Tt��"u�x��Լxg�� F|�#���	z���w���P���=()p�*�JK|�+j��3�{��?�W��g7|��UM�L��M�ĤQ`����xW���u�p4����}\��"��_�\��ͩ���������PM�񢚫~ߕ��~�_J��IЅv�Rr���Ua�����A;�ˎ ���?�}3�q�LH�P^X��u)�p ���ܿ+�Y&��|����s��	�z1�.lla�~�D�����F`�]�C��/�?+!�0D��,�iƹz�vI�w�_Otp��о`��!ߣ�D���O)eH�)k3�Θ�T��W���������ksc�m�D�w�gݯ���S�s�����1������l��[x�re�%��=Az���S�c{k��8�������:|�O�#�Sc�L�q��"������h	)�F���Yc1�&�& C&���j�hV�o�Z�RXۓc�*O�~	�,P̕�3&�rqFm���<��1
�!d	\o1��\o��I3ΰ��M.��H����@2j��s3�� ��:I��9��Z�4SB��>��{��,�=Gt8@ejOsP�;�@r�lޮEM%�4��4[�lqJ�S����J.���j���@5��p(a,��Q���W�>#f�J����9���)_��5�[�s'����5���<�c.t��l:��������a���xjNpYS�<:��
,o��s�`�g��;�|~N��JK,�����s5	������%�V�ikXV����������i���~�M�����M(�R��%	K�,C*x�F��$�*�Jt���^��	zO�F{��lŎR_�ABʋ���2�5�=l#C���U)f�2k�C���/��R`�#��^��I"�tc��$M�ueP
Hw������Y�uX����O~.h�U8��G f��+VfMxj���>��Ac8�9��̞�>8Ɨ\�{�5A�? ��⏫#q#� ���T�J�P�U,�����ydC9$��Wp~A����z!��\Λ']�U���DEsM8}*�!���	:ˤ�.�O/SfU��}��&~�c��<]��C�(!Qq�t�7՘'�����.��(g�Y�4> �s{I���L'J�������� }�~̍��]r��U�S���T'�pE�$�q۴����F���s��Z�M�1a&�j�j3Z#r_�Ł�c�$�vV����"����-����$������ylr���8!RF璮�c-�-���h����\��d*÷�s����N$��JVfGJ$� �8��+{AtL8ՓJ��g�v&�xZ�m���̥���h���1|s)�:X�Y΅�3��hei{����OM�5�{[tRl-��i�נ��[������#R��Q�-`���95�u��]~�A��\p�E�������J�"�!��ۋ1 aa������a��A[
�AZ2&��dև�1)w9�� ���g�ZX��jw��aJ}�ŎL��9�~���%ɟ���.:���I�NK�|��[[y�I4OR\NL���5Ʋ�sh�`��������h2YQI�¶�U�m���OǏ�&��=н�¨qZ`A� #��g��s�WY
|�J�*��!B�� �p^�CG6���'#�{Z*@�ڄŘ{bf�G��f���&��\�=�/�� ⟍���p�����\��͹��xu���O,ݺ�ʏH�C�J���.�E*�!����)'c�G�ɲ��د��E�edT˭iw#)7��yM"��#(<^����X6�}ph�$� ��6X��#��=ypX!�����U{�ȹ�G���}�2�k��ڳ�9���3���P����q�> x�Y���a�)[�~oZ�'p���5k
w�%:+Xn�0H_�)�$C�;�M�ٸ� LR�����.3ȟ�K���!�`��mqc��D�aR�����6CϤI�`�ʩx��SV]�jZ��XzW�[S*eXp˷�
����'S
�v�zi�&;���T�a��6O'|��b��3�d
�~T$;��~|D���#�r��&ǋ`/�|S�`낶,L�dĊ���h��l�A���Nݱ#��|��?����V�Q.�/<�����6;����r߱>sp�S`�z%25����p9��%���ŠQ�x՝op��&��`@޴ |Ψ�z��3���%�k��g�����?
��O���zm.��ko���
�K��3�lSy�Ѳ��z��H ��)�V��}@�v^7ѕm���#N�[H��>�a-�P(��
X>���;O�Q���o$
c��y���D�1�+F^~�g�Q>� \��[��O�0�\��[�uΔŊ�\K�'�a$W�����z��ڠ��>�]׈&D3���:�4��+]	^��ܧ6�18J̈́@y�%4k��R�u�@��#��=�)��E�o���t"^�,�avp�2dfyZc�ذ?��aK-b�pu��:�,��*��7�D��	#�y#����`�@c�
i^��3��0( N���$72u�+Љ�ЦM�_�8[�<}=��ͥvI�qn�z 㡾7�e ��2��CyS|-sE���87�@B�\p�2��Z��n	잃j�����yZK�����X��!�Ԙ2e��J;��;T��4�褎��5
��{x^bz���:,}˻�YO�� �׸l3tK7j|��ǁ���D�3��襔u�\�*Ol��6>���f�b�5:��'0k��`�����W���كx/k�mI���#Ō`i=������@W�����%*��]������$Uz���L��5r"(E�f��=��\Mp8)���'ޠ�*���lT�Ǟe�>ڸy�an�3�.(Ϸ%�T4=�ҷ�q�����@�DФ����p`ݻF�zS,L�5s�^���[i^���J;䎰���7fsjk���2�*�'O���O��?�I-Rv�稢;l�v_��H�Չ*�X 2�<� �M\3�;�Q�K�lB�*[�ӋT�r�����oI�<M#|���-&ʓ+B��:�H�Q��f�I6a%/V�N ��w�~E�*�ʅ��Ѓ(��$�!%d]ar;�A5V�V�u�Ҍ���ߋ� vj��� V���g9���l��+��u�s{�\��u �3�Kۊ�z'���椳�'O
����������� ���Nh�m��@�Z�S:�q��c�b�%����2[�[*9�T|be�m��}�h�� +΁_��I�c}E�O�m��:��r�,Es�Eg��}��phE�e�ϳg ��%��5�}��d����T��
�`����ϨL;��p���V������N���f�Y01ٓ�\���:�o`�p�X�_�z�v��~03��ҸO3����Bx^��cY�h�XBߵs�ٺ�Ն�i/�뾪�������<�(e�zd�D�D2nF-�)R�h�A��;$d���Ď�`XJO�����0OSA���t����%jkZB��f�Ms]�+��r�'s}@�`;.���"������.W6�=H�{�ŭ��	��C�d(���4���#�f���p��I4���c#�_Iz���ٚ+n�T\�SS͎n���*�I����� �(a��U*[+c1��F�(� E�P(�#jB��a��P���3�Քr�z��a�q
FJ��#$�AG"2��^B+f2����:y�K�V��w��ep��� �"=1���=J�T��U��r��w���Z3u��\A�$��T#$���4���]��L�d���418�A��do�����a��󡁝DeQxJ��F52��S�5n��~��I�WJl�S�>~�[�j�9l5^�]c+��er�<
�x���@�H�#��	�'ڎ����zd��ub�:JWI<__ \���X|�ߧ�A�@��Ƙ)�y�Y9�S� ��Q����	I�ٽ��A���+{xE��b^mW�D�5�&�E��3
��闗���R���7bD��d�ٶV_�GJ*N�W���I���ř&xJ$�w0L:�� �!ЈM2��w�$��l�䁓���+���h0�{5��ģD��VX
�I�0��	�u(�%Ƿ��t�l���
��B$ZԖ��q@GI��������~��݇K|5��m ��d3iU�t�Gyҕ��2���S��D��n%�{�|8�:'v�[�ESgx�+�.+Y�6OX�^���:���z�L4N�uČ��1�f2�~C@YMB���0�<���N��n ������G��b=�B�B��!���w���!�Uz�� �é�@׏{X��b�7�����W]a��<�w��>�k1)T������;�/�t���t�;{�s���yL��.J*�v:���������J���{#Е��,�|��:�ʙ����� �� ��,A�"��{���/��ߜs�C�4�f��?F+ޙ���`�R���#���8�z�ܺi�߂+��n%#����Ż�"C����lq���P�/�����P�}/b͞���
	 ��Ɩ��G�cL�{��rmˑ��E�W&I"�N��:���'O���Y����lFU��x�7@_$�BY�U����^Jn���2o��+*���K�!���v{��-��q�wT>��Y�*֍ykb����̟m�Z��8Yz%4��2c�ү"����x��ȷ�!��׏p9CoIF����p���p߉��,8���mg���j�{sn�%�#�U[��U���u�%-����Q{��7]�����E�\��0���0���u&��R��Ɍ�ﾎJw�d3M�[��·Lji��hvT�E�Vy/~x	4'� 5�D����b���T�4�WT��j�EM�M?���[�N�!'���%���^̥
�\�j����<���]5��J9��ҳSʺ|�<^��U���*��o��z�c֐?�Ф!���G���'Vq}
�7�G6�a�<.L�E�bݴ@��ۧ�J��ҡ��QgR9*�F�Jj�";�q��L�N/'O�kZ4i)�2D?P��Kp9B}��鞋$HE�|��09 ��H���[
��'�ق"����-���&8����6�J�����Ȉ�����I3��5[�1���X����|N��`5g.b�p Qy��w�x��Ǟv��@����3�ڥW�B��k�OZW���s��o8{m:�%�Y ���N��/�a�AY|���U#7��[z�U�Q*԰r�r���� t�K��z�:�����+�B�`b_��;54z���s>��_�m��I<�	uZ���SΚ�B������"��;��Q�M}T�?�#��r���_��3Ohjx&}ж�=��!��U�西V� +������kЕ��1�G"\�}#B.ǅ�Pi��.�h�|ղD��6u�y+��a�J�M(K�{�qE<k���]sŒ�wG�{B3���5���(��M�iRb�[�!�L }�;QSd��='Y�C�J�2����<8o��K�mY��r<ʼ~왔�	��W�Eikv�Qv_Ό3����{�`����9�H>�O�}q��#�����-�\Ń#���)�OO-I�}���0$��T�_��[��R<{��R��\8ސs��wL�R��r��)��5ߒ�(�;[����o����7k}��LT��u:��b_�.���!螱�|�%������� ��:���l[���Y5<_o
Rl�ؤ�5 �����_�ೋ^;:��#��t��y�i]	jшX�ϓ�Rs����P3:�PV������7��XV��K��A��+!��9�����jE�P��Z�������VX�-���(����U��2�� ���8|��T%/8_�d3k����$ם��{���[Q-�9���G#��/{���N����[A��R�uIv?�~qH�Xk3�I\�l�v~n�|�	xT���0j?4�/�&M��R��Z�8��]� G�Q�|r���-7��D��8���;�m�~:
��x�4&)�6���B>��SX9P���*r[�RC	�Mɖf�)�x:��n�~Z�L6f��r~���д���)����&3�!G�&�� ��m/��gx������5�P=Y`�7�N�b� ,��ۼVtpJ)����9R�U[��3Ч@|=Rh��¯N�Mյ�X�q�@V��hB_l���m���{�5�
8?|p�s��:���-�U�Y4�<�O<~Y��=�3��k�ݨ���-����!v
��Q�>�6׌y�[d��FB���3L���̱����/=���vB�v�S۔%�ֳ��ΑYni٦�����a��+�(jJ_��`�)͙!j5 �N��N���V/���M�ׯR��4�Ya��G�"[�~l�e�l�-�a�	�"I��;�Z��{��[2TIȠd�+�5�=�L��5MAF�]����cXF!v�R���ٷo��x�M;���n�־D�����������o�7v�z�t�WT]y�N7w��'�(�4f���A;X|AN*"��1����m:g��~6'�CQ�@I��(��ItW��&W,ç�KN��!G��w����$�>��jp"DfPi���١��9}�'�T�Y<�nU�yF��˜Z����!��)�F����B���;�@SX�ˆ�w+PB{	AX`,�R�������*�)�R��#�i�8���Dl��z���5L��#�����zK�&���1Au&�5�±���Ph@��DW}��2��D��<1�rP6U��[,	��1��V�Ӏ2wI�+E��{�*;��¯�yoq��4jT��H�$`�>j~�H��Jǆ��b��_n�NEy(2k�1j��:�����*혛� �o��cQ��}��(s�W�
��L�1�}Gvd40�,Ts����q� e�#���԰�2�r���7hV�sk�����M¯�	d�(�i�E�⟔r4�R+�7��n?G�S�`8���J�S�	���Bi�k�s/!��-9��~�:���]�l7�/~Ƨ�R��T�c�8�/�U�6�4�,;�(r�q0��63���f�o����˞(eOE�$g��w�t)�T�ݢ�b��8E�{��w
��d�#SG2{N �4uj��#)��G������̥/�ch�ʁocU�7oӐw�dsb�([���&C�.\�~Wtڣ����XP8~���S>>�5�q7�i�	O�^K�E�+�wq�C޷ʔ?Ik�<V���;��$�A,F��	���*�1t7I<<��&�/qZ�������~�%ͦ�]��ڋ�\�JFh��h�'Q:��������e�|�T����=�|���G�T����Ko���b��<�:
��I�M1�'f(�~�.rD�y1�H�K���W:ȥt�J4�N�\Fќ���*B�Q���S���!�Fo��+��d��m�|���ʔ,���?�X�1��K�b�����:���縱T��I��@��K�/d�_Y�����!���|B�V�k�B������g�7�!2��/k(�����ߏq'b2Aܐh�3NՅfge��X`UK�
}�ᾂVZ��dğm�|l����q�	��Q_�����D�)�:˘��gS����ۑ�>|ZP��?�=I@���ޒ�V�I1��Y��8U-����A� ���D�F<y��ENQ8)����s���*��� 3�k�W�#/ �LK����<c@�>"�	��v��~\��=����z-���dJ�{�.������#L��q��&>04�8=9L��ꋢ
��>��1���$�7"�t�MF���P�����L�G)e�-�#�d�3Т�m��7�!Rg��LK����+q��I�"�O���x�����R}�u�=��F�I�ToS���m�!sl"ʹ��"b
�L�[���íyW��Aҽ)����NK!�B�"V8�݀tqqb�*�x�)w�1�M�A�RcŖ?|��
���0O�"n?�z�؁�)�X��H�i_��
�*,�]_��c4Mnz����H�5x�1�Vz��85�V
������gՙ�H/�r�S�_> �\�V��&�.Ɋ���t�ًƲXdj��\�n��(�]��쥤� o?�Ù�[�^H�+����C�RHͮ�3�V;�X�k�(.��ZjUjU�K�}��F��/�z=���t��5�[�Vcfz���W�ͳ�%���U��[�4���`���裩x+���5U2DC*G~���~�s\�{�?�\Q�o������r~�6��� ��������P���kMxI�b�C͠�����4�����_	�8��ﺤe�3e�j>�`G7�a:���OSo ��ǣ^k/@�,��|d�����3��g��>,�V�/6� K�L��HO�>=�e�/uZ�y��9�m�"�X���1_� C ��D�-��ޓ0X����y,�l��ZG�r	D��%�[��4H`�K�N1Jv�}|1㸘��$�P�YbRڃ	p�E�7���۪[�8�s���]�o�J+���Dg7�h6��P�}��a��L����ƱN���O"�^�+��G��v��pr+F�N&��9L�lBb�����h��v��q�vE*�����'���=1/�ذY�4�w�����D���z�'2��fY �l$������D�°I2g��K�ζ�$� ���Mxd��H�!go�g��ſ�0s/��C�`ȼ�u�$���2 �Z�����2��n�k���2b�1�Wx12�	z��o�b����,��M�i��،X�2c|��!�$��AK3�ZS8y=���L� ɓ8���� o�'�N�ԪS���h��S�����t#��"�j\�p1���2X��$�D�핫pWʭuJ��殴V�za���Xa�>�CΊ�,xm�Wfc��BY�8	�k=��6��.zU��7���Co��:�+g���nB�/�Gh����'���Y�sUc$\�r�=�%��!�3�Z�U�Ba�Bn��j  ���Q�e���	�,]�ܙ��ZC2������V_l���a&�
mҮ1��%�	������2i�8�����R\�y��oW_ԊL�rd�»	�����t�L �w�¥�̃�(�^�(�jJ�$m6�$�\=��1_�ڸ
$��2�S�!+��Kcy	|;fIU��Q(㐁^ٮvi��lQ.�|��4��i8\�����*jēw�N��I�b	�Q�괶��!Q��f�f����|���}��	�)s���1�p*��d�^ŋzv�6M����i9Vbo���z>�߬=f� ?�
Ĭ!��џ��k����g|�e ��sauF�;��α�v�V@e�E�4p�⧐�U2�Hn���J���Z��y֑��[�o�᧪fU�і»L�	\�t�,vKc����S��#G(��U��r�j�\w~\��X�*i���w�9��'D��E^�Y����t��h��%�|$Q��N�6x�����2���㹑F�d�����Ͻ£�7q��{���������K�pJ��>u~�ݻ5�w�8?"x�N�K������}h\ғ�v+1 �z��%@e�eވT�Z>�\�IFv�����e���ܽ/��^�D��~�S(<�'�mӾ�D�v�����@�I�g�|W8]������T���*VW�^:�ɪ2;Y�{��Hx�N$]��ԋ�&�⻳���y�T�~����Je�m�Փ���ZA��~(A}��YwƗe�\^�U�wo��(�3���+�Ļ-�n��A��7:�n(�6�����(UW�6yt؃��(K�z��
��^*�W7P�2��s��^&g�������B�I�0p���&�����S��H+�M��������-�G��a���O�#R2.��=�^>��ݘ�
�+l�;���̩}���<&w�Z�|$ұ@زɢ>Fї�U�a��=��˺�_�����p�Y�cYvI\�k�W�[�IkT��]�>b��ʲ�R��_��\M�?���uXt��'E���A�5�d�">�&�/mJ�CZ�WEgBHN/&������ �oȥ���Vcٲ�]Q*��UCo����W.I�� C�؞�^z=�U �OO��7�6C�L���\W
��14��+#��~�0�?<߀YзB/W�Ϥ�Ѷ�F��+3Dd5��	�!�y�TB��q�mQ!�	�,��f��|�L�i�|�Yj�ݩ��,����L��2)���e����6�#Q�!աS1N�����Fuo���Xܖλ�s3��ԟ��蓧e����°$�|ݤ�7����i�,���[]�N9>d��Mz��'�K�V����H���6�UI�	�`o��u���t��;�/�"�l"�wo��E��(��mZ`#�3���B�5I�"y���X ���w��F]9��c	2 � rSW�դ��˃m>8���s�X��,��$w7��S�8p|�Z�}rq�1�/�.�#QH��jB���-'_�eP�}a3��~b���!��i.�dGy������u�%����2ᥑ`�N'ĈJ�g�u�Mw�{�
{�P��L�����1#�^��c�^��Wdܳ��5��t^ųf^�i��!�Zy`>X5���nYQ��݇���=?)_�#}m��S��*Z�y:�3��lm���V�$ś+�q#�
\��9�:�i�}^�痊ƕQ/�wL�߿L��7��9����*�xV�=��z-&���CW�4˻�?�b%X�ھ�տ�;�p�r��ٓDsո9���T�v-Xwl_��ɜr'��^j>���뵍y�Þ}�o��QZA�Ξ�?
M@������G���Rq8� ;x��C��	:�a>K�_t���(�ZV�{ktY��&@bO.� ����~����s�Γb��6Xm0i��6R�=/PS�y<�c���?m���M��#6!N6�1�J��\K�.�ki�V��Ov<�$�o���-�83jX�8��,U}�p˷��&�I�����U%}�p��������xɩ�`0(y	�A.R������(>���Ĩm���6��C�M�S�i4z���`0Y����~�J&��=RrN3'�-(�[�S����B��&v7������d�q
�b��،��na(I��e���ź�w4��E��7��k���pT�J�x�?������p�|I<>MtD#W�sp҉Lʍv��V=�}n�%�v�ݰ.��W�|��L�yy��I�������� ���3�F��zp8�)1� X P��LWsϱ�JH�^��e0:�=��JE��c����W������9zĈD���Un�fkٟ�r� H'b`I�!�w�Dx,��Y�(W}d��>����Q�4�!�7̔��R�DV8������Q7���8�\~z)��rEW�Ċ�^ܥ��7��k����[�-��X��+����_�V�hz�Z�S��lm�����i��F�FT���R"uq�K _�(���]R��>��Y�+�8�H��4=L��؄��R�ZP�Pv��#����y��波bLv�^/=��e�A��\΢�o��T87���T^h@B��8}Vk3ob.`�e{l�gmg9�Y��
��t�U�i�K4~�g >܅L����"�Ec#KW��8��%_=7�;�B�"vX.��8�U��듾@(��T\ ��W'"N�
>��������
�J�qj? �JW��J�#�D�N.��Cr�d9e:�ϪpL}�
s�����{{+$�����Ǟ9�|�O ʨ�W��:���;�Ә9�S�c��ǎi�d~�&M^JdƖ}�-Ǿ��魞3j�75�`N7���F=���{��b�Q�X�9g�tRӈqjE���k�{<��{�-c��E$��H����r,���aX;c�Ag{z"�5���u���X�af�h%��/�Z�>\�Yn�>�ނ+^9���� ���to�a�O^&�Fg}���Jam�ıMuh���Zob�hͺ��=���eH��lF;��o�H��;o�d��O�#W(c��3с`f�*H��4�Ru�m���x��.)DD�B�/�N4�o��?�J������kO7�뮫�	��H�:���mك��/:'Jv�wu�1ÉG��e�"k;��D�nw��k�]���o̞!�HW�}�5.���/�wPs#�R����f���� ȓ������A���\=;�}�j�ʃ��V_�j��bO_��P#��'e�_ ��c�ȫ�0��l!��qҌ��9�z���=�cû�#j"ޗgC{��Z���a�4q�� �p�a���*Dbm?����߮I�!A�r�Ȳ�y��]B�̞zר�7�qz��<;y=��JA��V�C�M�;4=�?��)*�#�:�̥O��Ū�%j�����CP,.K|�f��QF3��AD'Bt�Y=�V3�XS;c�o�����Q����Y��S���J���˓���;
-%�1�����4�V��`�Ͻ�	)���.��̳���Au�ZNEh���<R�4�`�mQR�Gɖ�ږ?�
���)	���ދ��L'�\�R�]�ȵ�����8��$�,�p~���
5����CX���1�K�a�![<��wiب��m�7a�kI>sW���sK�%��q:-6PRd�������;�D�����HrB����Jz�m�E�y��ojL��7>RgkuH^��Q�.:��pm>�cX�EA�� �<��.��=X$�F�^���%��WHP�o(����������~hܐu5�Xޖ�bO���K��0�&8��;�Yo�4���<Bp�>`�Ib��z�į�51�<��^���8�r��XR���V������FAw���}܌w�(�&�Ͳ�h��57	H��-N�̔9���L�i�9�k�8�!�91��ilg$nw$�@#�n�f$(	������(Vb�\�m��H��7^��צ�K�,ѣ�}��픀�A5����)��? �FN����U�4��8$ifV������|FL,�^	��0.��5,�\�����C�z �����w�dJu	]�)�w�L���M�24��a?2��	|�4M8)���x��˰���lk ��R �jAM��/J�� E�2��g�R�p�7!ˉ4��Jj~ҕ���G��^[�A���1N���#��L��H1�U���:4��4��@ ����v����������IHR�H�M���N+<4#Ao`��������S�3��{������`q�ù�?=߃�h����������T� �h�W�H��?�x�g�+�-��W�� ��#�EY3�j�@����[����)��NXj����3F��ۿ��,�¯��]�Xu؇��O�"	��a�ˤy�m �kʔ���ąc�{��%�Ʌ�%�a9q[�e�����L�}y'�وv]؅�֢�?�1E�}��EXQ��|�re㺛ݒ8gw׷h�2�K�)��iK�P�[/;
k}kN}��/�@<猶*yg��)b
([�K�3	��@�.`�I�T	Y� B
c��'@I��DMy�wHߕ~o(�<�'f}1�D�吅�"�ʳE]8a}<�� �E����}dQ���Ѳ�>�ԭ��@Z�0{���M�*u��o����(Fv��N��os���±�Au!'%�+�̚f$�n!�>e�쇨uɂQ�
��L)��i�O�f
X�ן'0A�QE����aP����� $�P��X=�֓G��@N�B� V (��f�s/���O��? ��;��~��}��	�f�8RnĐ�U��2?����b۔>� X '$:(m�l@�X8C������J�}�}�<�z@�~�{��*���6b����"�������E�D��,9� /i߸��;C���-�Gs�R>��=��ͻ��;Vb���*��*������N�*�����c��Db�*/�A_��`F[����+.2��n���U�kE)(��xƜ����q��S��'y����b�����>��ߙ�erG��������tZ��L^��v�.
0U�Gw�-��RRIw��1q�>`�!���Zo�J������i��y�5_E�g�E���UH�p#z�#`����~寁ו̌�[��v#�<����?����	����1�G6"�Nt$D_U���KH�`�Qr��6_��(����_�_�m�\*>b6�έ�^]�};2�1�x�ˑ��B�[M��	0{?DV�R7?��c�HP Pd�z�+�u��%jn߂�-�̘�P����a��YY����LK�迖�B6�Ad�X��}ج��e�$q�}4u�|�d[ ܻ����g�'cɱ�Em.��+^ɂ�C�	ʒ?�'��Hk�F�{���yٌ��?R�d��+Cl��-e�׬p�G����gr��ꦦ��}�v�?Ы��E���8�@,e�ʢ��dmb�J�����Ë�몒��O���~T#��` n`3��?�*�Gۨ�uK�cf�> a���^�j��^������'>[�P�!C�<��R�`�@Q������Tˁ�C�<_ɪS\6��!�H��$E��0�e��k��hӗ�j�N!���V�.�3���?�` ���I�ûf��0��.c��l�(c�o�b��tu/r��]CSmy�ы�]�V�ۮ86��9�r��dG��Nvq���B�w�ž�}�^���)~�h�f2�*����\3}p�78kt�'�Ψa>@�!]-��ej~zZ��h�<�𧴥$�{�f����1ok��]9E���0f(�~�赙��4N���5Z���u2��U�	z7���l��{#��`�⭎�fy醎��3��d�����u^y�]M&i9 ˆ����q�M�#�E��u�� *"mFg˚qL��R����}����DC��ަ欲o�8g��\�������K�94��Eiq+p��	�z`�����Ʊj酮�jFACn�\�:�� ̡�/#z�����k��-��F��)���¼/`s6уw7�TW3�E�eS��|��@�>~`���F�Q�����OH_j��=�h�^Ǽ���ny�3[�K�)�����&5���r/�JG9D���g��������`��x��ͭMQ��o�Q�b[�A�S�T�x4V�eh����2n %�v���i��:i̞�>^[Y���R��n+��8:�Ѱ�
��
���"^#f��N�qKG��5�xHņ����&���7�N�us����懲�<}��_������I	\rX�y���E���&}��p?�_).�h!��3�����d;�ԁl;�Ġ*���.�ڰ��s�ѫ����5sn$E����Z7��b��%�9��l&��9�[��&��0�pyuz�3� ��7��:g!���GJ��Lc5�===�.�����9����Ч���������-� \.�����ŵ` �..p���v˚_���]��ͦ_h�+�u�A�7��,Z�vM��n/H�I-��PX`ԅ�u�;�����'l{�F/V�Ӥv�ξ�'<�y�;'�����
W��Ex����ݷw%�i�B�A]o���gLR��PԾP��#�5_��!��͇_
���� wԂʜ���R¸+[�DK[�x�*�
�H��[B�z�����<aڊ;�=VD���t�S��i[�"!~�<�1i)��7��S��� n�4��.��۾�z��}��,N:?�u���ܗU�MFG��X�
T�Iw#gB�f��D�?����J.�}���ah(]^�N�2��|�J�d��x���Hf*$3E4�<R�A)�>D�M���������Υ+щ4�I�Ʊ0�0����m� �H��_�+ph��`-i����PM�)݁4�TI�K��݌$t���cFvDVf
j���?8�%qMk3Uwo�b�ޖU�8?J��w��D��P,�O����V��L*���	�Q��ͺ:�%-i��4]���k,�sޗT��?q��$�9�W���ȉ�/�b0���8|���|�sw�~�ǳa ���+L��'K�����AS�x�sr���肾͊��1;�B�Hg5]�*�S�����7���`i�C���{q��.)�c?��)���@Y�i�B{����|��'F6\�b}?� 3�~�Zn�b�*�1vR�4HXӺO"�8�o�C}&��vU��E�e�c`�H�G�-��(�~��L%�Y����Ppgo�v�4Z|S�q�1�
x�(Q���S'&����G�- ��ޑ�lxL�f���W�4�p�´�|X����X�Sp�2��>��P�@ӡ�8_�t�t2FB�R_�I�R�������'{YW�6#	�x��k>���˿����A ���-F|d+	r��q���T�@��7�
v�⢉�,��ؘ3���K�%�*��O6��mZ)L]q1���]L�6��� D�4�%�\���p�4��*J�ɺ�V��*�.q
".|#8d�ak�a����o%K��>��Juh�w.���^��"��#���d�(���$� J7���#�&O}�����i��S60�r ֧N_,�M�@�*��8}6^u��WJ]���o' (HB���l�b��u�_���<����߰P3*x����mk����'.K�|��wst)� �B�ĉ��7��윎@5�U�c���2r�	��,&�MI��=5��`wɖ�#s�-+�E=�-W���zi~�] �$���ۡY�5���QhB��Ih�����$N�i� �i2j�7��z��6q
�K��g�\ �Nq�=�z��>�z[��XQ
=��W��fἕ`��iƽ(6"Se%�$�5�ۥ���d�H�T�Q�-a{�\�NF�oV��d������#O�W�%E墴S���Mv�,bs{:%�J��x8�ifL�X8�#{1���&Ъ���
��ab�Xx)���N��o�!b��!�����8�%��w�KCgi���v�Yr�܀��=(�0\V�]E���5�c.V}sN����î/��c=�W2QM�T��l��8��Ԑ��<Gn�yb9�ܣ��uv64F��O��NKVQ�D��/a帎�)*U|�{B_y��[��l��l|��q)�]5�C��VW;jX�L�T*���n6/�o����!x,h�Z;uC��	Y����s��	?���N��9]b%��-w*y�f�{!�|]$�� �^[�I~M��{(A�L�D�����8��s���3����!��+����?hF����A�7+��W�Ð3���������:�5�4ө8YAI��t�c�'�G���_�o=�~��:NK>+d������d|#��m���#� |p��� 1�o�p�D�.O*�/���7��j▲�1z8ժ�CO2Fis#�I����BH��E-�G�ܖ�9B�c�W���L�W�� �y���jp`D=�L���˖bɦ�J���Hi�OI�aR"�X
A|������C��_ʢO�w�v�p1�ʨ�Q�}�8ތQU�j�߅u���$�vD�p�'ܣ���^�%|�h@L�_~��1da8!�#�AF�ؐ��0�s��Ѧ�o@���,�u�\��'�����+bov��(��_�&���W�m;^��fEL�ZA˵�ș]�����{��4目&��
ϣ�<o-��[?��/E������np1:���{rGPk��+X=��}���TąRPQty2��9��?(��`���^TR�|R�<�K�]�0� [Fb��[�pUc�3(m��:P�(��ʉKe�r	� U��n�7���e�X������Q
7i>Blb���Z�R���
���RnA#�o\;�&"�U[�59Yd�w1��H�Q��,�F@��S����ʟ���������G�|{���<58R8%�ǌi'q�t��s�O�Fr쾁���Z^"@�d(O��5�n|��jc�(�W�Go�l�g�����j�	�w�`1��A(��_\�+�r���?_un �Ȏ�z�������d8�I�Yn����[}�a�ZӍ]i(����)��8�J�}]���m�ɥm�M�3�����0�����|�FT38������VD]Y�����P�:��X�QeN�$oU�����F�	�&��tGI���}����~�^�0��bY��* �om�~y�ў��K��O����1���:ngj��X�6X��n��̑6���k��co�5|�~\G��:ozM4@K��ܶ,8�́�k#���U�R��1	�Z�x$&#�)�״ц�tA�80.��nkn(r��'�@t�ҭ���+E9�6��a�lҾC�^�M���yO"2�PQ����R�K]�4L�$�万�X�P�uf��Ytb�1�Tm�k�}����}Ũ���8��	me�(8p�%̨=Uz�EB-7�w�Gǰ@7��J�Q�pN�í9_p����fĶ��<��X�G��I�kj)iD�����r�~���2C�����X2��Y3��Kb��J�%�t0.l_{��xf�E�(���l����!�<��QN��/8�R*�;:�*\J@YH>�J�|*����R�@	oH9e]�ZP����m��7���(P=eH W&e����tff�!N���(N��BEBht�FcR#n�J��(���3*7����$(}�/3��M�x7�sM��~��rv��������}�yb�ӽ�SH���%�������]�-�]��av7�b���,q�д~њ��If&@h��b[8YȪ�q>��3l���@6�Ґ?$�1UC(�5G�y�d�RWݩ
�8�͛�[ޚ��:�o"C��X���MA�a�����ɵ�n��RDg�I׾g�0�l
0U�����g�g=�Ӹ_j˿��f1��v?�hRAJ6�鉠0��.ҲHTbJ��ihtb�Z�S��{%�眭���O�bK?O�>�;�Q���_�;4J\���0���<�D¼e	Ϳ�8A���&�s��������W�ƍ�
c^�{�a�VL>@.�~�y�ﰘ"�ђG#�?�{�� @jko2��
�Xh�`�4�����5�!Kw� ,�J9�Ж�H�#�g�����A��	���8Ĝ��挙�H�~�,�4F��5�R�/TL��b.���䨵=�t��K���O���,�T�8���6������VN�l�Y�u1/�`�#���)*�(<��$�9^:,�z��؆c�(�3�A��TyK��:^�Pw��ʁ���[������+�=�Q٩�"��rS'�n��>�AӦ�a�{�p��hФݓ��8f��@�\����\��vų��l X�L����.��������[��Z)�[�$�y}�&ko�,�f�Ϩ���P��?����9O�P�s/�|O:���\�dǺg���+ry���a�Ь����L��}h�Q�'�W���dIS`O4������C"�b�Z�k�^.V>+Ox��^���q�����U��Bi�>�Bԉ�K&�.�l.Q}��O��
�}?IV#�_@�>�:c��V�K��B&P��sF����ω�j���T5�Ͻ�B��0| �6��U��;SZ�r��,.�%��dZӘ�y�>����K���kr �y�?���=����[?]R��@�X��V�~i%�F�Hv ��#�J�
;m�.k��Z�	c���eI2��{�o?��x�1�p0s^HU�;~��!.6�Ga��&��M�}����������V��K�8|s;&�.�'|�̀ɟce��{��)�|BV�.�Q��Hь�Zp�ko��:L4�rlM��qEdbhw��)��4�P���7W�xU�
_�IY��
�=�ˠ�Z��vؑ�E��;.�
���<������_��u}���A�V5)_�l1v������p	M�gf>�jo��pW�mޞ5tl0�y�$ᇗ�*>�i����-$�^���W��F�`�V��x"P��EH��b���F���K|����0[���={��W%B�d��mwA�iq0%Rm_p팶�+� /��VB�e1����O$��!��H��2��"�	�|xKU�=G�%ȟH��B'��CQ͕#��`����S��kt�mz�V���[>Ln3�uFߕ�"E���p�f9��k1���<6J2f���+�1'��p��qWw0D:��m�Dd����O�<�NJ4��f�.��I��K�Y�q��P9AW|�w?uuQEj�Ml�G��&C?�V�k���<�a;��;��C���h"ǰ��C��J���	�����N�;��_��K��/&c�t��3�G�٤��Ā���_�.��:
����z���HA�?�Pe��}���0�I(�a�e�)��[W��*`������x�
����Z lm��+d)�%~�>gX#=���lC�&ݺ��r2�`����J�=��nf;�
�n]���Y�N��~���E"�I_}ap��o���v��4������Ա\-�����N�Ahv�2�%g�#7�����g��H'h���u����&��c9��f� �,����{:T:<@�w��eO�AD�J����-��ϧ��_��z6�Ɠ�/���c�gZ�}	��V�;݀�I/`D%z��a�#@��K�F���� D�蕂�@P���Mj��
{!���jΜ�Q�]��C��|����W'�B��|���TV��Q��B����[f��8�H��ӽ��{(��ur���}0�9�D������i���7r�?�5*��xW���Mbh4#�9r�ba���,#�-�WN�_���X̗i/�L;6Ž2�!)+�p�j���g��Vp�}�k�N�sNI|D�H��(_7h�TCi?��g�tEQ��x���x�M����g,]�H��� %;(�x��l�u�?�i��R�~��!O����k�(�F|�^�{'���s`5����}��[����/�L�X�cxTߦ�������a�m��j&�7��.�N�O���#�>\��?&�_TW>e�Ф�A5�2����iZ��2y6�!��U'�S���W� �&"�7���Ñ�޾d7���Ș�`K�㱐Ɓ:�?Śr�X���̜����dX����u�&���~�������x��
jS}���y�z��tp���?a~�l��0�1Vy���g�&؎R��U2�4	�ۘS�/F
��F��CNZ�Λ�w�'����WG�.`|�*�t�D�  ����>���9��SҷmI[̕s��7��m}$lC�����m��Ѯl��%��R�S���!8����JR�r�ܒ,is�֏��dR��,eRh�Y��|q*M�Q�SVHq�$��`��5pE�Nlގ����O�⌸TY���(9�7���	�Q�ynI:��hR�M��!�3o��m�c�Iy�����Bq���d� &�"��PHp�6T�C^������H��� �"g��+A̾�Nӑ�|���M��@��)�3����L�N���*�������1�]}��-�ۺ:�ww��F���U�������gt�p�	 +�o�`(��4`�Pc�S:�Q�cZ�"b�X�ﵪ}����Ōujk.r�5�2�׋5yzX�b<*u��W��.=�����<s�,���$�e�VF}�+L׻��2�g�CK@rW/i@9����D�]��*�|��D��c�4���]��?�H�<b��q��k��Q�Yǩ�giϬwt~j��ԩ/Ջ�-���?e� %�]�1� :�Ӆ��{����������e,��ݷw��°�E7�N�'?K�9�-SԨļ��Ͼ��8�1��%�`��\��v#��G�$_�m!%�6�s$E>�1�#�����t���z���&$Bm�X(FT8�1����mu��Ҫ䳜>�7o'Ed1�C��Ƈ��4�[X� \z�ِ�VrL�{)a�xS4w�7{��nr��?uo^��*�oF�.[+�
'�z��xU���3��:��D��91=�9D��DX>F��7+��}ׇFOх�^1�TK��\���f��"J�`i���j�ULE�p>�9��t'�O��*�Ѧ��툦� ���C4W�灳�j�w8X�fq1#A�&�{	�P��3�Y���Zk�zq�
K[Hq-��~�O���]���;��h�yT��ɾj�%�'�fU�S��jS��η�gF�'�=���맅R��)g��Z�Ep2q�Tw^2���ё���|kѫE5�]5_��E'�l�D�Fϳ�`[ >}4{y�)$ѥa�s�֧�}��!���(D���I���5�z&���#6����	-.Ǟ6 �����|$1OU5CfKg �v����o�;�����q��5k� :TRS���=P�-9�IU9�N+�%P��!��G�(;U��/OKJa��!��.�ً��3�F��G�}S+(���!腊��ȝ��Z�f^�=�Eӱ�c��sI�+��n��kg��u��y�L���P�ė��L�*j
��&/�8X��X�ϻ���k�A�Կ�Ї��N���V�(69ps�bj+n?$jC�˛u�~-�7;�w5��F,"��O���I��0K�qD(�?w]��X��ĥ��Ba}n[rY��#�ٖ~�G�d=S��՞��u�?�p��sP����܅*��B������ff*��.�2�V}���HPjj�Ҥv�(����ˈǆ�v50��!IFV����j?���8�}#+}�*>�" �$I�d&����V��^I޳�r�+�+ �Z�鱸��c����@m���3Ɖ�?��"���*
�N��FD���>�*)�V��D�͝9� @�eӐÅX2@�`�N�<��i����؀