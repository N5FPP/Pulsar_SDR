��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�uwC�5�b ��ϴ�	+�
Ct� "�J~���z����<
�����'k�z��ߵ,d�.��Z�Ӝ��2�x$ҟdL��h��ʔf��#
����;�;m�ȋ��[F��E� &'{=u�3jg�b�)��LA�u/5{<	����kk4�w���`+D+_�,Yw���Lg����x�*�����e+H�Qy�8�	���4^3�f�hOi3�Ø!��%���^dWp��[gN��U�v2�S���N�l0���V��IF&��c�eȫ��o��P�wH1���dm*n!��*�-�$���*"$G0�w奴���Q #$��w.1 n)��W���^���ϠF}wY�vT�A-7F%�j~���(�wu�8x7)��2&�'s��b_�zQ��3<duOW�w��kZRI'd�ᶩ�}���N�˱'<�I�hj19�]x
c�����~�k�G��[#���ʞ�M�q�N�y��ˤ+�ɭ���n�1�v��Y��Z��9�A�L":-S�+hj�y{ |8�sv�?9<�=�1U�'ݛ�i3��b�&�9G,A���wt�oy�����~ǈu�I���Q�y?h�4����}�#cؿ�侺���;�RE́R���y��mư���Y���2=��`7,n�1V�9�#$m����+1s0�ל�W�{�C�i�W��9y���y�O�w�N�1b����(Ò���y�p�#'-I�!��"9?ز�� e�B2���������0,[�?�Z�$\��t�\ׄ'"�	goR��dWp���M���2��M߇�eL��lF�;%o+���宂k��.�j?�2��ŖXD�>pwc�:�NPMҊ�Fӥt+4�_�v(DV�)v68�;/�����B�&.�/���m���+??���p��ߧ����(j=��7J����׌��e�Fp
� 5�Fݪ�r�t^��i����ӿ�[�;�DH�IG����4]��J�r����
�i[���c|�*"��ƴ/�B#�����!��9�A�T3�U�w���aݞ��P8�TL
K�nⲈ��?Ġ�ӕI�a=�.5�&i�r���R�33����<�W���Mh҆�m6����{��@�E���"�l��%�)��𱏊 �wA>"��3����.A���s�I$8�U�6HmAG/ +�2k���3��3�v����8Ed��2x�C�W��H���I�E��ʕ��.[�v�9��Qy�l����]�����i
��9Cؑ��t%������.�ţD�(+��%��V�

��=f��&�%����%�ޑb��#����
��*�qH�@@k6�ccPW&r���5NP�i�x��ZG�~�{�5�Y���$]����xz��Z�f���+��3]p���wH*��΢@��"g����Q�^��F�n=�Lў�o�sE[��V^�`g�u�%f�G�/�^�ŷlw	��O1�aǾ��T3�š9t�H�?�����q�'.����z���F�ϥ�h�cu��vŢ�)��U15���RO��|y�a���~�
���+��Y�~e�μWǊ�U-�`{e��Dm'��q72v�]V����.�B�+��Q�h���VK�$l����Fd��Ⱥ�J���':${��d_Dc8�\j���qy1��j2�O���:4��ƚy߄���F1���}�2+�u��o��������NQ���N�+
Q�͎�y��K��Ht|��������o|����n�Ԛ��23��S@��{��-s�cZ�H_��1��������ҰVW��\-����I���=�� �fk��u��J~��\��[�((艹��Pd���|�z_B7Y
�1v��E���8�F�' ��;ڛ���Zk|�h4�.��p�Z�ϟ(��S<��Y}P0L�+�'S�ى�p,t�_21��<���WoC�Y��+Y����LU�PV�sT�,,�+�_{T-�@H��5��Z
%a���`\�>fC1g�-!_��Ka��֭@��NE)�4����"R�	a��$½�U�K`�����9��imtT�G�6����Ҽ@�����g�H*A6m���Aw�M� [* *�?b���Q��8 #�UG�r�c����8"��W�	�ȑ��Ѻ���l�g���ǀ��5�Q��Ւ���iZQ�{�f�!�4���AĆ��&�C�tW�9@��a�t�o�����%V�%܇�H���!t�2 �I�e�݉=�+!6�˽Đαr�UA�;q�mM�AM�H����"�5��m��P����~&d������K�O��6\q���S����س���2]��14b1�&�):#�%�=�N���}�S&�/��Ȕ�V6A����¬m�<���7�[8|v��NpxL�F�Q��� 4ο�[^�H������$�e�b5�՞�o{;����F����Z�!L��2�nIxQ�CX�M:Y�����G�{�����J{�#��V{X��:���L���^)��a��N����u�:NcK,���w���Bߦ��a�{d��5h�b���Zf&0H�Ԋ�Vd�ni��8�LO���I��Ħ{���6�V��A����(����u&o��W�]��߰D�Q��O��·Aj�:���̜��(�l,�%�TyCk]�6��E�y����yl��֓'��ݝhjj"�Mc���?}ְ�|E*�f�\��_BYV�w�F�77|]n'�����OP#��ސ�bA��W��3��q_'��ݩ��k�F��@����ڈ1:��H�-���U�co�TDH���7��Y�<���2UⲨ��	?~<+�8�Z��D��%ŭ�:�V��|����ײsO[�+�'�h�3`�t�H"Vo��.wl;�N�>[ �,5���h^蟋t����ڰ�v	�l�6�^
;,x1*,��naHĬ�]����'��o�t�����l�=���r�U
�whr�k��F%)�N;􆿟��)�??���la����L����e��nd{"�"�+��8����������)p��
��F�hPX�x�F��uS����	B6�[Z��D�G�Ǹ��rЂ|*��F]�ё��6��0�"Ǥ�zO|�?W��?�x]*�?ǹ��(Z˖�����$���t�j�Plmi8N�!v��hӱ��8�ǯ�8f�C:b\vQ L6����t�����+6t�*R���M��K��>C�y/��+f�*s[o����ht��|����X�7X,O뙸��Mp֕:
H;�� �[��b��o��Ŕ��̰����[��*A��b�>��T9����P��8��S�����f�4<c,"2Jp�'�� [^tވ@ ���߶v� ^d���i��-�x��Z�0�!��s�LC� 9�Q$N`��@F����F%S�|�qG#�;�z3���D)yi�/]�.A{
B�\�1�bAw�; �	�!�ib ��řɃ�5|�#d���)���o� F��H���?Qb��{���/���1�j�IhA��/�urٱ���G��TH7w�(8����t���~c�S%
II�˪�K�yl�P����[�Q�Åj��5�a�)r��mGD8�iY�2{��A�^���R�r�㎥�aD�i���q4�Ʒ�t߰��қK�H:W<<���2#D%/�:�j�?C��3�u���\~��B�c��
6����{,5Ci�/��	Ľޥ���m �ɒ��4�f~��
���t�l�=�.�P��Oн�[����av�й4��\��Ef�i;
�˱����]��|w��]��8��EC�37�.z��I�!f���5�� �����?>QAA˷��l�,�LzF�V6Kd����N��"����o�۰��Ɔ�j�`�p�3SP�����w���r?�VՃ�b= �RF��@xV:7&�K�ɑo�G�ʻ
�C�pJ#���__�;�ע���wR�u8����׮6CK���AEV��Z����^/�p�߇ʆ��o�5#� �r��Σ�¡N����[��Њ`����A$�Î<Ǔ��',���!De�ݼ�߇�`S� c��)�4��.�n7��k2�4���X����>ܚ���&���6�F.�����U�fGǉd��j��a�*z��Q+!��5V�[��ɑ�@y;'��$��������Q�k���
=��^&�+������x]geE���0f+϶�F��p�X�� �,��NiPU��?��>j=��ܫ�엏����<E
��r�ų?� )�8S�nѸ\�T����Q��� dY�_�<������[����3�i�t$�$����ֹn�d��c��^ �gȟ b}:Z�Oe��]__��6(q�O���7�Ih����v�
��xE�hK<=oQ��U��k�(��I>��uC�f�;�oD�9;M=���f�D��ݼNy�8Bx��ք��\�� Da�Yϑ:� �>�o�f������
q���[�����y6`�R�}��������ޒDmP��Vufs5���!� ��o�h�B���?��nl�|F�DD�������&�rMa��_��f��%�s�)��UX��Ƅ�`oFd����C��q�yM/֊aA�}y�����0�W�̿�f��b@��5�D��������W�qY�x���������xn#��yz��b�
a�(�B���s�w%���g��j%S� �C����1q�86���b��;H�>�M�j���h�g;D�3�l���eN%��9!ww%��H������0�Z�f��q��*���F��߾q+����e�V�����UB�U7p{��-��Fq�$��juGۦ�`�v��lۗ�/����<�%2pg�P��ȵ9ٔU�D���D��[�KƲ�������i-?�/���JKB�/�=|\;V�����ysY#�2ym3�M��2P���Z"�q"��66�[�9�:��t�.4�R���Irr��y�>l���%������P��x����I;�UM��o�|�}V�}%�w�cK�P��7�`�]q���F���aw7�À��k�>i�	>��ٺ-�H�Y�7[?_���PEM#��p;��� �h�aj�4�[�O��W1��>OJY׹����������58P�n��~L���=@���V�Y�eU�ƃ�e�}S��a�����>2�rW�y�^�f��f���_yJ��Yl�oX"eIq;Ѕ3bzX�#a��[��� y�-MEK��5���^E	77�9$fK�H�*NJ�(�|���4Flz���QDq�NST܁¹u�"�T��r�2��Ή��o	;��O�}��*��B��1�e�Yٻz�w)���1��t�gaks�5to�����M�g����_b{wakYCg�qg'IG�ܫ1D'
��A��"�	���������<`]
�[IZ�A�D�$�>�7�K���RHь.v�1T>���TU+5��T�VԵ��>�̈́����Բ�d@	�qwU�#�=K��9�٧S�h�	�.�W	�c儭�p�I�;?�
�R���L�J��i�Wi�|�G��y����x[ ����CS��`p�pˉ8۪;�maf���]E�=!��@���;J+� #=L�4�>ͦ ]���:Z�?ȭ�:��7��9 M�5����G1W�
HW&�)��.�L~5�ήK~��~4����t$Y��g�.��<��&�����y3��'e�0����k(�_{l�y�5:,86>������9p@Ȗ�b��:�x�{k�a�r ���uz�bt��F�B�q������xq��=9�J�LZI����N�B`��,B�;hh��vu�9����2u�&,��'�ꖋB���WP.�d�Ѳ��^�aaO{�Ӏ%
L�S�v��J�~R� ��ٙ��I
(�R�Td��%鮬(g��1�/�M[���8�2��w'�[�$����(;���� ր�y�'�w����XԼKY
�_2fV�'����V��*~Qk�dJ��Vy~�|�ȃ>k�����v��1��	d������OJ��u���@Vhp�gޫ\�amI��2�W���"2Nnm\�k���M��W��D�d�0��uzvD��9禊��@�Z)d�4ɍ��c�N�����O,��m'�$��f��W��Z&��)�#�p*�l��n����D��f8���o�Z�AqbMy.�a�~�?�9������U�"������R�R�ǂ�fֻ�45�_�>�5Չ����,�&Fص�3�x%�D�b���2p�s���-����~Xۗ�0�U�">���(�N�s���7N���Ӆ�L�X�I'�1�R�F%b7�KO�����u�y_N���D�\��r��Y$���,�����]�~��ț���Ӭ��X�f<7Pr �竾f���E5�VA)���ȓ~cq�3?�pQ�<�����ފH@q��Φ�ꇝ]��̆���{��˹��n���%�u��LL"\��x�}m����"�mNAn���|���0������CX����[�,�����q>ҡ y�����{�x9WcV�z0��V��{@�4 �N�|�R�8��g���X��*8?�t���=>H��7Q!5.6�|���}Ɨ���ܭ�������[�Uy/�e���u�����fz����<	\�o�I�F�������+���8Ą�}Ĥ��.ո{3��"���|�OX��q���T��D�nmҺ�}�Eb.�8;�f�b��P= ���y�RrTٻAN6݌/{-0,��ђ��[FJ�a<x�2!r�m��4�l��H��=����,G�ʱ�)��������>���zZf�k��b/ߊ3�O�li�G��	_dU�x�W�yz�����f��;��9Q h���J�*����_|��f�A|~��0�6�2;x��F�<]g\d��G�_����������e�fd��S8�
��P7�pC@�d�~-��ski�Wn[����̐�-���&Z:�7RoD�4W*�X %��]��g��5�P�@x�
�xAc��������x�0����C�M�7Oď"�7�)_�'<��KI�_ $v�w]��}��]2Q�k�?6š�yH�wI1ݢ3+nSNs���&���C�॑V�D��
R@�Wq���߹���!Af���;:�K��6�r�999vb��ac�=e�������Vq�����=��3��k ���2D�KΚ��(vJ������S
�g�g��.�鈁
\��z��UeD�]�@�PJ�"0C���W��g�E��h<�T�;�֖K0����m�+T֥���L^��h�|Xz�\i�݌S��������}�����qG�/�zx1D^v�#ßbx\Ϊ��D�_�P:0k1�9w�]��F�<Y�c�X�jOůP�S�W"͛�2'����۹+Q�L� 1��(z��/4����O %�+?�L՗{��-3f� ��fΠ�h�2�I`ir�cnOu��Ԍ��H,"W��m8��Ϛ�������q71���rH�����O�x��t�+��h�c
m��\�#[��a��I�aXҺ{�r��W��3i����
J�!�SܓA�P�}Q�<��������v��I��E�8sG,��
;y��/��e֙���`�>��aI��Ʌ���q�W���pQ=q.����b�׸gV��~d9���%#e_���.m2d���H�_c�B�> ��w�ٟ@B�z��1M��ؓ�ׁ�Q�xr<m��I*�(S�Q!J2Ϟ�g)L�����WإG-�&�k���Y8�e��^3�ܯ&���%�0A��Php��R�=�/5[�������7.��Q��O��dލw����lrS���[i�Z:�צK��2,L�7�_C�D���3�hĳL7\/��

 ���&�bR�Nz�,��DB|2@o�Z�aQ�T���3�}���0����
U��yz���W�����#J�t�	�F.��*��K2C��Q�Ȝ�����dA͑!���負��Ή��r*,b,:q����j���x�+�ĵ=��U����yx�!�[���/`�1}���~�B�B����B��DXn,�,��u�"3t8`w��
-�{��кw�|k�JID��K�g$��}(���FB���fŌ5��u7S��z����b��T}x�s@� ������`��/��<�(d�S�2��V2�n	��9�^��e͓�>z �2��߾k���ث�7x�_���p�,�������S���v#��|��Htw�!���1 �z �gD\+����#|ag��U�F.Z��Dxw{�oI�4�[b�'~��䜈)��N3b�rRU�1Z|��	>8;sC>��)% nW|��9ޠ��Ǫ���zu2�--	�������@G�2_X����`�N�ZBg�g�mR��A �[M{��G. ���N@h��>N8r��2i�e#�^,k��b�c�df:�iG�:�c}ԗ@EbF�	z�҂?��h	v���.[�u,���]���	/����,�lj;�-��$<AVeCC���Q�{�
#��s�N�? F��s�i-J�-H$�W~؁�1��c�<�{�U�m^�!�vqi)����eȁ��qo�É�߳I�;��6?&����R�2����v��;�����=�$D��
���&t/�i~�:�It�*4�k.��_QѾ���+���K��3��WWk�o��*�i�>���N�?��3� r�"p�暫���oF~�!lT�F����ś/{o[8 X8+�ѹG��KŽ���_���~$]�>/�����0%֧���GYa�拱i�Y����\�����i�J5�;�a��ll|�yU2p�ъ�nt�Y+��rB9�Q��_��C�Sӛ�ݯ����S� Q�e�H�0�v�j�Kø��9P��gr�"o΄�n�B�~����`�m�ip!ռ��ć�ڿ(Z�N~�
��9N��fz�٘ �3p�u�6�	��_FX�G��!�i8�����V�2��}"|�T�t%���uQ���\!�%�C�^*���XY�\y���T�C�J�  {��_=����}u_J���G�M�t��;��x��'L,#�ORG�W��Vǫ��M�0�n��Z鋽ۂ�O�[6=QX)Y�,vq��Y_�aգ��An	�v��f����$��r���8�Rf�a���F?��v���F��C)f覂'�1q�\*��� I�G̺�����_��N//��#&�n�I��u��j�B��;2tl�+���V"�ⷀ�e �
�F���dB��,�2���ܗW�N�I�H[3S��,ċ(�u��T@�#��?� |i]~{0�#��.�y]�u�[��h^�F�:�
��@~J�/���M�u��:M�{dr4�@�Y���?�|������c���|���pD��V��W�R{ �1�Xӡ8^C�_Z���#������=)��F�sN�A�7�V�MqD��� `�P۱5����R峆��K����0_������������5�;?	�D-ޠ��8��}B1�{;�
 �w�W~:ge�!���o�K�};S�E�B�!�s�]��"�KOC28�t�w�\�� �C[mR�A�ƀ��HD�����C��!��4����0��4r�Է+q=!v�y�"���ᆮ �7J�9.�i�z���� i�|�`�ᬺvH  9�a__b���WN����@Q]+�����v���h1��@W�׎��8�� �(�7km��vy�f	,�ub���vp��� }����I�Q�����f+KD����B_Mw,�=��mn�1I�Z
?��8�\Y���'����}�WG��ߗ)�Z։�q�~�eKJo��w-�-�Z��j+j>���[?9H7�x<�z�ny�duV�?�)Gr����B�j������B���É��A�V����\�2�Ҭ((q���������n���;F�B-;6������q�!K�.XҷVn0B�G0�
� ƈ��J�_���eX�����% ��/�8�*�~j�j������Dr�ɀm��^ �%|�Fe`�
⺁�0t-�4���}Bظ��%����2��	dd�m�Wxҝ��_&}�N
����A���q{Q-��������������_�3Sq\�_>�-k�`X��^�P����F����V�V}%�B#�倵�_;Ms�)��̶Ӡo��l�9�dR�F�'I�,E�K;�>i��7�[k��yn�`b0�������B���WJ����L��7߹���\ԭ�k�"R]]|��|.�irC7�YGɢ0TKH�>݁��L�e5�3�_mp/'����8�ۊ@=�U��K�R�oZ�th��ڄ�n�
|٦޴��j¬�Ahak�,b�;��b�g���y�^�����s��R����/�p�{���<��x���M�J�۱�X\ Ϸ͇�T���x����ާ�a�{e7���26C�q�N�0�5����M��M>`�;P�e�)�Sx��H��]�ӳ��0aLaɜ�" �3/@�C1l_�T�ݻ��=%��h��S*�;E�L��!)(~��N%FwW<i@C�&�����q�H5�9tjc�X�` �b��?��w�|�w�}�pS4��q�!�`� �m��u�1��d<�E]d��G
~��G0F��ܿ�'_�S���,����If2�����d�k�p�#물��A�p
al��ajG�#����EM[�k��r��	�V3oQUSh�V�(s�:����|��@`�&M�W�{o�_��oGe����z�4�pieM�֏T"��&�8ϣr�4Ȁ(��oK-`��볩�'��]��Z�E@��{�@��;��	������P�a�u_w�G2F�D���3��a��xe���ԜYA�p�V��G5q`EߐS�t�On��YDL�.�+2��n�l��*e���N���H�	%/�G:H��7N4U���Z3g�V��������:��m�Pn�u���9��Q� @�����%��@j�^a�Y�˜t����N?�0����,澕7H�8DX�Bs��ꪽ���0D*/
��b��eE�a��.C��gFؗ@'$�4��$ɯ4Wo��}�iO�SF�mA�[��.}��9�
Axe;6!�Z׸q>ܓ~���
5!�b����¾��Ȍ 0�k}���d�ޘw��5��Y��} r��<�$�� ֖�!aF �u�]%��!�V6K2d��������i2l�zԁ�k�����.d�����&�NI�H"�(K�L�A�/���n�߿�����N�����]$�+�ݏ�����|,��� �8��$�c4�_p�p|��
9������|��=*&TB"���/�m��A�Mx��凉�)��Qy��/k3u"�0L�	Sjc�n�{b�����چ��Хf�=�,�&6��|���Bh;"�zR1�>g�]/��b��z�..n�C��ʉ�M0=e��󠐄�#(M"��owD��.m*/��o� ��;��{`�\x@���E���h`��'|�1P�I!�R*[�f##2�&Aq�G�B�ɻZ�{��$�jV�ђ��QW���b� %�&coz_��$o%U�Ur���<��"�[qL6_���ߓ�C�@�!�~�l�B`�qc��Kw�t���=�c��B��4�
 �WW�>S�r��9@{ǨAe2?1ͽG��3��ȭz�ϛ���<Iԟ9�>2*���@W��5�5�&���S��� ڒ=��8`�^jSOE���˂�,ɿ�$�.v��$�/3��q0���b�yN4`���7���&���ߨ�H䕟���+yN:y���f:��S�Y���O��I�K8�bJ8���@��u ���a�BJ��e8)�!K���-��|5�}��>�x����!�[�J���Z�G���]���ޟ�Bb���Z6T$�.�q�6@���������@�'�7C���UPiW籽@��P3ԯ
?����L�4���0��/C�x�x="&q0�����x��oܬ���⎄�:��2��*�qG�M,��4B��D�˾� �4-�kH�֚���K[�:��4�7Mb1{V����x5�Y�6�0&��$��";"G�o�Ox�Q��t�ǚw�ޏ�V����L3�]6�Xa�.3�#��v���Q<�J���"Z#�E�z	�Սêe��k�-��Ji�\����2����c��Q<B�5+J�@�Ot?�%���D�W?����3Z�U�J��y��s6��:����p�fF������vvF�A?8�)$�����m�q��%xn��Wm9�ޖ��r�����ă��lG���=�ƶVv����h�X<�!d�P����/���$�Io"�3o�?�H�>�H�<��y'�
��iC���0��SG��{�"a(a��a���s7Ӗܥ������ټ� M���.���s���H���u��+�ﰥJ�K��z��ތ؛GDb�LJ�X7��Ab�{r�|�2W�s�JS��*�-�6���%�J�~M�٨"j�k��{Ҡ�r)}�-�$U"0���Jo��r����@��P =Tg�,����H���.�U�T5a[}���r��y�{�^(v�P��f�W�#�����c�Rm}�� [S\´��N���7���g��q��@�ˆ������O�V� :��C$��)�,��u�4N{�p��!"� .v<�1'�%��G����Q���̆�:;��V�[W^�T�8ؙO��"\��M�'_�7��< ��/�j�cis	[������ ~�t`��_e����t`�Y׾�z�l�h���󬶻�$��.�)��	�>�dg~���F�z(���jSod��cʁ;2��͌�@
�2'��l�୏j��A0�(��Jj�k'��%c����rm���!k�@�.b�lfr�qrb������ ���BҖ�WW��Þ�����zTN�����U����	k��
�H݆ x�'v�	^�����hmߞ�p-���O�iA�>���XM�K {y1�)�aN���~���-�IX�R�0����[�+�Qz�j�_-Ɗ��J�#�#���}-�`@Z�"0^זH�ΥSB�����M�� dB��%�`�꾽[^��X.��b�A�x���H��!���q���k�5~skL���,<��t0�kS�$QL֐�lޓ�8���C�Y����zP��X���XƤ�'�F���L�t����id���n������*�K|�\DH7�$�O� �u������Us%�!b�(��wo�~�>Zd�Q�����D0`�S?����ɩBBD��QO�*Ц�U�B?�QVސH���\��HS��q+\���ЮH�.����o�~ r����>�;��^^����_{��� �W��6(�.C�jc��T�-���"�MLE�c��z��Rw�t�.���B��y��
����ɟ��:_� j��gN2���X��y�JbV���V�*��[��w��w�q�<���hRY����u�o���!QԻ"i��y�����nn3N}��|D�:���OEV@�t���{g��{C96��q�҂�aܲ��� q���	���Zx�k�{���^j/Ԋ�!�]����5H S�Xi#e?��!`T�
�|��[k���U�|�X������!�F���U�� ��.�z�*���k�!s�͍���s	���#N��oLc��J�Ǣ�;}["�I9zX $�l���OZ ���n��������EjƖ�;-�$6����n���s9>�DN{�Nu�R=�o�8��CA8ޝ�����$sm�	;��E��u�;�JwM,GQ�;q0*�m�(xƒ��JM���p��} ��
���gef�3\��� �H��F�@�MW��!��1�6O�5ңo�O�
�7���$����E�>X��J��{��
��F�y�O��.+)�b4`�����$X�v�go b���x�6�A�M�9�x�D�8<,��a��2�
��cI��wmJ��S
*CrWj�25�*����HG|f��4/�ԃ��Zd�0΁{?�	+�1����$����x���~�1�t��~�}́}��&��i�B%>�F�W��@�����6�U�o���ۃ�����<I�#yIS�a#���W1��z}M��������=h�
+�T��t2{�ѠG���@(P0����a�"h=V�5Sp��J9�@_�����ht����H��
 5s���ٺ/�������*t_`� {�*��������p�cGktu����D$뎣ؔ�8�ܨ��#OW�p��Q7g4�63���s�s�FT)G�4�R�e^8��Yf����Ի�&d
���s%�)	Ъt#uל�h�6U&���
��W}F`aN���,�!���*�t��.<�Sw���
-E�a��*0�Z�]8�0���q���t��E��Yk�G�8e� �@��p��XE҆�	JxI�[�r�ZfH� �><�0�{
@8�<W�	9�T	MM(v����BcmE������y�󡺧h��S��tk�M"lV�JS�M/E���ݶV�(֍7�S!������P�0#��d#sX8��!���:X����E�C�0�*�c��}́�Q��f�����0I+v�}�b��דH����e7oj��K�itʶ�Q��'G|"5�LN����+c��#��Jp�ϔ7�����(����U����Ϳ
L�h+#��3<�WX*������Ӊ[ �o�����r�D!��Z��>,W������b"4�S@�F|e\�K�dk�%X9Wt�!l��{�O����?/+���՟n��Ҙ�Et��R�ֳϛ�����r~ٗ����Ǹ�{����<ƪt�1�1|�b�z���Kuc���e����)[�z��0�N�%����b��˭�����I>������y�h�7=2��]xe���^�o��0�
�n콴契�����/�V'�9��o�QW��
C� }j����-�o��Y04|6����r�g��l9�}��޸�ʔ��kT���1�O��V�/�>�/B7~�7��3g���obL&z�gubө����ThSf�g�ֺ���ωD�J�*�v��v���� � y����I�M���{�\T��2���oD��q�����;Szb]��c�Z�d�+�ע���B0]������[}p8���d)kj�~�+�ʕ�e�)`yP����ba�~�%��\Z�vat
-qA���E�	�>Z�:H�M[�5#���R^r<WX���E9���iܴ_�lF�[����T���-�sR��h�	�>�	)� ��?E}L�;�^���`?���E/I�V(�3L��ϊ��8
���3c��K�w��̈v/�aw2��p�<��t��cˤ[;�`� ��~w�>�t��w�,&�SC^I';Z����v���v-���f�3Ý��`
�J�-�0����J���z���c�L��݀��o��G�b���Y�g�t�|ܰ7�t��/�ED���������i�Q��)j�￹D'��@H� ���&@�U�ef��x�VM0cҝJ�p��z�>����EQs�I�%�R���w��|��� �.�)��fx8(}X����JE$��N�b�h�b:c����(����8�[nkQ� ,C�UL�
5��N��^�7Nl[{�)=�!����5�!a�,�G��x�$���%"�5����o���x�Xm����oF�������s����N��2Fv�k�<B_Y�?�m�Os~��%0t�)fx�a�q�nٝ{/S$#��]#�� Lƭ����9�>�J,����}���O�h�:+f?�v8�=����Ϧ����^�:���l^o��Q�W%zy�Sф2Zwh}�/��/�xF�y��Ɂ�����t�/���E�"��jK���0��d�|�I�__�N@T��	h���&��CƝ����Ubؠ���$�=,$b��\tk��)��ѐh�ET�T���/2���(6�{cU|�F�z��y">TF�#�D�%=�-�]��>u1H�ݸ&�|�G��>���l	z���-�OF��y���B���VH���mӂ✧2�@� M��ҏ�<�KpL�!
��T�Bh������ubZ���ש�6�b�*�:K{�7��9���@x�!C��nU�Q�ȑw����o�r���Bq�p@ʶ�
�X�qN 	�P�_��c?	z���u���P�� J��{����'Tӣ��"�$;��P�����[��'�6���5�8����G��9H�}1�>E<�De�������"���ڐ/1聢�Sk%�uH��0=�&'��A�g�o8�*$J�S�f����HSP�wS���V�&!��ķ}y���9S�m��	�p�a�:�b�6�T2���Vn���d
�0�%��::�W��rZ��6���Z�@�����4l��Z�j2\��3S�u�k��d�����D͌�$�����פt�<���߀�.��������?;�p�� ʭZXӦ0R�F��QP��Yr��7�c��,�S����'E�W1�7���WkT��
��	3eG��?�+k�A�`]R�~V{0��������J���`���<�aw�Rp��2��ˁ0*dU��>��g�@3\���D/�O������]�e�0�G�1�FC���<R|��2�����������ahkƸ���먑����㮀u�6aZf�{:,�s�������[	Lo��K �rT��V��p��yɞ>۸d�|�n�p}�Ib�ޱ|�@2��̭��Ï�״a�D��lQ�h� ��1k�oؼ�K�ܕٷJ�#�O���.��.JC�ty�,��Mk���E���Hs����.��x/�,��4pS$��F$d�SV'�@m����N\Tf\憈�~u�y_���I��1�I1��B<l��3�j��;�W)|��D�6kY�cy`���
}�8%.���[g� s+>�i��d�?&�m�Ix2�|�W��n�%7��p�ˇ�2�1G�M��W&����a���Z��{�#���t%���˹��8�>@�ӻ�KҗmTROf��%d��'�(��w�%J�th�PV���1��0uX���@�괏��J"-�G
Xo����Im765�"�M)�Q}I1>*���LRwe&�!K�:��j�@�d�w6w[�ն:�6
U�*��@�c�O��U5����Ͷ�c4R�ݟ�#=�3��)�Z~E�g���a~_H0�A�a�}�d1��^�Hܧr(�S��~Ħ��&r�[n�=EIl����6��'=��{n���o��4 ��Q͈�愥����Ly+��
0b���D�H���'�}�tF9*%�}����X`�Wn��ќ������n�o�z7��F�&�@�|8�=y��=��v���:�T�2�?J_���w�U*�%�%rY%��,�$5h�0<�M��swJ�OİR�U�E�g�έ2�V���@�-7���-2�����ۢ\UN�&x�^�HZ�C���;Um���[�#�k�WH
P�?�S��X�D5�9����{񳉈�3��K�4�BUVVn\G�l�H��Fe??{䉵25�pI\����jLl��5,�2F ������ڿ�l�cT�Y^.�T_?_�P�������8KC":�=��<����X�?���ԡ����@衼5-{UgK
lpb���������1���\��aό�[S7lvu힤����/T�Oä8����p/���5�u�2���S|��uRȾg,�a�\�(d�����h<?�*K���?L�Yq}kQ�}w,kM}*B��s��pmv�	����� M~�Fr4��k�bJ��z�Z1���Ns��ʀ5I����[�ZI&���~Ƶ�"
�#�%5be)�&�P����"��3���)�O�����}�Q�F��[��Y�� ��	uIPՃ$�}�I�/nX��)��	�%����O.��F��"b�`W
_�gG�`���Z��eq;�)�楴Z����rC�����1�u��HܗQ�b����Ua�v��@^��4�-
��2dY��
i�\@U��Y��cS��I�N���bC�(^W$�~%~�<2���/��+$NP���\gX�WCR�[��<�<��dD7��tE2�m�;hoܿ���q)A�3�ܝ�$�#�O7H�i�+b��ܶ���{1�v`�ݶ�D���Jp�hI�A�K��i]��
��@�����F�8l깍�X3�&�@'?���C0��BH�� �h�j~-����(��{}�I)A�7���#(���x}~[��@��v-h~�;o�}T�����A F��H�=��
QW�������̙�hj�HK�=o�ܰ��V�0@ral��C���#��u�,w�i��_[l-ԑ�ڧ}�q���Ӯ�4��!��ڎT�Uկ��sϠ�\�@�n-)J��N��헃�p��)8{����!��������R�ï�Bn��Xs��^�n���`|b�--U	���IS�*�<�!)A �1ٛ�H��e�/��Z��eq7W��N���\�뚻WI���e�Z���KfK���)΀qO"�A�9�84u���5�i�2�ԇZN��p�o��(�~w[��j���2��|��~�@�����Z*�xF����\(�=-�:�!�Ր�����x�n�AS�<&���o�U��h�+ni���F�:�$��� �o�A�O�I!iWM�[�Nxؽ�[e�y�b��~���s�rT�Cg����d�_���Ö]>:s@w��u�9�r��?K�a��x�����be��vj���c��2�!�[.�m�7k�S���{����~�"�&��z�	Ѻ)�'�{Xk�R�A6g$�S����:R.˭�u#T[ދ���]�xfҽ$��}���r���e�܂S �rN������:$���`���!՜�l�5�t{����m�ٴ�AR ��L�=(d��>m���i:A�X�J2�Ӗ���,��M9LB��$r�u`b��J���BO}'�^mQ"c�A�L7n���E��n���A~;�b1�+��];_E�$�����^Wx�pI�9cs��!�Bv�/p+erst�������№�&���`��FڪU�Z��B���2³�rrQ���շ���~|Υأ��:���S@�)�TVӝ�k#$�:G�c ���̊��U�6�-~ӆ6cg�>2ӛ�����7�m�����]�&Ӫ�q�$}"�0I᚝��?f<-:Bh�� ���¾��$�A ��^�u��P��H���S���zL�����1��ѫ�m/��aq�-~wc�T�"C���xa�Mg#�-R<H��T�f��H!ųz���1�2b�b�e��ۓN7*����G.�7z��psO�ځAnԳӣйc��W���޹/$���8.n���V��֗�[G䉁7 �K�uó�	�)����kl��&���&�{ �v�_n�\��9���Xp�qi�yJYu��Ž5����!�|�kߔ�����R�#c��d�Z����^���b&�tߵȈ=v�u^~�h)vΕh���u�D��O��'�����^��͉E����K- <bn��R-#��d{Qy��ը�Q/\���?+�$L7 OI�΂|�\e����>��_M��j��Ȕ~����̜����K�����(�cR&N�����pu�ʿA���v��a���F y�B����&����#��s��/E|䪋��4^A)�Y6�����O��2���^��i,���gg���!/��5��/u�������'�Q�dݯԖJ��:��ջ8P+�5?Zw_:����L�E}�� (@�'S��/Ӻ��ɋ��D+� H�җ�I}s�`��Y_Q�$�G�M���)�(�;�.6va�����͈ҧ(�Fy/w)^��]?Y�]�����,NvjXi`x�d�˪�P�:,=�]�&i�ŘH�y��؝� =y	[2�V8�v�����ֹ�أ�4���<qL+�i,*�K����3\��1J�PmmW�qi��KR���ܡ4��R��g_�lb;Yzſ��\F��XZIxI�	a���qX��|N���ĸA8i��|h�}�n�-H��g��Y����[�sKf��,՜ٶ��0��5"親��6q|�䑀Л�c� ��2��g��Х	�]���4&����Ae6�͈�@i�:�0���;��H���B��"ziZ$��a:63[jo-n�r8x�'�I�}�t�e�u���=M����B:ɫ�z�{�����=�]��;��F�7�����TGX�n�;�����;z��4ˡ0cKX�VK&��A'�ܺ�(р����/PB�҃\9��>´�d#����;���t>�F���O��:��*,�*J)#�e0^��b)�]�)>��StCl0�^�����~I�X�s�]O�GK>8ee�ĭ>_�~m��Ti1�-/��[�W� 3����_�bF����_.��$� xK�s��Yx�N�Ϻ���0���e:�.�qj���sx�wEc��*�çϊ)lve�2'-���.�_-��K4�ԩ�˔��s��h�����|�_R*���M�j �
�ie:
�������h�Fz NGa���L{U���4"�k�eo�r�"�JS� Rhrť���`���F@d�Y�>7_C�����ɪ(*�Ä�M:§�����	�������[���8�'ze��~wkT
O�X��Ȧ�Ba��4QOu�R���e缓)W����r�QD���!Q�j�F?{�7�ybz��І�!�3�N�wg���Hs>䲼���/�l/��3A/����U������b~^s�D�.�&�
uo��k�x�x���s��nW�vWy��~j���P��SZ�l#� G�VMֵ����"�>jUW�/G���smXƾG�����}��q��_�I��iP��ƕ�ey�D&�?j��;���Ru��@6�>�~���Ɉ60���D���ދ�EU��N萆��'�a4*��C���ς�{��ڒ���Hh�[�m��0�L�寻��n�Md>*`��	;s��-�3"`���M����?�s�"����j��T��(p�%l,*TP����N7�cb�W�����m� �A��y4�]�G��P3Ҷ��6 ���/z���ûL4F��|����!�u����3[�`
`��H�7# D���/L�v����(bH�ޙ�0-*�3�t�����g%�ڀ����z�f��&��O�"�3B�4dҤ�0��Ue��y��SH��Ղ����	����\���f���ԏ���&�ˑY�ʹ���yΧ���!a]"S�������Ɯ�A�P����Z�*nrM<E��mm�:�'8�iN��d������9)��)�gCئ&A�k����61F'5@��H��C?���j�ܓ�د�x=HR3�n����՟�,=ɖ��[�����h�c0w��8�}	6m,by��V%�A��yށ�H�%3+ ҧ�0��p���&����n9m�����J��_3�@���/A�.��վ[�!�8��t@#�6x,� ��E�0�5�k����H�O��ɺ*:ZB���>���a�s�~�w�<������A����ƳLCB��*a�t��c�L������o���LU _s+� �uGt��ˉc�>M3�M~IS���;�F��a��0�d7h�6�Z�H�=��v�:"8Й����49(]������f5��Չx}w�1�қY�jf���*d5��-03#�Jz���C�*%�(K�i��������Km=$�{GF0Ux�@.�P��"�y�N�b@�;]B�Fm��{t�����ub��a9��y_):͂��0q��*�"����ϵ�,�\S=�yz�����1C�����Ԣ��Hۜ�&L�}�����]��6W���{p%���c6�u�:��*� �<�Y��>�����yv8(�A���*�H����϶�x�ַ�&���e�_��6-վ�*�����K�Z��5�Jj,H<AF�C���u�#�o��i�G���>���]��tk�� ��r�d��>����t�+�	f��e�_�[���&�	qs"TY��p�{�)�Rԓ�[�hd֝�@�/�<��XD�h�c/�	PMr3>5rR�z'{`;?)��={ �"^ү"����l��u�/߆�z��H�Ũ�b�5d���Mz^2��`�	ۓ��E6j�g��ڮT���T]qb�2�i�GSy֪@whX]�g1�8��9h� �4))x�SW'N�J��u;q��.�E_[��rm����˄SD�B�J����ڀ�vA��D��|f{�d�`E�F����B�������>6&���T�1��ء�����B�8����K�xd�9�Q!���f-��.�*o�%��P���[�'�;���2��=Vj؏�/�5K�_�Ϛ]2@�}7N>��2����	h�����Z�R��<��35Uq�c6��	�ħAu�t0�Ś/Xwҽ������L��?1J�����$c��O���K�ں�q���*�=́yR�}��u���]�uS��Ƈe	��3�a}2���=J ?\�@����[p+,y���ٝ�آ�rY�}�X�0�al��7�*�^�st���1]�������m}Y9/�B��B~�
�V�*�IԺ#��Y���~ �X�1WǙ�w�6f��
���{�(}}"��E����!���n�� ��-"W.��q��g��z�?���ǉ�H���Z7��!�FrU�C;�RR�Ҧ�m�W\&^��@���@\J��\E�W�1��mhcs�r��N�=�oz&��!~ ��mi��0%�6��1��xͳ��%�>(���>���nh��ŵYJ/)8�K�]�(d;���"���:iG3E� }庿J�K΋-�d<?W�W���9�A]��W���oٲ�"H�k-䑩Eӗ6q��R� ����ƻ}&������[��h�<P��&A�5=8(����4e���{��,,��l�,0�M� +舜���p�U�!{�W�ٿ�:�z���c��jR�P�������)f<-��Gq�ov��]�Ϸ�r�iSbQ�(V����f��0rE�ِ��_�rj��Y����y���U�6,��eA�*7���� ��|�?R��ӏ�Ԭ�r
3��<�g���S�f�ymW�3����������xнAةg;؜^X]'�ט�1Mۑ���>�p˸�=�� ��>��K���N�Q0�$+1}�jD
�Ɇ�K]̄��������ܓ�*F�)��	�Bg�Jp5�UՑZ��ƄKؙ�|�
 �Ƴ��(#�<�Y$�7��^K䉜RJ`MT�_*��� _��Y5p: _��7�_��>��'m8�P�E[�����s�8�˹�Y�^�,��ɶ�i��Gou���@������ ���AL���w�;�Hr��l�´P��~_Y��-sXf4"����b��Ӵ'�;��N��:vd��.Ѫ|j�q\������(��꯱;�/�=��j����]��Nn��[�;L{����e�-Gf�)�&X���������܅��U��f\{{�9H�I�����C�G��؜�hV���Rt�x�֕=�!y�����rs�8(���g`���z-0+��*(���>��#ͮ7[����tn�g�J��!�#�c�Ƃ}��<\J��mqM9����?cM႗����A��_t����	$�Q�WA'B�o`<{k��ֿ7f��]�/���노S����ښ�.�"��;s��3��fdZw9F��V$��
�ǘ&�ib5!!cb�}��/*m��XR9���䄢 V8x륒�rY�"@��	���]���wu�m� n�C�W���z,���,N^ڻ3X��ӄj�ף��l��ņ�S�e>��2~e���!��}�oi;-�h=[1��
K�E\�'6�.�[�]���Fb"����W������){q$� ��A��:oq�	�6l5"�P�ھ����	:���&Bw�Or�t���`1C�z�`��p�f%��Zj��ֈ��0�x/�~RZ�c(\<G��T�!ЛG��ԭ7�RO$����v~T���4uе����1�4����*4�qg�F��ؑ�Kn�\���Ս��������-}�N�7؏�w�-x2+��b��RY!��� QͅO�*�W�X7甄'�kh��1�m��Գ����� �2�-����00�����?5U4����?#��R���,��#�ֻ�Iސ��꡽��St@@�0[�C�ۑ!i��d?�sݦX����tÈf��t`kF���70a�qF�Mf�?��U�3K��eYL���#F�v5���IV躯�
C�u�}LY:����a�7%T�����:���v�U�+�$]C�6�r��h�c���S[ɿ|J�#�*j���W%��Z$Q�l ��t�˞���8��5h���>�P�=��ҕ�6������ ��x�=m�ۀ�U��ű�<('���f�w��9�I����X��� L̩�f�u8@uQ�ɦ��lƘ�¬�ƽ�m�'{���$�p��L\�@���8vq8���F�wաj����+j�l�a��?d|d-�띻| cw��������O�l&A#l�-%�
��L�bx�+IM۠��6�I����H;��ek';��wo�*3������#|�Q�d��G�`z�c2JR��W]�s
!y-(a�6/�^7��`��2�F�Ҝ� �bR�P�UfzN��V8<�F-��m}D�P���;�ͮ�ͻ�x����Ը�I�|]f*� ��kܮT�}�)!��x�̄
z�W�b��q���x�>��<F2�reF6��hn=��FԆ�5!�E��7�>;�bo3�<y�sg�{l'BZ����Ӊ�$���	J�d��|�|�������G�*�;�󍰴e�K{�����M�Unx�o�=�~	sw��ٲ�)riB�_7v��S��NYJ�������n�������u�Պ{Xu૕���k��=xX G���F��$!�Y=�u��^��'��\�u5>�)��ţ^��|���*�dZ�ؑn��֗z�z3�#P`0�'�%��%�Q�����C[^Ix�$�w��ؓZ�J>�� ^oO�i�;өVn�*m��etH?{�b	��}�:1��K�ҡ�L�� � �/��7P�&Ӯ�ǥT&��Q�٢x��D�Bc�"�,YJ�Z���3��(S��O�}8apr������G��J�_X�x�ʫ�!��"���AЗ�?[���h�̽�S������"����(�VL���g�n6Ÿ	@	�@��Phh�Y��	��k�:�=�4V�(p���"��*.-a�R�3�)�B�p�w`��������w�N�H���e%��@��:��+��A��чϴ;$7�Pw���mW��/K����r���UjI��m���p���uE6W_K�ʣZ�i���/T��Ǹ��׋ ��Է��\�y�T���Q��V������Se������@��/�vɨ�5��̩�=�y��囌K��GC��f��8��L������mX�C\�z֛�]1A��8�I���z�s^�#�������:�r��s���@��݁�����"�9�j,FD|�3�o}�ah&�Z�� �T�S��Ԋ�E�N۴`�N��)��X�X^�Y����0h��_֍Рˡ�2�Y_�*���#f�.�^5���W�WI�*��K�� GJ[��r��B��B!(����Ō�3B��®(S�k����~d�C�nQ��Gr����Z��=^V�⯎4�v�IKtc�I��M��t�G�܎�V�b�B5��ș�_ѵVEw�C�]{�d�6'm���3v�,��^|�<���	�m���!�%�E�#ġ8���5x����_'w�X;Q͗$	�)x�Bh�o<��]E��a�F�+��G��0Cbn��<!�{�)��k�Mm��$Y2bI���a�L;]�@����ൔ�K71N^P�#���p��&�I͛��8��L0QJ4��[�sIu��'0�F֓��Ln�/yyt%���8���:�]�o�WFpbl{o�cm�����{��ϕ&���nb��Yv6��",����5���Y��#x�JE���ڃ'3��hS�z�6������R∏��\��������)�4�.��D������N��[9�Paa]߾�
�3jI���p�韪�׍gΞ
��6���h{IJ{4��	R��#F�W/��j��B���GQ�5E��Z�R0�
���WG�7
�2ĩ����6�L$HfRǕ3��f��p�4�]#���qZ��O�p�}j���v6�C��^7�;�1:iN�ph��L���B��)��!J��%�:�(�)q��:�>�iSWa#�Or��Hy�+C�[��KD�ֵaKY��	w>u���x� -c=&4'�ȟ����,m���ą�>���\����*��we��pqgR,U�Z�B��4Aa�`��� kO �S�3R�cq|v��(OS�}�X�M|�,uG��v��+�6��ﰊ�5~P"Ů�N���)ǐ,�ȕn&�x�����&����H?��C�����P4hb�I�n��}��~�t�U�8�7���]sc�6JV��l���c�*W`S�B&ʬ�:>��N�*��X��33�fӓ~�6���zP�cU��kRT8jVJ�6�K�I�R��z�i��\�jP�>��4�!7,l8B�=<O�O�>�j	��\%�F�3���cs�
����y���s~���

���^yA������_R�F93yX��.��p�ٱP%� 84_�Ma6`ߘ�#0��?�9���1�E�Z%o*W�Fצ�=W����Vu����E�t�߂��Ʌ#�k�*O1/�t�њ�i�L���Sg��/�3*��lF�p:nY;ڋ~�GyL�Pu��?��4�� 7pKM`�m"7�zy.`@!J0wjC�i�~����X<�iߨb���0���R��Ҕo�6�L\[���T2hT��S��gQ.�Q�a(w�m�Ĩ��}/g���y�w$	@M�l������s��k��7�m����u+k��\��ղh��R0A��0�E��1�2Gvo������"��6����J%
E	:�|!\�2l�M{�O/��'<��jh=n�v3z0����@Á�!���N�����ߚ��B�L.<�E
��"���H��|�[�~�y���1NG������2\G �W��}���)3��U�u�gm�ǔ�I	�P�%�R��>\L+HL�O@7�����-��˛EO ���W2=��O���F���E�{���*{�W+�n<�36�1��z͆s��!{v�>�U���Υ�$�˷8yt��Q�C?X��hC�*ٻ�D� ���c�_u9$�s�����ꯈ�������)�<��HA3t��<���d�~����U�: ��Y��1��q(�Z�Y��������k��A�(.f����$(x�\�\~&�?�#TO��ґ�h�(n&�U-�#o=��E�닦g�座,������/^]SL%�Pvh��Z�	�s�:����M72�PC����:󳜗>}Xf��/�b�Ј��y�~�]m��"u7��Y��DƮ���}�Ò�0�F����Z�uP��:���O3��}ts1S
�u�����U (�vu��������b�٫�k��Qo�Rt���g�Tsb��y�u�{,���oFtV&3L.1�l ���d�j4�fxy��X+���r&�P���8Xq���(R�Q�pUz�_<�I�v��-(�x����ͫ��Y"^9D2�~^�a���b��K������A�|�ة1�c�w2�A���Q��l[����(�����$f�r���0z�����F�Mmq)��0����D�Lؾ�X��W�^/���y��b<n'�l��uST�?�ٙ#Ր����
`���q�r��;W��0��j
�,�L՞h?��Ug���L�w���0�֛�~�a��A��jVa�����{+�Iő0h� �k�W��e��'��G���L�}]��=�i8��l�ު7��a�w%������F�p�����E��{i҉NnObʊ?�e^��?ӡ-���}8P%�X=)�!B��J�A�>�F3�<ڢ�ńU ҉�Gk����9��,��tL��>�Ȧe�~��]?>�} ��D��F�[I���,�Ä�ɬ�IĤ���!(�
��7~c��Z.m���������<��jA[|��i�J�C���o�G����ikD�CՎC8��W=y��o���Z`lo�CVH�Ԁ��1d�F�%�zPpR�j�߷���G�k�˛~��t��H\q����f�Jo��\�#Ѝc{D����i�[Rx��E�8�e��Y`+n�^ǔ�����l%+��d�70υX��ޗ�u���Z�HeW��4T^���{�\�A���!��٧����e-�=�@��#G*�6��¤W�<��ti4�󝩀ђ��ru���k��y6�k5�#$�O�ސ������~\>�_�q`���	���:��m����]
p�(]���f<���0�̗�Oj�Jb��� ������8�fJ>.�T-�Wh.|�@zQ�����=V����.�E��1����u1w���Z�X�+��#5�=R��8صcA��s	Y� ��*.��	4`�DΩ�sjZ�(�ڌ���:�0����HԂ�L�u?�Y!���Go���ņ�&�KnIi����o�R��N��F�q�p��L38e�HV:k���k�]�<n8�x�Kdf��1/��r��@�} �h&�-:�}	�'��<g̀�?���p��U�S�v��o�H`ɱ�$vX��t���7z%�5(�Ғ��1@�Ħ�}}�����@s���Æ������B������|�y�OiÒ2�Q��Djl�_>�y��\-�Sr�8\��j]�Ulڻƪ�g�]�32��E�%�A��N!��Na��:}��ڐ׉�����P�6���΃)�'�5�f����6ϛ?�_4���wЛ�����Z��+�V���6�)�7C^d4��9�OL$��5R%����l99�y R�3��@`C��Pk�8ƻ�|5#C.D�;5w(�n���|����6�"��ي��wZ�j�Ɠ�(Aٖ�"o�sο^���naZ^
ռ�@w�"ɑ�eM��fB��2W�[D;b4��2�+���wu���Ɋ���"��������.~��}�S5:�:��(�Gp�l[��>r�Ґ�D�D|�
�d���z�LY$��I�>�;�*�(�.��Y����G����&�$�;}�՘՞���J�|�?x�S2�hqy㼥9^�IC	���U0�}��zC��Y�Tp�!	|01h�.|�]4�Ws�^z 8��=u�v<�`�;̘y���1���k4���U���W]�n����՘1+�~���3M���}�Fm�Nj�;d�W��8��"4X�L��'��dl]���<0ַ�����#(0��{c'�B
t؞�!�i֫|:�h���q\��(�uLB�t<�R��G<�A�-|���Q��%c�_q�M8Y!]f=����^����=ŭn�X�+�'	��eU>�eB�	q�V�#\D�2rX4۩ֶ58����8!o��-ׂ8շމ=�q�E­�_ssߗ���v%y�~��%N@~��~��r���4[}�׸㮓xt.�cN�����;iqGY����i�&xg|��2c���D�L��'V>~~�73~�p��r;�����/ƾ]xei�$Q����ҁ��N�嵾���!O�=�5�'��&UzlS���Wo'�S��<�Hr��*)���7�9�+���x?(�{�:�"R7Gyͬ�&�(|S_˻��%��Eڞ'J��+4*uH�5�Ȃy#�끢_h����w�[	�+ �m���ĩH~f�B\���\r�����:�*���R�����Zt�㪒����Q��0���|gf|Yvv���zܢ�W��Q2��B��	i�)a��زnl0��xv�po�4��R ��E��	(h��N�~�ؿ�2B{D�����e��&X�
��J��x��uh7�]6z�u��<~q�Br�u��V.oh�R]��_�wJl�,4���V!����ﻵ��]�wp<3yW��(
�h�D���u�۾�ē�J�~�l�����NIGJ�t��O^���:J�}�A��8���T�]���b��^������c����~Oa������0��nf���s;�b�
A�Л*t� �@eX��p�l���`.z��6��)��5��*Y^^�ע�TΩB�A>C�b�-�x�mh{(/a�H@>��<�:�'�Xk����(>դQșo�p�������6�n�:kf������T��`��5rCk�����?]d�#1���ь�8O'�FZ�37�o����F�1I�.��&R��el�n7�1���9M�6K�����7[k�I�%�Ƽ�J�k�P5��0j~��Pq�Ц�	[��Q�ʘ�)�&��](�Ԥ���S��quXC�ֆIS�B���E���wJ�[�J� =,QPZb��U5q���:o�c��h`���Ow��Z��ۦWǲ^�8x�c�֓3�wmxvz�}7���������\\@�,��nF��m�o7�_�̡($[���c��D��'J��UY���J������,1��ei;�%��$������֞�vI�T)p4�xm�,ֳ=�����3�Ƣ&��� 6��O�H�4��b����m�����b>����-�aH+�Xt�=�HS�av��#5m���A$LX����JD)����W>l�A��%^ $�����r�-$Mb:��z�c�Y,G�����)�ӌ�$�"��*JM��*҈B���!4nm��@�Z=im�X7�ס��l��N0�絰$	X��-�=pR佹��c��:�?�7S�H9YbC����������8a����f�d�w��rГ��M<��tA�=���b!��֯
=�[��&S�L�)ڣ�y���k�˧[��8cj�0��:#�;9L��a� ���k�P��ͅ�8��'C��拃ʁ��,nMk�}�r�)�?io��ߗ��l�|�'�~��r�z�$�F��?p_�!���)$�@g��a��>f���%�A���(�8��߸�<~�=�\��CV9�2��O�W�Cqn�/�j��v�%@�b�vnb�jv�"K��"#j
i�<m�L�Dlˊx2���h��\9X��4-�<�8���������ߡ���&,�_��tĜGOݠ�&���_kj���0�r���u�ߝ��t�ҕ=�Ua���X�Q��K�^�v�(���4$%SG���[�`�h��\c��
@} ���m��T-VlB%�$�|BF��Fh-~�[�K"?��s��ŧx����2�41TӼ���1��@��n�"�s�o��/�O(<���#�w�����I��S�jڹP=0��@�̅x���z?��|̴��}s<���8�I�hYd�K\��dy6ٕ���Ѷ�@���0���WI�}-�&V�V`�W{X +�GH���P���o���s�>��>X���+��h�������ژI~WH{/�#��=�V��7�в�Vg��odU(,����L�>3�Q~"y/M ���H� a�����K)��K�42��t���[ڔ1�6��L�v�Ca���G���g*��G7�"Ml�<��i����X�����7����aO"`�HX�!�/�ᾌ�
H݈��/vqya\�aVj��\Ԋb����ZÐpP�5��1���-7�@���g	�V�D�S@��� "��-!��H �ܥ6�^�jl�=;�#�m|~��
M>�,���$��΍o��ĸ�N�Q�c�(	��WV�*պ����T���2�`|mE/W��J�;
���S��2���y���}���}R	jqR��&�.=�e�+!x�_��6�F��Ex?M�:ML���`5��S ��y\YԮ(���j���i��َ�S��9��-9��u���7��5�e��6Y�G^�]Pm�gA0^<�k(��`��h�?"�� ��r��?&Ŕ�)���k8W'����=LQ�D���~ ���z�_[Ά�dV�'�d�(/�5	�6۷�R�NG:�0B*4�K����~	�������&�Zʈ�ɺ5��D���'�|�x�.������޻r��A?���apE+g;4eЏ4�mհ����H�)�,}.�9FK^�k%��LRYEc�ˑ
vD�y��NJ,�6�d=�"�2",N�g"�P\̚4˧�����I����������"0HW�1�(��ב����{�C��#��PXn��|Mn3	��hg�urs3��L}��(���J'v�)} lJ,��?}�J4���2S�>Y�\��d�Cʚ�-Ux�����3�����wD��q���s�0j���j)�
���:8��Ɗlc3\:D��<�j���(�x�5//�����vi㮐f]���ѤF?Vw(��l	�:��=�q�"#�A1�9LNT>�8�ΔE�l�.��t�n���Z�e�4fs��徆�v�S�Q�)4��~Ս��j�^�͑�a�����n'"�-~�j�_ia�\��
�iD���}k"bC[�Z��72�Z�a�t�<�e�ۘȈ�"������I�e���S���j�~��߲��e�xM�0'����E���RKYy���LM,��խ���t����3��	�<6{a���#�%c�ô\q��0e�!'�X<��vo~����ҵ��Ͳ�t�����$55&u��W�5[̶��SL�4���Aɼ��qBp�{ �)oh�U":�i�~���$8Y�d��^G�>��:����Rk�N �1
��+ 㱬1�3���vL�\X��x�H�2�@8L�5Y�RcR��+p��c-�|�O#DZ'$%�Ř�zHn�>wO����B���.:��<!6��o)/��i-�7��s߯u�ʦZ��p�!���45"7�<]�^b)����*&b{k�d%8 ���B|���l!�].�Ċ��.LlA��,!�l0������'��ft1�$������}�R�8�r�͡m?�ZӜ9O����qmfߛ|����͡��P]�<2k�k�qk�F�3�v���"
aӵt�ě��8w6���Gئ�L�+GV��1mS�oklm���e���m�z4�T2�yu�"�'Ʃ���J�=����ن������n�@��|b~I������k�Mr�O�)��lpOE�␢<�@�sve���W9%�	�*7��1*�{:r�`��MG�.j��ϛ�R�/ew���ld�$�Pw�7S�|��A,���q�ш	����4oɟZ�!LQ�>����\F���Icߕ7]t�o��i��T�{��AUA������\�b{_2�*N�:UԬgk��#���7_M���U���3�[ �D{�_�P��v�|LΝ���Kb���e����5b%m�$�I�1S��P~	�D��V�r���2�X5T�Z�G��<�\�dB-
�֛X�K��#�5@���H҉�%ٹŐ�G4.WgJ�MZ�_~ǵ����mbF�i����ѻ&
��0���$����4<W����Ʀ��;��Gdzb���R��I����
�?�9���r�or��lv�(�nQ7�xDG2�ܟ܈v^���ۘK=��Y������NK���A�rO�J>��}�F�9��N2l-I���Y%C����b����3p#��#:�C��ty�`��tt�;�������gv���o����J�; Q��c��"n�,�2���@͎&��j҆}�Q�S��Eg ��C5~8���-N m�r�*�D|֘bxO)��Ȃ�ɗ�&��Jpm[�q�)i87K$���s���vn�����KZG∁U�jj̎�	�ӱ\�-�Ͼ������5s���OsK��i\x�_�6v�"��B9[�L��V�����-�^�uJ�Ѩ��-GSo��E*��1���`P���5S�ɝu/�H��1�(EZ!VQ*��ꄛ�ݨ��y.^7�������'UY[�0���'E��^� y.�j��\�
�����a�K�T"�������q.�Z�]{o��l�I)��T'�p�i_l6m1�㚽wC�ܛC#�nY2m�0���-H��Ѷ�`^��[e-���m��.E��ڇ���}�z&G��Y�$9���ށ����$OB�W��n~ec�ܤ�~�]%~x���,�4����c�<������}"�b>ˬ��ł�U�z�m��BA�p��ز�.�j�?$Errv��GC�����}V�h��W���`D �d��f�bG ���gn:`����4d`����-L����H%8d�>�\we`��p	��43�*}࿙I�J����2���)�Z��U�^kvuuBB�w�8��z���fJ%Q#�mn�݁�0�U�y_��u:����w�ʋ�&n.�:�9�ϥu�@�[�q���%.mCU���ȕ�>���
~�;~H�m�mK5\2�~�cԴ����ޖa��u�-�{����*�=;tǪ���J��-���s�B4�WA����w��C:�=���}m���D�tW��?���b��oz�q��8��Ch`�\��JXF���x�.Dʪ�氆cՑg�ѩ���x�ms3���u��څ��U��I���\e��k�����Z�����~�Rm
�:j���?�L 5��u����B!�v��X�~
���0"�Ĝ�c���9C�V�P�èq���ހ-�=����R��B�*��X�v����:eF�#8	_�>q�������I�Ȟ�~�(ƪ��eMe<<+�CTc��i�#��?��'j�E�+S��8�Q%��q%j�K�зx�W{Z	�T��[D�wm���cO�Y�$/4�W���8������6����~���H���nRG���^�b�����2����f�{ӿ}J��]�(�u�&���cUv��0��wOS��HH�G��%et�p&��J�t �'�q��}�׮#��`�*�t�znkg}u'\��M���}f#��	�S^���SU����5��Qs�]?��I& �r�qhe����~A���i�~C�g)�^DS�6Ϯ�N�	0�g�tO!J��M�'���u8>���R���[t(���`�o4��{�l���me\?@[�j���ҵ� �àLp^����|��$IH��ܶ)��{y�ģ�ڍĥ;�|��,ſ�b+�r.̰��
y������u�"�	O�������ۦR���-=�������y��8�'�X׃%�����MZN�\��r�!����Y�GL��t5��0�?�_9�4�.�^��~딬7.ʒ=����J[��M>^�����y����7����0�u�4E�=���R����RU�}�99A�F�a?m~���D�(���1\,���ovJ��Ȩs[!V���hKrR2��J:9�p��?�q���`ʃ�Y2Ȳ��\t�	-`�<� c��Dy�#j2�>3�=���uV8����p�C�� ���Z/�A��km�g{MC��Rј��Ʉ� wd�? ۬�Ieu�~��p.�,	@���S�s�X���M���]�8����?z���
PǌV� ,a������`������I��[a���o���#������]�x���5�$�S�����3����3ԬM�n�1�wm|i��u���#;w���鰻<5��$%k�z!5���K���v�q�������%���V�d�rh����>ТS�(z�D�zr�+ęU)Ċ+�iro���T7D=�$>��%a�g�mEE�"d�F�q��>��[u�O��NlUEb擈��Q�Ͻ��l�I���Af�V/P��W��+Rէ}�,>�=� x��t=��O^�IND�?(gI���g?���T"��lP�+P|'c�o�L�XY1�= 7ױ��\n�o�Fq��Y���4���j�^��;�Lˌ��6:0�d�9�:T����j��H�Em.9���	��PV]�|��Y��_� qt��d�����Oz߉�=�դ��^úWz��,�+Qb������sw�؉��Gx�΁>(��g�İx�����O��� u���P��PFCes4
F�ґ��xVO�Ai�&&^���7��Z�8��x9�<��91�u��/.߽�\�@S�hy�gA8�o������!�ٺ~�
��U�>P�PV"L{��!]��zd��x���q|m=kʅ�:p3���˝���{�b���͞n���7樚��If��e���P���e�Hw�`pJj_X�`1N
3��?9�����zϔ�F��N��������n��&���'�nP�/QFav�ϓ���Gɛ��7��)��B�˭�ѭ���7\��?��v+�H#�L���=�U�=+���]e�?,�:��Y�`�n]�!�s��+t-P9�%]>��Ν)�]	��_$�����hq��C�k%�a]:T.V��v-�;1gDNX��Rd%�:��p���1�F�	�q���lt����}�DƷ�$��61B�Am�P��D�Z�q��Ƈ!����%��W�2�`?�D�������3~�/�C��ܞ���v�ӎ�w�~�<��5��nK���,���E�Pfl ��m9���ߝ�$�l�V@"5_�Kp��S�]v$���/Z����Oӗ�Nm�z-_P�87��o��G����
�w�����C�5��s ���&4�RN��q��0X���_ ���2���w�}��R��hk2��O�^���jA �r/y��_�47I��(��Sf�g6כ�i+���g���D�ulp&�^T���/P���iu�4zu��p5����T&>eg�A.e��]f�
�>vm�t|T*�U��u�aw�*�IwQ��%ĬH�|�<RLp-���kL�<�T�آ��U��g�E�c����H���j��:���H�l,7h��6V��jT~���M�0������=T����>*�c��[���~a�V纜(6� ����Z@�.��:Y6/���CG	6�s��WOO���^!w��Xb��#^9��B&���q2)�y&d^��Gx���x)Q&��G�뀽~QY�t���]���m�q��FF �(d+ed�s_�U#�e� ��W�.g|ʫ��f�����)����Xɰt�~�y,}�*�̇˕����b��B�Y߶�ɟ��P�Yj�fZGpj�Y����e��̥������s٦�ݥ7��	�p��	�M���(��Y=�L�{a;�	3�-]M]�b��*4zu�d�l_�Z(O�c����k�6�[7+�3���!
3�x�n�j(&�u��|�)����/�Z�zeUk�&��n/w�g5�^lT�2��r:fU��ً��F>�x!e#T����9>TQ�G$��k�<�-0�!9i���z�λ"��0HGK�o�N&�����E�).5�R<������|lu-�b�	��wmeJ(��%Pb&�������쾱���������`�rv����y��v%^�Pѥ������Z�=d^�
��9"*�-y�r`�C8��Pq�'=|�e�Д$e�gS�^P�\��h�{��Y�=iZ	�h�,(#7i�f���M��*m���H2[��%�HwP *	ǻ�޼4R���C8�J�RR�1�+to�Ӥ�6j`������|RE�tR!������-e��P����y�c$j`���X�6�Et�cN���lc����`z�{?1�����[C�Ǔ���"T���^m[�p�z�f�Ѓ����Rs�Μ.nuv�ǶK�~�`k͓g{