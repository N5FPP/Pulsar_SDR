��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>hs�*�U��Q�����0<���ij5�f=���n��Ŭ�po����-��+J�j��7�0γ#~PF�Ç�n�~\ݥ�����I�'��nn��a���+iB�o�mp��O�C�HnO��H�bМ5<���\J;��r���:h�"0�z���7�=���Hs0���@B�[�|4^�y�(�< �,&OF1�G��b�y����&#O�՛��.������Ok��ePR��C��`ľ=K�18t���IE�����y{��`tp]���SQlc�{��r��Z���+2Z�R1�'�e�e��H��@S����|l��,��<Uz�ǵ �״��@*�'��r�=�f�#�B*���*^�IO�u4P��l3w���JP0Y��Xo��ez���"���9��`�S�,��]$��ͪ��ot�U,��;lO�\�v���|W(g�3�A�__Q���dT9�N���+������MVū� ����`�)z���G�P]�/8��x���u����.�$�#�^����g*��k��S�aǹ�mTBJ���Z�Ӧ�x���r� ��^٢����#�Ew]���}�Ο�=؛o���&KAT��J���	'��?�E�}Z��>)���@T��?.f}�@m����.s�k�rn�oOg�AkP�2mH#j7W�j��g�6�
DL���દ�]#�'xy�Ѧ3����������
0A5��%��o-�aspy�w�ٙN��"o�9��r=?�c��$�\֛�	�5lsf�reُ�}��}N��w�]Ea]���2T����d1��`%#6���� �^v{ϒ�綠Z:�K+��o��(̲���hg����X���!2��H ��\��Rc��c�u5�{ >B|��X�ˆȋ밙��T�4�/���3�h��0�{=L��$!�s�σ�2�l�T��Щ����-��W�3�HA���cZu�-�&1�_֖B >��|��Mц�}��6��s�&|�g�C_=�A�+1��3=����Ҡ^�:}y�oO�=��'hf�UA�%&�sf��������$��K�;�խ!p��箏��c�H��_ϰ��˿2��MZh���-��hX`b"ޥ�#�����5��A��q���	�H�|{��MK��
7x8�[tџ\��!�%%J��z"��e��\�1��d��k~j������nDc��@Sr{ŀBg37y�v���J�$����NG2*�&l�=؁5]���v�䎬���(�!g���i�x�����&t�[ҟ� �J�T��T�p�e�֎����L�p����-ìOB�C 2�
�B�cZj�H0�t+�@G��+׀pVfc�2��g�\z�;�����OQu���y��ڮ�X@w��!-�ox��
e�oY�Uv2~pI���b/|���Kz�Ś�b��`Nņ^iML�V'�w�<�@��)p@�-"�N�������D�Wg��;���}gK�Y�$�}A��pr�F�>��xV��Ыs�Tn��'͕_+a�Lv&F�c"�EvTг��d��M>��&���1�R��n��.��׮.O��ͩ%�2���vמ١��E����q	��ǷT�������É�{���l��;\�Iأ�O��I��^t4d�~�8'��ʥ|:��{$�u���k�(�`�;�!aJ��N���[�V�8=�h�U���@�:N��{��cd*2�:�Uk�FIfw[Pń�r2W8(h1eZ�k����)���Aè��!	��5r;ƟT6��_=�p(���Ѯ8��t%	�W��_}u�:��|�@f[/RjT0���Ъإ_��U�)_&�3ycO���/Xg̘�j��do��_��@cs۹��rM�@]�qU�H�;�Kd��V�{�M�)�N�nw�66Ł�J����+��q��/Mf�NR�-�7e�Y%��%=�=h3��~���Lh[Y�J��	�G�ӬJ�,��-�t�N����8,��9�VԀ�X��pUý���<٠�)8{L��}D��u��86;�k�v�L�x�N��ߠZ7o������= *����`��\��8�gD�T	��)<nq�ڄ:<�%L3ꉎ��x��VS6��X�{�������̡���4�L�6��|+�	��y&����9b����Tp=�b�+�i/G�>��'��0M	�	U��n�mD���ŉ��R'l���� ��u�m��ּ����ʚ�C.�����O������G���6l[pf�t��wL��E�S�����w�)`nN4���3gM������M��.@,��;H����.�hy�����	����
���`�m��&׳��T֌�,�� '~Em�?M>��"�Ҁ�P	�_ ��.�0�,O�1��x� �����n=GR�y��Ҕԡ�Fȑ8/e3��ۇ�%�)H�}V,�n�\���*�Ӵ����~��i3yԻ
ʨ4z���C_[��dh>'���G�5�/���ĖIV�σ�G�(>>�3�$�&���W۩����b(� ��#�Nh��J]]��U���hvm"�h��J��a�e�p�2;B�8�c���c]7��c���.��cO�~�{�t,Nw�[�ARb�δ��qm!M��Ă�a���i!��}.xQ%s����ի�׌���xŌ�I��+�=�u}y����.���חv��uK��$KN�n��)-ʛ�i�v�~3��c^{_��Z��l���r�U#�NB�h��K&����Eok�Z�
�'=��HZ�<�)`���p��yD�K��2}��ߌu�2(>��k��q��h�b�xO�_�ɝc���j<��v�~��:#N@u7��N�\ �����v��7(�3�M�9�#:��i� K6��YX5��q�l��9R&��{�\� ����op�F��v�KL-�2������r69���v�3].s͓��5�p���)���+[���m0d�8�(u
xm�K��E���@�:N�q}�۷tc�7"�����"g��k���˂_u���q[�x���78��������'@Q��f�zJu��(�:�Zw�Y�`��Q�o(1$�3�{�M%�䤿�l�R+LOveJ.���ޘ��ŕ��Y|�dI$�|z�墌5�s�A}&cȫ�S�|㺸�ǒ�IN�,�/�w��;[EU�#
��TE�֠P	�ی&����� �i�v�J8@���!�2�vT�������K�*U��� ������ߚEm8�S�za�2i��Ӈ�{Э�Х�^��[���޶Kshb��h�|�����!�njJ�W�;��埣��:��8�T�Ř�L��8����m���H鼅 a��x��,K.!Z�9�P�K��ѿ0��41ES�R�Tӳ��;��v�������_B�^P�x t��M�,��F�QX���SX��v(yO���&���a�z=�m�Ξ�gF���@��;��65�/�����nvZ'fmЦʦ�i2B2�,������[�2�K�z������������w�W����'�,z�1e�ek��x���JP�Z�H��=k��i�a/��X���BiR�=\�O���~��*_9ٔ^�f�ҭ �i��S�1�x��
{[.�N近~�رwVx&��6آ��o�⾛��~F��Ͳ(�~��3 ����G?d���%�Is��z4���ބI��3��]��`����wu8� ��p�8 �3�[ff:�����[Y���;>XMl�՞��>�2Zz����yݭybpy�X뼤�?z�Cxe�yl�V��ܦQG�0 T�$��@�Z�~ i���$�WdV�sG;���ڀr虶�aЄ�[-m������/�ˤ�؝p(����aT�����!]�����lC�pի�<3+�W���{qt��`^\b��j(�ׄAS� ��l��HMʚ+"������MJ��M�#��>�r4��X�T3������"u�,�儉��[��2�����<�|Z���XZ�ʇ�W����6�Ęz�(�ne���KL\���W�8+2�˾kkPBH$a/1���ۨ+9�v@A?�N�C��YD
 �fp��"���D�*ڗ��5Q���m7j�Z�V�(�����Vۂ��m��J�	;q)��?�Ff2�p�KE�'��C��e�zY.`-4��b1��YK�0�����""���Uhٵ@����7~ ��Iڪ�����;Ѹ%��ʣ���S����ƫ�o;��n�������Um��sW���J�nM�bA���ڡ���oj^�:	�q��x��[�&|�`zX�����7S���
�VN� r�_�O��T�hM��]o�{����y���!���ď��9�AT|��=L�hl�d1;��	�Q[�6�>�B��H�t�=�!"ca~G,J3n�0U��0���5��h�K��VȔ+�Л�'9e
a��XE�E��(�l��'Fg��\����(�qph[��(B�R�,k��9a>F�E���9C��b�̤n�l\�kY;���-�MeC�<\Sσ�)��hN1T]����p��x��/oV���ft�^�]CM�T7$����h�,݆Su��:U��MW4>���)���L'�D��ț��^f'qZqS�˴
悢��g)Gni�ÿ�Zdk�jj'��C�ޗ����8A�OCi��&�muS�V��z��E-̎��3��eUHp�H�=��d����"^;��`�����ʘ/���M2�)�]��Z��ě��[��F�sn�������b3Q�MS[� +j�V���w��8�	+P7���J�UGG5���-�j�^��w[�'�}�U�N��yH~IW�1{�4M�)�?�UY�D_T���nק^l��	O��/���p�%��z�� &
[To(�Y��A���e�$a���T�|����л����j���!:ޱ̆g�O��ݍ��<�ތ�
�(��=e�[��d�MZL�κ�K�8�
g���Z0ki"2�]E���jH��A�p��c����½�������5Ց(���� �'�	q\�H	���*�/�@�'em��l�Ɠ_���9�ɶ�&�b�b�l�ts�\��o���u��������A��f���w���[VW����d��5,��w~�is���՜9�C��/�B���5��i��L�jU~-���Gt{�����q�/Q;�mi�3G@�L)7~�r�YVW5��͂�0�'姭��(�ഉs�E�������g
ֱ�V�����9Q�ڍ��5�?�쮋\e�;*���!���>B 0id/D���xKᢤy�뽕^İ��{~�s�t����,AE_��^���U7�	���g�l������MH�y������T������S2�ɞ�pڪ���hЖ���&�����0������2���������8�У+u��k�0B�dME!	иr;�ԡ��д�Ԑ��7��5G6T��f N Á=�E�
��J�ƶ��+p҃�dٚ)Ic����[�W>���<r=�0��C�Y���V��:�����=Al��M񿁾x>�}��a����%Ǥ�@�,��b{` %\1q��F9��`��G�d�c.���ꧯ�p��:��~�À#�R��PD��Q�s�8Rc�څ�����"1��u�NVc�H1(���T��v���.[�<�,�������m��MZd�0�>G&�����2B����0���v.��(r ��
O�N�ԻJ͎c"��TU��F:�T>������W^7���\��d�F�-�������J�&�����r̹�&��r�3�c�xŵ90�`�$Gۜ!�h������C������Mo����#`�0��w`�Jn�G�2C�}T�IE�v�3�?ͩ���ն!p�d��5Q��_�����!%�R����1p��b���t��e@�jك�t���bk]U�/^w�@wX�)�ncAm�|x|��!�4�� ��ag�l��!�@[OMC%�]2�G������9oE5{��vu.߰�����[��|�̖kK���(�>�Q2\���a|m?a%��o���"�3��)fՉx�y��8�ǆ2�$W���a�#��HcE�K di�a�� �L̚�f0�(�@#?G��1�p��&�_�<���%Xmx���
&���H]�L�+iCB�kaM�;8�.0p��(�7YУ���-�ΙA,m�N����Qы�b���Gl�調)�f1m�%Q��a{旻� ;7� �]���uo�')��N?��e[x�i�����b�i�M�k Y�����D}k1��X񂢤x��C�o��/��_�Iye�j�42���B���9({� �_cY�cC4F��t�uv��o���[�sn����f�t6ts�$�O#Dzz��S̞��x��˔wIڈ���L��n_F��G���Jg�I�%dY��;%�Zy��`�W���ыc��Ȥ�Vw�7O�N�0%k��*
6·)#[po5Xµ�Hl�/o���Q�}<���a��/bەM%C|�k�s��K�x�Q�ˆ���+��3coplWµ�v�ͭ3�'Hq�27��yn��y��������6���EcOF�H��q���ϖV���AҾ�t�'���S�|' ��ͳ�ۻ��f;n�1>�x,�h]��o|	�pϨpM��/hxg��M���M&�񍵭^��j~���F�8b��^�]��I��I//��n��y�Ef6�w�f��Q�,����҉��=�Vզ��[r�<���ܴp�u�֎:BY\��;�^�1�����'�;.$�|qp��/��k�-��A&�ս�Lw]yzD'@)���v����X�Eێ�P�쬠��a<L�-\���c�.ę�鿔��~̋~����[����\W�
�0*����Ygyhj���q�ͼP���:�_ד��FL��0�H Ա��ݨ�f�y�B���Qg�O�͐ _�GvX� ��
�Oj��('i��%�p\��*J��J���N��mw4o�e.h�	i��%U"g�����P7�P�b`
� :�-��?չih����t�f[cw ��d���O���t]2�&AC�!OO�4Y�;�Y,�jJ���a�"�Y4���h'�Y2��R��׺���a�i��B�ק�߽UcQ�Ըh�_��}�Y�~��v��D���_/W��
Mv�`]>K.!��S�uN�j�W�D0u���lE2��8+6o߹�M�Ν����"`C��\��3h�W�<�9��s�#�u�nXF_�-J��6o��I�V,�<%{��5	"B�E�7o1:��CdZ��wD~�H��=BNT�|�H��ƛ����`��� A�S��Y��l� ��٬�4�g��t�GP���c
�EXPۖ>?=(�,{��$��cG��J���]L�rD&��i�l5��o��B��є'614�����u.���D<=t��p�6�Z��qԶA���F ��XM�L�^�v��x�k���%|�i�I���3�20���:U-]d�3G�;�E7�\"�X,ʸ�*����>�]}�|�m��jڧ��هݗJ�����8��^%Kݽ���$h�7���@�FM������<';.�-��DәM�Pi�3/I�s� �YB,zl4�Ž�5/�
B�,�3I*l@X����ǆooH�1