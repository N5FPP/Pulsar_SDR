��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY������@S�}��@jm�Ȓyp�w��G}���-��_	�rM1��cP�'�)gBq����ww�$u���X���W�7�实�ͣ�59�����l��xe�8Wf=H؎g9a����&�y���A��������G�տ8&��a�U�۴K��(�I�.(�����Mto�T�X��b�s KN�x�K��z.�	�n�K�1�N�*�>�P�C�g�J��b���+�ҫ��xfz%� 5��X@YЧp\:��^�5'=-C��Ԉ�s�A��4����
�<���i�!��i*Op����o��5RK��ee.� Sf�sW��d��ߟ�h��>?�&�'�=9�ы>Ue��̅Z�ސ Bj	�"�/�ֈJ���>O�4nym�6eY[Y��	���?MAx�'u���{�������sO�1С���!<_p����}�\L�Wd.�S������#5�=�"�7��|)Y�Q�1�s�k(�vݨHl����=[�/q�J1�^U��Б(u 7�ٌYb�_�#h;�>�JNj6���K�^/�5q;>��L�u���B��Ȑ����ʪl7�}��Ws������Cn�x���<��ם�.�R`{Nh�g3}m�K<��)4ye� �Z�s5�I5��Ǝӳu�{f�aPVsi+������A�`�)��#�|4e���*����~��x�G�ڗ����io�xn��?�y�&6k��(~�'���):����*�J��ѹ<~��!2�����=Q�.A�&�ئ�8��g�����h�ӖY�z؞��*[��(��-Qӗ}�d�4�F�������p�Ւ�f�a��X_�w(Y�D�/.� ζ�+�Z�9��G�]N��Ɍ�E�z!KT&�Ƃq˄q	?�%��w[��nR��0V���4��<@�,�Y\�}X�t�}�{.C��e��X������|,��(�����z,���k!U�������`����w�T@�|�S(]lP�B���/=r�b��#�'�-D��]u±�H�F�[{�VGf����|�3�S:j�k������I�-�����߿��btx~T�.�,��aG��3'�!PIO)����z��UhJ�L��Ld�(SF�Z<��kXe VXᆾǛ�lLr��u4����n+����>�3D��f��R��W�����%ޝS�R��k�(�@E��]�T!�����Cj�=dO�ѭ�lXJ�qU�k�xRN�.�{��$�^ʍo�Z�m�#��X^z�7&�3Z�j�a���	���9D�$J1TOg�P�N*(눴�"���&��bn3�K�o�@0��ʹi�������H�ɖ�:�m�]���_��R�=�H{OV�E>�"r��-5Zv˽�⦲�^���<�Jn>��[�a��xl�B(�R��ӆ
)�N���N�r�:�,��u=��A�-�e�/�1�� v
P��a��<z��c�]�Z@T�S Z�B�Uo/h0|x��BdWIŇ��jB:��4�'��<9~���$��a�ϼ�1���e��-N+�m�Q�!�� Y����:��6��w۳��B����'�Hbn>�2�|��U��>��+��MvV��#*���5�&���X��}� "��%�J���W(�r�i�`��Ɲ��K��f�]i'�?��=���M^��O�LF�h��mG:���.��>���󈲽�����[����/�w�>�*�3aǮ�N N��(W�j�HؖN&d/ ��?�����˖�G
ve��ʏ����R�c�B���2�4a�G����[����>�m��<��Z��O�U��e��y|������u�>�Q_�&qx�A�s��Ry���lbZ�.kf�:܀�9I�\��B����ٳ��<�\�����c��U�G�7� F~�S8�u2���^ ^�H?�k���j�l5�=_GR�ˀ�~d���O|�!�-�O$�Ѓ*1�����8�y�͑���+Ʌy�ioJ?�x����ܞ
���x��w�1�1h+\��{ �%��y 0+�)������.~^����� ��Q�!��~ȍ�]��G��������+?��N$	<��%�`���_���$Wk�����{�#�u��g���2��G������Teeܨz])1�ѓ%~�]N��cGEF�9Ps���1]h���4:T����K�:������ˇZ�q~��qi��s�t}�\���z���b2ߜ-��B$[8��D���4���⁋�`8�Ѭk��:�ĎL=tD��\����D�E������?�Q)�,q@R�R�I��
\��T�����8H��l6��l���к�1�-�	�|���L **!Hc�ȼ?�Q������~`IRs3��_a�>(�	��")�tڶ�GR:��X[���ՔF[�R�X��f[t|䬪9"�U<S��u��]/T���T�9t�'rOd��wGi��q6e����ݪ��_&T"i�1��ޏ#u/q���	��i���I�iPs�?r����y�7�Ћ˖�%�bg���M���5�RK�?@!N������0�yl[Ȳ��f��H���Da���9�.��a���ǽ���To�!�����T��.��(�& �5��d�6l��6���F���5�ލf�	)4�C�U�K�ٮ��|`���K�O���P�5��+��mD��j�P��dU�^�?�P���UjQ��|^/�����#q>����n���5>�TE]3������M����ZA�B�{s&A�K	���yt��a&6���ai�;��:�I���+�a����,6�kE�l <NOŌ�rײ�W�㠕q�3�1�V�`��Z~׶��Q4n���+J譸���|d�*W����b\&�)fy*�����2 4�=�$�����������×�[G�>��M,I({��W�Ҙ�A���*Ҡ&�����Ѽ��<�2��0='��>��>��%h��Q�'�+�pB��#g��~�I(m"�C�M�?,����n�J���J�i�s����Y�[h�Թs*�����Ȇq�H HLJtaY���:��
�����g�D��8»~�P�'A��{�d6�}�`�+�S|��p8��S�]H"es�`�'0�B����3��K�T�WG庍�UG7��1��N��G�������>�k��&����w��z������꘺��*׌ޕ!�J�^�9�1́_wc����"n��de|�?��5�<�a0�ɣ�c�dN����!BhzEvQv$�)/!9ʍ���Y�����i��`�!�����X��{�oR���\xB�_�:t�hD�>���~��*Ɗ>2��Kp���߭qtqx����[Q�a�T	
~˕c+B�=rtu����D�L`8��P����B6��G��|�B�⭳=5�%.T����_���D�D�T�̿i���N�Cd3��۫���2� 	���"�`����k��?��{�X��!�](�`y����2�ul^7r��x-�[�,0C�ٽ̀�������_����dۏ�����1�_"��}�iN��)�J�(Z,@L{}��ã�)�Z��d�<~��>���	��{ �C�*S�61�q7��������`����f���}�/�%V_<������;qhB���&x��	L�w��P�G�%m�s��#7��������m��Ư,�<SgOS����؝���f����dw89�$+�ֹ���'�k���S�܍�Ӑ�WA� ���;Sۓ��n��&~hw`��J��~�E<���~>D�X���u��W�l��o��K��N���Vn�YR5w�)?��F�os��D�	���;c���<��$��X�X�Ȧ�J&�آ]E���ټ7/׾ob�"����5���߽u�(~�qZ'�R�P���Zv��6�������%�:�\�ݎ�`�h �hH Dp���d;l48�S�-���6}�U���p[��;˙�sW�Q�A�Z�j�v88���~͎]ױ�@���l|����e#*�}�Z����~�@�䡘��� ��\SW�FH먇�l����m��ؠ)�V�m*�@L��=�a/6߻٪��R��6��3��k3�h�-���	I����,��y����Ǜe��N$a����+�K��4��U�}/U˃�������w;���V���F��`}���Z{<	�4�B3 :�B@�E^n��+����*e.�!]�uo�����>��A���	-����'��C���FD�;U�.p:�=�����?Q�}\o������[��	H�ލ�ñ�!�+b|�6)�?�r��6��[�{�z2vQ �Ŵ��ۙm��K���U��d��WZ����.Ƈ�+��ǥ����e`�I"㧖��|ƧK�b��lĩe�U���tDV����K�yK8�J��?����b��ǕV䔸��}�:*�"_�V ��
B���C���zF1t�\�0��s���Z����&%����U��d�6y ���k��p�h�y�+�7��Ts��@��$�zS�D��x�L�y����>�}aI辐����j�tu<w�hr�?$ہ�ԭ�&Y�X���.�f�Ϸ�޲�P	1�� �kQϳJHQ�|�����!��K+�p�ZX3�Ҫ��e�4�H�x�:j��7^⇻.lxXu�mvJ��2M��^A��{1s�ށaចqfE�s~Z)�'�wU9�W��{DU��dG52��{�Z6�8��˾k-�o��\cr�K�+�E{���h�V�e�Fd��ٰ����a�z������N��C�N|���@��w��.�j+� "^�³%84f�`^O��h��h���κ!��E�0���;�+�erg Ĝ+N�����m�����矦�)&2�U�r�AXS�{9&�S"��o8k�X�8$�X�t��� v��(�"��{�F/��s^���B�Vr�h���p�*��n�F�PTH�j�z�d`tt������������_	���������۾��̤߭�
��2o����ft�(Op16������j�Փ)9�Ua�:�7��$�0�u�V}�U��QNj�!�.q�p���>�)|ϊq�v�܈��T���L!��+�!�}P<z`tg�AbaCq<���U)N���>�2V�,<,�F0�A������^�Aq�l�a�$��,)�W@��̬ �� ���d%,,�=�.ZT5��=�%�]4b?�m�3GzH��$V��z�Ŀ�o��o��&�r#,�o"�2`A�tK���ek��3,�����;���n���Hwe��
���uώ��y$$�l/�gï8��4�r�M�F�����
G���5dKY��2=�Mo��-ۅ����$��H}"._2�#�#Z����|� ��J���<�O��F�$c8���	#qIK��w|�MK="�����:L�.�P
U:9�=��@2O鯔��-�#��>h�R�$Թ�"�;F����o6Z&7G�l(��R�kړ- �j5E�i�̫�	�3�r~�٥X�N(l� I|��M����hٴ�t.�!��z�@/��*�`���cS[�5>2k�/�W����O��p�@Wk��h���T�~&�ț���\�E)�ajA%͟!ߐ,�A:����v�=E%��=�R�� �?c.t�4�'j�w���_��OG��V�~(|���O?�[#)g�������+Ұ��Mh�o��P_���`x�9���е��]��9x�׽o���`]�:0���2��V�w̲�3)��Aĺ��cBl�ʏE@+k.�l��"��h(�T	�����N7؇���Jx�m܌���� �+Z�6�0d˱h||M{�YPo�ɂK|�������UԂ]���"5%��t�Ux�e���hF�R�a�t�=���]�kK��dR�4�/��!20��������zu�1��a�)ܥR��6��1f/��Xʳ,�4�A����y��Oǲ�h��՝7�ԍ��`eKD9�C�K���^�H{%\�z��g���(�[�`�a�N�-񕱆XɈ��#.�����z߁���_%���$�	��s�ٗ�f-'*��<�ah��<�*���)@i�*F��^�{0��x�g
u����ٶ�R:~��[��0ӣ��}z	�/�Gנ�_��Y� �L�W��I�����ϦP��x_��'��w�8����볃�ƞ�v҆R��:V%3��tFO=?�G9,�f�/�F^� ��Z4�L6q'��-��<�c�A�9���]��]��N���{�p�������Q!�ٖ�hj��C#�acdP�2����8Dkk�C���S�^K��@�ve$S�4*xhE�U���e:.n�:�KOK(^B�#���A���s�D#T�����i��͵ �QT�v'%f��J�Șu�t��mI&%Z�'i��|�'���������i�(I0#���B���`b]hp���Pk�3��x|���Rd_6��E��ǆ��b}�*O��:)	�>�_�Z�\�=�ķ;��I5��'���v�r.&U��0Z�7�#����[m	o�W���1Pۂ����JB�P�x��Z�����,w�4���s,�j�P���\�5�1�"\�g�i6���kg��km�i屦����a���c)���r�ib�|'Hr�����#JQ�IAV��@TUF�IC����w�Y_\��6�G��y�6Zܤ��;;�H�'�J�9CH �}�(�m�\�8��`���{��IH|���bM؝�a�M�7H��5'�cd��� PeȠcm��b^���}�˜��<<�^)��t��,�[�sV�]x�A,�c��s�6�>�)(H���G�}�}�a��S�}�m��RQf��t`lg����{����3���,!\�&]jc��Ҟʤ����X|�آ#�������o|�Ȏ1 G�ҏ���u�� �i�{욹�xH����*���@A0�D��:2t�	�;^�gt5%T���0iGG�w3��n��W�c��J��3�T1|���U��Ȇ��N�=Ő��l}	G��+����a�Տ����N�ݠ��%M�*�J+f���;�I37%m>����VA��rG�q�ҟ��U��&���E�|έC_��/0)��-�&X�n�q_NoKdK����H��\��"Y��ߺ����.~ڻAm!�&��}��S�]�p_= ?R�"��=�Z�,�!�A�Z����G�H�z���TeR	�<���/�4���� ��E�T��ԥ�@���@��fT4uU�W2�w8;X��(��e��C�.��ʆ��~~@�K��C̹�F���љU�N�;�Hwف~��q�J���n�h�'J(�c�m3�4����GI����8�?h�s���v����~���y�)��<��>���'S}��\u�,#s�Ҩ���c(M1���Բ`��G8�U��6��Z��kF��~�+���m�5jZ�X���"��(ϛb|������P�%s6>������x�j��(,@�1�::�Z�M�PA� ;�3���
�x|�(�1`b��;��B�^��e�������#@���`n��-��dI��f�g�}��ܔ��`c�qF��*�=JK��,��h����1O�����*!gT²d�;(Yj��k�	����*�:uE��I�K�{�߅KK�7iC��0 ��
j6�E�y���{�d�(��L��'n���[B��&���X�@E�;��Q@X�E���e��c�~�d��V|$�a+���O1J
9�(�o+Ɖ��4�����H��>|`��h����CRq���6.朠k'M��
�W����L�1�#���ԏ�|�H���.�T���U��\������x~c�SU^�D�2������yv��g&��/':f�0V����[��U�G����AEχM+b�&��t�!�3��\��_8�f����|�#�#��rS���Tz�5Sf%���/(-��H_��
�����t5N�Z����aq�P�'���g����%9d_���)tY��3(��5iX�k�u����ֵ���������� ��L�F���XM>��o�K1�_F��A�~��b�O��Sy�����:I��Ȯ*�x��<�H� �� ��@"�
e�㫽���噖YYY��2KR�u~!��/VDH�T��!Z*�~��=�x�Ww[��ϡ�����Nl���-�.�U(�jV�}��Jw�,��Cd�%�e��-�پ���aa��ü���3����ǖ-c��8桺�0ccN�@��7��O<[�
�Vki�ݡ�oNJ�n���^��ݎ��2�E
mʏD*(ӆ�Q(Э���%��-�:��`ڔ���a���7^����hK�R�C6PA#iӀaH"5Ϣ�-?��h1G?�R��>�; �8j7�Z�D�II�22��X�
{��b���c�����5�?�ĵ���ǂ6u`��c�
�*�.���hV�l�B�;o�Z������Π��pj�tu0��P����Ĉ�ӕ-��G��ӵ^�3���p�=�!/T;VuX(&�������X�C�Uң�&�5Gek�w�\��Ǿ~�Jwhv3�DK�:5�{��}E�W2T8�<=ԟ�
��tD6gN4�$��z�[��y��l	Ϸen����`IH.��h�s�r���yDs�v06��yW��b�_���hlH�f�h>��-~��|��V��m�U�ter�"2.����g��}u�w��O��������$����u<�Nn�w��@'�*⦕TG�=~vY+>+6Z�"@`��ۣ��7���:Q�N'�s��6����F�H5�6���]d�!�_�ȷ$:AX�`轝Q[&v\hU/1�Pb����_�L���N��l"�<�ņ�u��Q�l���S�@����G�	� K�E�zJ;��Of��Ԑ����{x_O�� =O"8�!1����=P�z��>�`�iT��я���p�� �7�y���&W�Jΐ����&m���l&�s��������O�Mi��͔�Phm���k�+;��~�h�y��aN�ٳ��B�4���NW�)}6\�|'�. Vn�.Q��e%y��f��5��Uxq�O�nΤ]�'Ԑ2�s׏�*=dX͵
&��ZzД{M,ʧ���iUG� ��_�7JW5M�.`^�܍�)ؗ2�7�\�4������*���]����<���x��Ҵi_��Ga߼{?�a(�0"�u�/�5�ږ\��H�y��������u�q%f��l�8�?�Pn�}X-�Zo	�y]{����
E����ܛ���j^3z�ds�f?�� Ēy}-��dP<Z̳��\���됚ãd���Z�A_+͜c�����1R)�Pz���f�ۋʻ9鰍��^���Ďɶ�X��Fɡ�����j0�ҝZ�w&!Dc��[y:M��[�Z�4��ou�n�N\1ݳo�_��-q� ��R=u�
,���M�Q-$�;ԧ�q�8%�I�mQ,���MW��H��&��#�g���)?$�'g�gy�͙��s�y8tjM!(�hޭ� �?��{�@�B�Zw:3���i��wN��u x�E�:t����@��CF�a�,;-ʢy�U�8���p�+�jt�[���*�Y�E&������Hu^�f���H��-'	Mߥ4�!6��W�ݙ�q���\���?����_ߋxA�v��<�!��Pyy':~��:.�!(bN�o������,y�� �Z���e��7|J��>ǝ�[q�'�۩�wV�ؖ��O `����0�JM�� ��Au�q���@�K2�Cp���5� ��a;��Y`�	�+#�g��.1?]^���Xk{r@!��_��k���8(����x��7�=�o���~�t!?�� -�z E�l*Jh� ��9)�gY^D����W�A�U�\y��a��s�|��f Z�"���&
i�3��E`���k���FJM�	��N����T^�w��OR�'��v��#��3���H�G�1z��x�"땸�1:������W��+��-)um����$�
��GB��
z�����LqQ�������c�ZX9���c���rP����{Yn)o�%�ӮL�m,�����`&ͱ�38嬚��V
�{R-��w�xY�^H&��k�q��;�?3z��g�a���\�I�;אT03�ex�߹��[��}�$J��և��f�?w��qX����N`Y���ȉ�.�U�6qFc�h��1/�Đh�,���3� ē�?��+�^\[]���.�	dұU�*��F�Hy�	%��hv��sR��7y@N}D���a[Vs�L6�
k�G^�(0C`M���RN���^d�c�^�Igpq#��#��h5�x��[��`k�G���"�pfZy����˳�rfoV�V�Ҡ���t?y�o|,b
�#t&Bߎu�R�$��MJ��K��-Vi�:�	_�_EG. �33%p��
���k!����bjI���Y��R��G'�yC��u���AR�j����,茂��(��!�����,��hi3`9/�jëUd����p	��s@:�u(�O�I��
��gTJj�P�4Lo�G�il��M*/}�j�{���n��*��*}3�I�����2rM����2���?�a�i�lv�C�l���}E�7oH�2�.QOk��6,E���&t�����V�M:-��C5F�7��2��B�R,�W���bEz��i",�m�U�����?���t����V�j�vBg��\�z��@�p�0dv ������9��n�B���-~�N��zң/dz��4�#ag��L�i#7�CNgmGy��-gA�C��kQ����<͓Qh�O$hխn�L�@���k����m�����Ju�ի�K�iZ�C�����H�z�->�w�l^��V���u۰Cz�9�Dt�\���6i�#{�	i������+tO���MFݜ�m�K��bf�3٣ѾIk��,y(�Zn��;�4�;M�-ϱ��*�1v���N���Hr���'I���s8�vݫ�܁5��x���8K!� `�>Љ�ttB8�YdF3���:}���cZ�v�m
�h&��w�F!:��ݘ��S{��B|�8G\��r�S3�Y�S�c��%ؖ�����)�b��#�x�F� ��&ň6�N!��|��Ǩ���؛%%�o\Nn]*gw�Ʃ�x#e9T��]��)�G�%R�m˄��ʑd�
�
��tVL���Rb��Z��5A�|�Y[$�`B���ULY���GO �-�\wme�l����g���5�!:*�8-b�u	}�k-��͡�7�\�C�h9ﰪe]u�v�.>�0��:̘��ῇ�r� `&��
G���Kc�zsސO�OZ�����^�ƒ�2�۽�]�E�Wq�C;:��
�Aƾq�Ŋ��q�>�<��e�pW��/#�	�O��K����4ܗ�kE�9ԙԑ<���Mv�ڥ�g鏇�Y^��P���ƿ>��N{E��w��S��eի�s.�?�dTV�,9e�k��!�e��*w%gL���MΧ�����C�n�/�D޻̴�˚�~��ضW�c�L*��ӠOm��=w8���J�~�
q��?n�T�~�uq\�H�j���$���k��/���`|���,zvoy��^�����s�ܘ󩵮c����q�u&Z���⯨�^�3��s:9�,.8��o���Gҙ��{ln����o���yJ7l��bM�!o���NԅNe	b�Tr���>�;:�/�uX}gf.G4������ ��w7@4u�A�-�]�PZbv�J���H�҆w����J�Erˑ�l�8���^,ޔ� �"�b$+�4��9<�}� �w���#U��n�7"͵;e��QM�]�N:'X�@,|�����ь�	fAgy�4sz
�l��SU#�P��Y�j	'�����\����o���ϰl���:F�K�M�5���)���Ԏ��`ܩ��x�Ԙ4�����(�_�3�{��ϱ�O3�L��aǢ�uˊ�	�J�"\��F���ے�l������p��%���?�"E����������ƢL�q�h��F^�u��e
�B��oW�cG�Ep��	�RY� ��m�f�N@�'���jx@�8j<s;Q<s?O���qr<�w��{p^��~͢P���x�`�y�U�hv� �c"(�j0�k0�]D���`s�+n���#���e��<q�;��\��>D��aL@�qʯ��VK���N'�j46#��s^��-�&꜒O�W���\b{���n 7���b����G1������˷�my5�n��mZ�6n�����|��͉�ϯE&��:�ۯ��M��_F >E�9�:a�x�*o8������ø� �i��ܻ��fag���-�����;v�c�|/���`���v\�m}%�(}�T�e�ݱ��Yx�S$*�����f�$�;����-P�_��=�H3@T�w0_,xVy]�oo��k���Zr5�#�eǫ}�4�%������<��wȋ�<`"-rI��ަ� �V��S�����M�pD����hKm	����U��qa�$�t��V��[<$Y�C�=x��
PD�W&��O��q4�J�A}q)�٪^#���ݤ���h�l
����Ql������; �e��0H�t|��"oU�މF��� �KvŴ�v�(�|3=ϵ���ʖ��ܜ
ϷT#AQO���p�Q� mtw�h���̠v@�����s��^"��2�n^�r���������bu �G.�6����4p�CWu���%,~��F���	iӂC�h���WI��5A�OĩSaYy�a>4yT�0��TM��,�*��Mo���L5kO®��R�/X[� 	�'d�J�
ǘ
��<�_�7;�w�֨4�%&���X�kB�W�S'H�#�o@̿��P�JG�y	��W�(
����Z���V��	�H[�Fz�-���v�um��A)�xOh[�Gb�&K�3b���1TpZ)�,�q��"ݓ=~�]�}k&�{>/�O}7	�!�A��d��%	�N��U)���.Q�X�P5/M�ps�6q �n�0\Q^�R͒r��"8�K����#�JPE�g{�(��cCD�y.��I��� ��l[�:�Ob*�/�挌5�A�
	��=,J=�&&��rN��V�pl�HxЭ��sTE/�Gb�;�DG,���z�e�5"!�X��S���^8�ぃ��{�������v���>��2̌���io��e�C1IA�M9F������<1�ʹI$�� �X��1X�c',��]�s7��(t�CB��Պ����@���S:���3�e�e�U�K�`H�"L�^:D�P����wډxoaK�صʏ��C��(��d�P�Ws�v�󽎿��b-�jD�qx_�Y�����M~��`�~���S��ձA؝�$�d�h��PR��N��H�}��C�;���o�*o҇�l X��أ߭��)� ��*�N=�+�|L����1��HɢKW�����};������I*��T�d�ҷ���g����f	���{򩱵f�ׯ��E��8�A#�9���OR�f��s��d�6�6u��c�If�a���>0�1���`fx	-�(����1�z"SG#��Ml'�&)3
p1��Xpc��+����~7��[����}�>ˇ��m���06�EH�R-uk1M��֊����� +n#���ߴݍ�k�	�gBO���f�k=P�u8D��.��*"CK!�Q�s,�,V�+$�o�9�Ϸ�d�����(��ό*�A�}<���ֶyQ0����6��D5B�Hf�F~�Z��wY��D�\��=����v�r���"�7��QT�~2jjmF��ı3��QA�E�QIGt�^��o$��[��HV7�k�%$u�ړ{�
o�@W�<�զ���k��$��pS0�w_�5��}�8ز�JC���S6,c+�c���7'n�P�e�XX�2��6�b�y_�)I�ѣ�ԁݢ<7/g������UY(�1ZwUZ� )J�)���l���>�ɥ�wF�,����Oh�oc5���% �O���Ϗ������;g�굨�A5��1�����f�fH�֗�*6�y�;D�ƈ��g�VӴ�AGq��!�W��+�b��wZ�+�ɻ�vjH!�.n�^���K����ݦ[}:8��h���l8�{21z��w�W;Z�u#�	��f�0��c��}@� �,�C��Z¸�*}�	Ebr�����I��5ja�"_g��< ���%��ƍ4Cj3�f��Yt��o��͚J�庥yAVw�-�c�I\b��Y�ˎ���d�K��V��?�xP�|�-��W�{�ۣe�+�/�[���HǁP.j2�C�ro�6�v�7Nô_�Q6*XA�a6G(3�e\T4�45g�W���U�t�\ߕ+�G\�<����8���?�d0x���?�2U���6;=Iu��t��e߈�~R�^C蓟3X�v���t�,ɷJ�5Q�7m�×x�F����Fh�ԇ�
�E��nl���Ԣ��[KUGΣGor�í��ڂ&��c	����&=OH6rۋ���%��V�m>6�$'��[Z�rʜ�y�+�ƅ��?�w���ٟ�L�R~T����8�:�S{��i�7Ǫ�T�!� ��gO���Ɋ�`R����:
�4�tfa�U�Z/�G�`��MV#�������O:�5RGВ�Pl�/��Kk�p�g�c�?|H"�V��X͍+O�f�󅪋s��d���f�m<Sx��t����zn߇�B���T罱��A�:^��{:��Qq�����S'�xT�F����{�Ϋ_,4�����V�� �זl��*~ 7ܜ�1����ި~��޲�V�I��f�8��,3����|��mb�RDݚ�ew�Ⱦic� K�6f:�R�Az�5����ήl������� �@"�l��s��g=|�]������;
GuW6�����"��n�?wy9M �ek���O�G�Oj"�EX�
 ��&��R�'cm!���)���k�-J}oO���Ob�M��zɄS�x�?U�����(���+n�	ؚF7�y�Z1�<�N��e�+FQ����q7n����4Dn魢�FS��zI�p>��t�>�$˜1���/�ol�`}n�19����X����=��N���[ޔS<��'��g�.�ԙ"#�B[��a�϶L�6%KяO�Gm
2]Sl�OW�}��.(����]<�ָ��`JK���q���c�+�����[=��%���u1�ʭ�������6B�u~\��!��?�� $�CA� �e}�Y>{�n�Aʼ��J�)B@oA���$��v��j����.�J',�K����[�'��oaz�n�v�����������]�a�����ԫ��ߋ�j�^6���H�R�ӹ�U�vC�k�<��W>7Ew̳6�~F'��K�N.jJ����'e��8�Fd6��E|os�
XeP��z:3��7�fov��'%u�>$�N�� �,�=s$�)L{��}��`��ћPo�~�<
by�������@u������?�/�K������Fg��<zQ���Ř�Z݈(���N�!]7������ik5%&b����;�0���{n�b�-�y�|�q��O�\5��t;v\y��,yQ:��sPԍ��K�u0~d#�/�xr 2����?�|Ў�A�9kl�'�#���8h\��!�ܪ�9�x��zK�Uy~�7��1��h��0I��/�gX9E
8g��E���rಛ�!���ٓ�/Zv�P�$_dkx=����y��~��Fe��ί�h��_�p�l'�j~�%+ZH��2�G4<T�J������M�O�^��V�~6y$ 
�8�!~P�EnP����q���rBx�EZUu�&^]N���K�J,_�R6���#E+!P���#�I豲��ó%�%�����xip�69u9����|�;9��<��Z4������J�/�b;�*�wz �Zc/	�_7�6Fh�K�m
��"��e�A����Ǫ=ER�s�"J��P
���>xY���]��W:��X*���Z3��0cB��3	�������;6�è���ǖ���]h��^�;8�Oo����̓U`W�xo�BX�Q��|��'J��8��ds)3k�����8�	���W�:�h�w���U`k�o���9����H��O:7q:S(.�KF��*1&�spܖ�ˢ�Fۇׂ"�gR֞}A�1S1��v�bF��їP��<��%��kVJ�XJ���Ξ��P�$Y$3����"�X�yP
�L�Z�ADt�K0@!շ� �'Q�Ғ���X�
�q
F����g���FnAs*̾����ق�[U��q�ֆ�r1�n�4 ����aF����ޅNYX<���D��w��~��[:o*��jWR��� �
�h�7�4U�m����%�vcc�}��46�5�E���+U�b�ϸ]��,-�rJ�x�^�d�a��?�������u�/d��=��kB��j\gN5.M��	m.@5{��CL�U��Z�}�f����ϋ�]���,�E�B�L��E���>�srn�����������㞊S�*)�Ub�	lbuQ��O�5�˷�MT?�l)�?xtV�%a+�}��w�؏�jU.��������o�c��jc�)�����4K�nv�<lq�M�L�����$����	#���7lrQI�����N����8�5�
}p�x��g���{�~�Ui�9ӯ���=��K�(�y�.��K��]�l�
��@"\�S۰����)`�`���|��}~�sT�� ?k魯#kź���nA o��j��������P��boee��G�AUB�-��<igs;�o�Z�Դ���]!�,(�\@�P�\��ʅ��y�gr�v��+���yw��J1[vL�NP���>U6TIJ/����)�h;h}��jVy�����C3�vKM�NPi�f��|���B��A���n�J�}��ު鴷��JAk̓�"%}M�s�i����(N���n���q��io�B,�ٱ\g@fWHԝQ	C�!4��fwW�.���6g���X5Z��Rۅ�f�?]s����m���W��f�Xn���w�8,���#�k���nQ�����yvF�~ɹCࢾ���+��x5�![�|��ǐ��Z���j����ڷh��IvW��tK+k6q�Qtm>�5UϚ�W�>�qB�X�+�����0�m�����������qE�5��B��x��~��!r��K�;�9{^k�cQq��_`�D7]�8?i�!���wl��:��w�S��n�,��@N��P�Ve�K�E�D�K�	*S��"-���uj	�j}T,��=_����d
~�Y��2A��!<�B�lg6��&��?"n�4A&���(�7T���RN��K�4���^4��:KG�˗T�.��<�.��E�䠔5VR[���ˁ�n\�4 �dg�X��zي�Tl 15dP	1�u6u)"55l/7�%�E�[���Z�����{J���@��G�\lt��5�78����o�\(g[Z�uV��(Cw� �*�.5�n�����C4ŔB�0�('�de�9Bl�m���5�.8�<�⁁��V.㊮���z�ױh�p�?�q]������J(�_�C�_�+���r�tFL�:B�!�(-�Fi:Lٿ�r�L��ZY��j�&�Rq��S&���0�g�͊9��x���W��j���.
�h-q"�W2���7�AZ���Ĝ0�:Q�ۯ�<@\����*Rޚ�/���8�����l���&���i2xo`�;��m�D��k��2�������C�����T[�D�/~����N�֖�/*[���P��K�d�C:z��Q�dz������MOkR:�P݌K�R�Rh���5���{�-!?"a�񀲽u	y��-��ԄE|�(�����t)�L2M�r��K8e��gV�ː'���Kc���@+ Ϙ����P��m��V�3*�V?�*��[���O����ini�zD�x&b�IQO���� �";�7��b������lj��a&��}GM�JK%�?��d�]~��ܞ�ș�I�m�!?a�����[5�N��SE�F_>)�g�b����=����P� e�bӧU�ˡ��1G4�+s�="�b-&�.������G���=v�fn�(��Ͽ]��5P������/:��{雳�z�S��ot�0P�I�*\w�}V������S��I�_z�6tΘ�,oFΐ�&�����I�?��ݑ��_�A3��X��h.Qݢ2�qi����2��x�MƢ3c��~�%���~:�9����7��*�O���
�e;*N�,���V�`����kf�zn�RiGS(�����l���ygQ�4��������۾ټ�����?oZ*'6��#����9�	���L�V�t�����2�����ՂM"ҪN�a�ɹF����l��$��@����Ln��s�C��4����D����	X��o�8���(�v�oʙ��R/>&=%.%�7d�@:��p��y)�yq
@�>b=w�M�B?"�!-����fT����K��e�����&0��fx������X����Á�~K�e ����k4*�s�n����4�쥕Y�V��G���]p�l����Qa]�K���֪�����~X�v�"�ۂw�Zi<�_�S뼯䵧�Z{y�)ß6�Y&\�08uL�_W�'���
��8-�:��/��D�Z�4o�� �6U|[���,�����kp�����L�e�'a�U���f�2~p3ml��xU��;�\l:
y�W��	%6�	ކ������u"�T��"yoK�Ch���(��Ł���dy�\4Y64�`���R9Ͽu���>���CW�-����ԾƶWP�%�j�h����js[Ց#��6����o�
��y��@Y�7R=��1+ZHg�%�)8J_���l[�� i�M�S��5��y���z?Bh���bCA��a<�A�S6��6���y(��V����T��S�fĵ����[��t0m�>�e��Ȭ m��$4���K�����Pl��*����A3��a�&����_�V�x����'x�7���������R�\�9/��⪮��������B�+X�,���Q:k+U3EN?&�>���0�_Ųi�ZM1�s�5s�ڎ�0ڨ�{�I� ux����̎{���L(�o�<�H���i� �l�&��U�MU4���I�Կ���+[���Ϋ�-��5-��]+�^<5XJ2]bl ��셧*q�^Ϧ��Z�_^����N��ło#��l	���@�F��(@�1h vw��8�4�)�W��>~�v�.��+Y�[��/n&���i]� si��X���:1�ZҌ�2�����a?��à��E+�:f��ɛ�@�z
�ֲ'���C�je�?.䋉4Y a"�Q}s/-�|*U0ܖ*Z���%d@�7hr9�5Cq%�^j�'��U���W�j|�9?���6��j��5@G��B�є���=j�����:��D� v��i��cC>���~#V�"�K�/�B*���V=��Wߔ�Ⴁ��p�7���<�l����c��e\j[o�p�o4c��tkƱwo����XgP��IY��O�1��,�+
QqR`�(��[�?���E�jFӡ=��zFG@�����'=8�;�X�&�zdG�3_e�b�M����
��QKU�'w#�_A���j<�+O�/�7h�[\�����΀s����"�����@�R�e$��\��d*N=\�%SAI�x�S�'���$���D�TM� �3ta*�tb ���ټ��d�K��P�Y�0�ު%�-��;�$ˬ#�u�T�[?N)n�9�D���u������A�ՏXa�mٛ���.�S�@�d0X*q.�����Z&²�O���۸����b��V6H<R�8�`��mkAm�������Rd����B:�78�F�&9�){�}".�� ���VD���j����yjA�5	�yw�ǀ?,�=��A�b�����\P�滩w���j�EÛ��=���o��7���'~����|��
�1�p�.m/�!�I=U��fb����m�3"���sfk���o��b����+Z>�E��+���9s�.�����ǈ&A�p��0'I@V���
C1˹���h�7gF�s��!,��n3���zd��$�񘓌"�0k�$�8tΟ�R��Չ�ɜ���g�J�N�_S6�Ԍ��e�1C��ª��w;e�����WuR�M�$�������G@+gx�+�H�� ��'�0+���Y��&�F���f�j�vc�Ш�_)mG�cl�V
=��܇����訾s�IU�_���Z`��A�菆G��̆�S�	��٪y��M��D[��~C�F�Ы �l��p(�k�lƧp��l��9��� �W.�
t�B�!M�-�M{ta괥&��END-��=Ez(T��}�NB��{ ��n��5�8l$�<�����_;��q�O!��I�q�-鏕��QP����:^��Ӱ�֔�n����+9c��&��=ꝟM�o'^���ݢو��ݫ؟�Qe�����g^s�<����J�૬Mq� �aP�{��y����D[��i�L�
�3~C���Rh���9�S!m%����.�h�z��8�2���>"�	�!���yk���ej�%M�}h'�?�#U���L+�ps�,-d�Ɍ��r\����+��;�v���	�ĉ�4�]X�ph�p��q^>�Ae�E����\��a��'�E��vl۳�� �&��_	.E�����٥,	��Q@XM�X�w1���7���8A�s��B��s%�8)S��
���Ǡ�6亭#����<�d���;�*�+��KBe�e��E.�xȒ.L�Oj��O��K���_���A�<�4"rݧ�฻�"��֧�6S�ħiI��
��"�F̖I������(�̉p��}�}�.U���
���H�ʲ¢�jh�M!�F�᧭ϫŐ�go��6;�j�I��ۯ`�������@'�o��K�y���6�����][?*���o�*��g�[�Y��R�?;�&�3꾓���~-�֍��
?�W���N=i�(��p��B"�2g�)�8W�Mp�Y�'l^n?K�IJ�RR[%���
�R���"�'���W��z��>�e3,C��Τ�)�o�u�E��� S|l=�6�_ς�c/�~H]��G����Ў��	3��[Wc�|��k("���9�㓁떖�5_��N�0%�K�D���ҹh�H�`G~=�];���+��Jv�Z���H�O.�)�>
z�g1l�+9�}���l��'�*�	Q���#ӡ��0f���S3���8�{��a�����w��>�9of�TIv���";�'! -:��RyhB8>�''�B� ��z|�Y�x�p�� ��ro�xF���YOǷݜ�H6��ć��'����P����j�>ۏ��S�nT՜�7�+�`r]U�-��(Ă%q	f��ŀ�����޹�:t�d$��Dd!�e(A��2�b!di�֞T��|5	 ��˱��G�*��ќ˻�P�B�l�SںW��*�����
��#YJ���#+��D%��t�H���7�F��ז_���A����=���F��B�>Bz�S��LW�]rC�C��E��+Y��]1�r�� ����;�]!T2�S\si�x��P���2�rhP_d��$���c��1�M<Y��3	�)�J������	7�GA�$�����u�^U���v|���x,z$����W"@����)<ш��Ǘ�w�)�L��?'�M�H���d��#�V|1\,����Z��ձ�ʂ�E7��5~�V�R2����g�\�C�V����H
����͵4�!��)y��貪A�Γ�Oh�߰��ct�u��޿�|0�����  �ը�>�8|�*�V���d�!i��;і `��U0�H$��h<�C��ߑs�͝бqd0eY����X2��XLY6 �Ʊ�dY����HH|���\��,�	L	�1�Y+FD�O�w��u��!f���[��(��]Թ�4lOW�!��ס���ҏY�D�|L,EZ����f�,�ec��)p���<�w�8��$�?ɀB���_�z�9t�4/�Ap� �.�X=�f�0��*]�5Fp5GV�'B�DZƱ�2Ԧ��晳�Xۤ ���L�&n��f�f�s�c>$�m�77��DTZ R9��=s	9� fiIKǹ�ȹ1�̀
|!���S]��.4�ԁ�o ��Ƹ��y��E�zM���]yf�5K���������/����H�	Zήo��ꋛ�(Һ�A@�-�������� �7|�_�נ)0����ʹ{h�u�My�l_��c}���5�Փ�K�߯�	U��L��"�@�!ɣ�fGd��\��f���U\�'>ۥ�S�R̘���u�2̉���׶�%���3���*"�@h�Us`��F����5��$�։��5����U�%��q5\�هc5�����3�Q���Y�/����l�N=�%ڷ= ،8{?"0�����{*�Z8�A���P���:e���U���j\�?Y�T+o��Ŋc�5����@��j���$e��b\� Z�;<
�K7�+ᦑ٢�'�^s� wC&���#�!I#3����tHY�܋��A!�%�����M��ʹ�B� ���V�E�p�\�E�nV�O4W��jץ��[���s�k����A�!���Ġq\~Q��O-"�m�[Ɇ�$g
�?�.�%�$�+��6��.iǵd���}��dC����4��?��o2��5�@��e���\�1�HL�V^%�W�W��w~ Z ���d>+Kk�"�׾�������4�m 3��`Q=����3���J����&K~8�ޢ�H���1�TP�b'>����ֶ��Ѷʹ�L�T݊-�&K8i��f���?4�ܼ�1/�b��� e/v�����a_��s4�(��������I@���r(�;��+��Q��稄|  �A_�n)ѭ�������/0�}hP=��'(\�(4�O=�c8��'��E�rM�1M��xx/���m��+7�i�6@&���;f���>.�tղFW$�`��z���f��H4�#]Z>�i�O�*�;�»5!��o��w�݇%�F^��̑��x|�g9�IP$�)d�$���uC�䚺��.A�׬�dnz��Eb��n2��y�W�
�j��?zrb���!��pw���t���X�)����t{��ϲ4Wͳ��bbF�J�~$��� M�=g�X+���j���p�Y{i�g��a��ܝ��!�5�/��6޹VJ�{�)M7dk��,���/;Qg��-�(*�8T9�	���8���t����t�J�f\�M���v�1s�h⩚9���+;7�e��ͫ
�e�����-^r�+%��K0S��d�n È�j�p-�� }OL`V�K�8Ε��"M�z~�d�8���y2WLH�rM63:��yWj0����(^s̘��E������jukZt�ٴ�y���=�.�؍��+�2,���=!^�%r~,tje�R��,l�>�D�?��E�/e���l��ߚM��Q���@��,k��<Hl\�8�=Bs��Dj�
��~���
}��/'dhۀ��\jE+jl��v!~v�P��{�LM������2�2ɗ(�&%�>Y�ֿ}9Wӗ%���~jU���%~�M���Z���5ܥ;�|a�8Hw<�k��xir����T�l3�G���˞�DC�}u~���`��bB&X��S�.�c ?~�{�ʃl�	:�7jM6[�9
;>z ��W��]��l����>���/Jښ��i�8yK����a����$��9MD�`�ͥ�}\ϗ��޺N�R6C0��d`��D�)�$���Q>Zj���y	�	��j�8j�7�GX�.#p蠮�?�s�"�ۉ�Aʽ����{�n肚�Vo�m�gG����j��c��	tBl?/�H��Ih��->�ӀOAX:��%���P�����⯆�eBb��\R�e�*?����C�8^(����'�n���Q���J�[���BcNЏ� Q0�y�~��d}��=]-FI��"O�_e�8s�hf���S��8����L��	oU���;s�6�v���'���?���o��'��<�R��mbQ��"{}���|�fe�3����C���<�Û�W�������ir��R��%��Wy����Vܽ��QY:Kݓ�0:T�"���7#�!�d�b�ߣ�\"P�|%�Q�G�
�ԍ����3�# ��ݑ*�z�èڌ>N���Ә"�����9x��n&1Ǥ7�'�2�.�<S�^��e��;�&��#��i=(��Q���.�?�O����ֹ�.c逪�Xh��q��y�m�T��}o�3����ŕ��tiW=�����X��J���\?ZI�
���eD�{&�a��E����O
W��@Xs&��	n
L�;��b�� <y�W.��#D_`M���)4�"��{��6T�:�H̘��=�1g��'/g�
�UH鐹d%���*���Z�)�r��Fkr����S���UsgP����%�K��������I� ��'�[p�B�"�#���I3�Q|��psXC��~�ɪ�S7y�{�xSԄ��7��@�a� K�un����i��5��Q/�/Աć�S�}�u��*<�Yա%��� �<W`Q�f5���"�k{��}Q�Y$\zU��TB~�K��P"=�Ƹ#�����Օ��oRgm&��|s����|mQ��M����4��5��W�,?H6Nm�V��ssq�2df�񸾡p�DI�5��b!�����Dݣ4�$�[@-g��w�U�3q>@Z�og�I,m#GU[�:��H��U���iv����:��w�V��o�s-����:�e`��hs�	��	���*�#y$J�){ �HK����U����a9�q)����cd�WߔRt!��*�J)hpq��֞Q�4䗥�	9X��K�79|���"1��D�Xu�oxu&P̘>[�;���T���NV��)m&x²Ta��G���{14v�rfp�cws�	@5�}񥪟��s�67�����a��ύZ����!��Y�^�0V���n�����+5�v�%�Z�q��x�Ťd��й��#)����=�h�����W;T߇5�(��h"�J�	f|�����#:`\��P��d��1�eڐ���1��bGc���k�?�j��� �k��Ƭ-iH�'��!���\���仂�i7\
��f�R��j<��?r��e�4�(Ce�9��O����ΙB +��L˂�_�;Q�������L⯐�P�5�~����ٴ�$|@�xL�C`�1`��ı	���R��-��Y�Ѻ�e��Ǳ~yҡ�;��l
a_���݄ω�m�U2�9Q t[��>�0�����D�^���l��:, ��H ���a�����Lɩ�n�1���<�}N���Kp�K۟�:�Y�Y�� 3�M¨3��Η�\�Iq�=M�ﳏ��=ƩI�!S�&a(���I�X�N����S��x���dz�qs%5)�F�o��C���'��Py3�f�����p����FW���������,��J����?:ur��e��Mv�����-_3��J����	2����r�*��/��B=�L��S�W�ы-�b�R�4��!Bxp�:'�������Dqdn"�ND���)�^�&.��\k�z7@3�\.�\��N��v-�[����J���q�Z�2�\|K�a#���/sߢ1��.�s}&�:~��B�
w`vx+g<�f�����@.�^v�G��R�R��=w�&�Τ����B{\�B�<ũ�h�I�D��?+@+H��τ9�����4!,ͰR��M�gWg��[G}|>7-��D�wh�:�s��GG^��d��^��q��lu�7�z�}85]�+�%���.��>�62�!�M�=���ow	6]�* ������OR���/U���Ҽ�^=�����t���ꬶ0��o��ʵ��Ȥ�w���5����UL�_T�TZl==���r�4�e#ګ~9Eǵ����8`�����<eJ��Z�P���]H�1�;�f<An#��Q¡x����ǀ���V���-@j���U��hZ5&x$'/G�*���ʨ���L!)+!^ @X���E\s��vA���ꭋYu�~2��v���Ξ�Ȗ_��:\�3� �2�&s�H2J��1�0E1��x�)u�F�e��������3���P�s�Pao���X�v�n�<�Le��1w�� v�Zb���n?��A5��L��C�_/��d��V����u��UA~O�?�J�����F��2�[�)@k)�v�H�hi�?���#R��Sv�=��i�f�Z�����(&W����ޏ�G�#WmV&pԆ}���@�Dz]*�����.cx忚H�L1�.g�<]�&�{8���P�$%�|v�W(\�Wj=��1jp������X�r�ɧ>���	&^|!tm������@:#M���
w^��o��2�	��Rއ�1_��T��1s�x���4��*"�J��.&j�փ�PzZ����S4�Vv?��Ym� t����+[j��P����<���.W�C^�,�O�t%�U��SYǀ�B�ib��V��ydm�1M��vsB�u"yT��s�����I���\zA��b"�P�Cҵ�љ%�D�H��Oa�r!�v�Wi�Ū�gQ�*qv4E��u�菒��)�_?��T"/��[��?Ҥb�e���b�U��0w�S�)�Ȱ��;��S£U8�M�@T�fx�B���b��;<�|�b"G�7��������p�P�v�i��sb���@�^C���ƈ��~��<��P<�7�VVƌc����r>�C����	���y�ʒ{ۉ���Rӻ����6T~�	�Z�<]�x�g n��0��r�����Z��0�s��S������|����׫�3~J�n�!ζ�Ć}�)Ų�˪�������O]�ʠ�;HË�~{Z������|i�����ѝ��]U��[�L�0"�\?~7wK�	u�V����Z��P�y�V�H���|Mq �t��_��XH"!�q���%�~�t�Z�/�Y`U���� j�|�T�#�e,d=��2���T.`}��NT@Ƶ��)\��E_�Qz뾋��oP�̡���vc6��TJK��z1Q�=���t2���@vW!Z�TDV�j=2��L�����*6�.H�Rv�dg�I��͉{WlDRk�ơ=�o��t%Bg���>'�:|���TH	��D5�R�x�eɃ-�h��;'�����ATΜ�f��Կ�_r>��\�Q�j�ή7eU�/��J���q?��EsY���a�� M��7?���g �6s^2�����������\�更�j:jJ�X���,�p9�U�oǈm#Z�)DO���$SKv�p� �=�aL{w3̕r3�,���Q�Cw�k,�Fy(��",���s���@H�R��u��3���6"�?�����?x����9����#d�����9�npR,����4�"��g��qRU�9�ڱL��F�IQ��Y\桲'.G�F�~I0F�n�n�-p����h��K[��[d�U<If%,�&��o�����~DeX
�25���ш7����f����x����ۧ�������;݁ԁH�hx����� �ǈ�dz�A~���q��حqi�#��}s�gQ��)��������f>�4:�>��ޏ�m i��.ژD�P[<��wF�Ύ���m�`��多>8�p�"�V�|��@�����3�c�-��Q�����!ɿV�Ps���s�8?�����?�,�=ٰ�j*׷���Z���fW#AK��9�}������qb�U(~V÷T(��D�1��.쫥�D���ua��7�-���� �0��gS�%��Uk#�5���!D-}�y�zmj��M�=���[�&��)7Ѽ_��p\0�͘zj�&AQ؎}�s��R��f�)Q1�av�#�(_����f��$��Q�ǀ����l^�p˰��	>!�.s{-b,���dKF�;��c;4
eGkr	/�/�lz����&Z���hOn����� l$P�����>l��׌.UO�OQc:���x�jK���)�<��ӎ��A�C�O����eo���2���k�|:$���A�v2:��8�e�YY�Di���j�����U��!�Du�N��S�i�l-f�@�ܘ��zsq�)|j���	�ɝ�3�n����0x��dTzA*��ʄ/.OaF�`��:#2 �J�Q�����s2��5�S�
��dfs6�s�C1�A��հ�Mݖȗ4#t��ZZ-TM���F�9��MF&��(�A�mh	V��
L�C-?�BATP��114�{���P�|e;ڐhy�	$���,^�v���a���HTm�@w�~��73�_=J1�O�Jc
�p*�"Y�G^ Z��%�����f.rZ�Y<��M��ͪ�~�˙����:�e��W[� m�n����J�1�����x��'Z|�ﯩ-#�}^���e[���E��7��9I�����~��EqP��
��vz�{'�?�����lQr���Aʼ��ˊGy5��p\jnZ��V�w��"��[Pr�|ԙtXw�E~�Gc_g{k��]O����,k��*ج�H]��g	�!�I���p��°. �6��c��]�H��Sg�Z���M��`7�s�깺�����,Ԫq,�ɠ-��P)3�����9��&M>�1¸+Z�9��z�e@�xϽ^���yc���Ҏ�p�J?�B��4h�+��#�YV���+{:�D|�)�869���h�(<��Ņ�B����� �������A�߄$�1X��S�q�Ĝ����$��R�C8�8��oeGc��ǽ_���P������ٴ�ףLY���0��K��v��_��˅�dm����C�7m,a�o�o2�� ES�u��l����0[���#e�>mM���x{ͺ��T�t��lb0JȢ@r	
��V�O�-`�����\?��P1���s��Њ\2`UҼ�"~���f#���������[��8ƃv0���$|�T# n���7"�3S�OX
��������
Mݠ��'��Ob�P�����/���.��iu��7_*�p�\!�`σ�,6�_sk޳#���Q�EN���'���Y̝�>ؖ:���ֲ�k2�E��A���,���F~)[+D�D}�G�$�Չ�]nL�Hn�0��Q?0�����* ��w`��̎WscQ��b~9�p;���T2���Ս}&Y�8Ayq���$����Uc��y��U����#1��B5霕�Y��)V�D�Q���Y�R��SS�N�0[�
)�4��3�����Л��6��f���g��t����Ss��͝��k L�w��99�����cu��0����_)J�@՝Սn����-������q����%�k�"��5�J��xQ���4��η���h����H[u�HIe���)�$?�(���"��pFF���?�)O�a��vf�5� .���� �9D�׊�~�Ƥ������u���^k��?�\/���s������̔�NK���[ٌP�ix�S�J�i��#tZX��w8J���k��"�Z��\�=���R�g�P��6��h���M�5�3jm��� �����o�.�8�^%z};�'��y�H+F�w�]17��Q�RLKǴg��� ���{X��� ,EV������(��å�S�/3���T�*�fծ��Œp>hDW]҆�����U}�&	������D	�����

6|� ��/2�U*�W���o�3���fA���������A�d�aZj&����?�Wd�ęd`�K�U�cPJҰ�f�ޯ,��y囐C-Ѷ�R�o�tOF�i����M:�D
k�y���%�ߢ����	����Lj\�(G.~�a�4L�;LbOv�bM�Ѩ)�P��w�x?_b�5���9O���`
����*_;P�Xp�Y,.�w ьM���7�Z�B���* e|т͢��ӏ��δ�@�ʼ���D��uA�j�Oe��B+ˋgF�$-�ni"�G$'v�'y���$d�_��1��Bz8���Qʅ��N�N��ڑ[��qșe�G�3Zq[D�m}M��t���\�Pa3 �M�c�2�{,�KLgQ~�kܸ�t�o���TK�~��˝�j;������*���\�+�y�8�XVw��j�k%y����l�Z�JIؾ�D+�t4�9�/C���	W�x���X磾�W洍.&�fU{R�͓��*�~l�<C�u�4\-���`�������\.5Wт� ��<�U1fy�����3�������i݀�2�O\z5�����a�䳍H�r��͉Ӫ�1"�2�u�<�a���D�r��d�{	��%zq}+���)w5T���Δ��<��ٵD����� =��
�?��r���m�jIэ��e\u A�XU"/�Jg5/�i�ew�̑~#�W������
��dT��iqØ�MF�����T�(���!��Z-�wʢ3&���.�_E�7��{<T42��K�ȡ|���H�&��V	��`������b�..�~����p�j���?�ȼ!��6���X[�&c�#[�����k�!��#���醌VB�R�[��)���+t[\+����emFN�.4�<�U,;`*r��V=5����Xs@7I��9f�4k��M�r���ۄ�zu�卝q�u�i���b��i�������u��	BS&|ao�Q��:Ő<���5�Ѣ�f�M&*<������ �!V���~�p���A�?��5��ݢ|B��J���0Om�k��;'M�߶JV������A��"f@�#��s@0��U:��A64~Z�۵=v��S���Z�qq~�� }�~���0u��v�E>��ߢkyo���gJ�Kp8W��>Y����ںd���@�J��[�R:�QZ��y�-F�f�LX���6/��2#�H�/dX��K���z2�J����.�5��(��Q���r�J��8N��[뷻�"������ȥ�"�G�t1O�^��s�e6lA�S��y�%*�P.*�6����;8������gl ������ݨ�z���Ф����H`G��}c�Xȃ]�"�VklW��r�f���!|z��!U��#p��2V��w�1�@���_Bg�3(�d��v���RBt�w��=��I���5f�s:�zM/�ޠ��''�R��Ye�<tX�%��Pg}�e,luxo�GuZԟ
��DJ����L�bJq�C)�bΉ���p�����EI\�&��&;�ǿ4 �#��tb�Ss�lP�>l���`<��ywY|d96�|/~xֽ�ڊ�\2��%�*��赨R&�%��&/
�پ�D�!�x�l/��^�-�.4)V������#�NI��J�6F�q(���-ى8�)]�TG�.h�]�@"���n�<Q���
Qj����W�F��Ӹ��&S�l��T��V�B8����C뜻���!�T.E��J�S�X2���e�������.QO_D��Y��>�"���@i�2�@yN0߷�F���*c�8�֊��W�16��vx�p�F�k����=f�V/��������E���Q�-:��'9)=0dF�Gs4O4q&KU ���Z��W�Q�<�W���ۊ\h�B=�%��<�){�_3W箔�lԀ{j����"�A��O�۟	�@x�H�
�E�����~猍E�/��^Hjn��q����GfGE��W��'�����%��>�[�ی�'<z�g��	L_�`'e�������&O�p:�T-1�A�����F�^���� ���
�7��� �����g��B�E�v��lq��-��3�Q�ͽ�X���
������ut9SR�Ϊ$�N��T��}j��\ ���ͷE7����c�B�=�d�Sld�Y���U�����׿7�oj����������|E�:�ǝP%���������b���T%�a�����Z93��Zz�i�_(��ԅW��6�{rh��V��g�G�s:��`��_�D_oW�7=�݌UPC8K�n.�!b��~%�+-}g����Jk"�f�. ���$*I�C��ǻ��'U[&9IJ��〓��k1%NJ�c�P��r��bk�_y�69�W���m�[�V��`�@����A�̹�?ǃ')t$�.c�@�㊂����;�Nh�wt�^Xz���/���0yn�<f��� [��݋������]�Ϊ���/s��AqK�.�Q��K���8+l���ى"u��6r�0;É� L~G7�z�����c?�_�ܓO_���r�ICH�X��K��^�|5t����%����,�
�ą�{���.1��������޼²�>���LЦ4�X��l���ԁ^��O��,d$1�W�:?`�����ӂ���t�G�@��Ks'H�h��f�'��7��I���:��Û�)��Mi�	�gU2�g��t��E�A���(��x��3fo�@�R�cx�%���H/<(�>�%�S���PPih��x՜����i�&�d �Ks�T�ָi��\�t�%v3#�@�#�,tЋ��Q��K�RΎ4�6<���%���[�`�k~��-u��;d����X{Ś2��{v#�T�>�R��0��܁h,���O��a���Iȭ�`&ĵ;.ٙ�����.�
JK�F_���kʵ ;�j���{Td
��/�?Y��&�0v	�>���ٝ.���̃فtkdn�=K�ך����'F�d�A�r6��߹I'-@V4k�(���(��`�����N�?��m+���?7��I�n���@�o�J�W�N:a1Y�YGJ\[E��FV�=�P��~h[�X��!��
�>�i��6b�q�,�����&_��9����.jvqՑ����2U$����c!�º��ݏ���5�7~�.��u�F%���Z�;{u=l�8f�1���o�
؇YI�B�qI���g4�b<��~lߩS�aY
��R�i3�f�
<���i�:��E��܂�װ{ߴ��}��j�$���W��	������S�[m*�PHY2�!��j1ټO���͖-xI�5�g|�v:P=]}���q������Z��ĈKHQPQ�D׿��%n�f��Ǧg���B�p"j-��?;~�w����=#4�_"vem�yT�*-�,Y����V�t1��%������'K.��}��o��8f5�\M]�jϕ~��� ��\|w��%G6���I���fV~���42L�����d����P~�b�:�y��[�8t���:��-�Lp�nU��]�VT_ʌ�M�D�x���|�2�]�b�"Z��9gא�2���"O�8�I�e5 �&C�%r��N-W�rW(R�i8��Z~����'��Eig����p�#��_���+�W��/D8���f?�����."^�#08t��
]s<���~�y��� �+�V�$;�*CS���5�݅_ ��a�~������YD�S����ڡL2S�ʜ^/�P����B}�� rҡO�G�r���e�ܟ��+T� �i�:���mtI��u� �EkW��2�m��[��j�������b�ʔ  �vt��H����2��Y,���G}h�<Y<�(x-4��VR�Z&�h���E���+O���}��ڵQl�Z�� ᵤM�(h��,E���ెk�"|��Y̨g�'�gB���Z�wCL7������<����Ix����>ѤB�q���r���?��6�>�����N�0U_^�5j�E�@�x�K���96Ҳ�|W\^u���`xP��k�Ծ�_{�t�+�X-��H�w�~�`���+Q ���"s�3US����N-nE�7��k����6E�ɗ���?:NB����>�N���'���=�4�@ؾ�X��j5Yw(ʮ8u	Zw!�t(ZI��r/�`�Ùp|����ٛHH���˱��Q��?�_��C�盈�6;O|����#��bk�e�n�T�i���>�_�2�}��|�P�ե�s�7#�1r�8FC�xzcsu�|b��Uk=�w�8��$��;|�[<�j��JH�������F1w�2�ɴ�]��.�^���i��{�N�w�P�.��<HbK��N��'X�_4�'|�n��
���(󄥶q�e����hѶq���=.:�u>"���J�ʓ�UX�#\-��d��[7/��w�r:Ô���� �M�t ;�ꆸ�Gs��Q@N	]�#��t�S��!t@�N��C�H��a=�X��(��\�2-�Xםɋg�f�T�PX/7[gF��f8p_Zn2���_'L�'��և���<�9����)��V���؇�R�ܣ7}իJEӿ��T�i���I��A9�OO��_��Г��
n�o��L�BO�=Аw�UtDp\��^~�ݸĠ��X�h8j>Ig��{@d�"�+���~ɍh�A2�7�1Q8UK6pl���1T������_�����<�A_�:=*�����|�7��3����?<�z�:� �`�[I�� `wր� ?F�sT2�̋���:T>W�ϕ/��׌`�ƒ<~� 9EƏO���S��y#u�)��7f���7�����^k7ڳ��#Ϫ��_�u���+A���B�����Q�M�M@��!HI�!F�"���}Á*��]�6��m�,<.�9���xq*:�=�34�R�s%E��(�&�&�m9���F',��z"�8bU,�!2lI;��XF�U�M�z�@��Y��#��������>�*����J�Q�O�HnI٘��ǐu��g{l��n�N��V�3�Hx�P �W
I���-�Sr���	�O�\5�
^EC=?�Q��[���sC~�e}��]C?�gJwQbz���UW�G�O}&" ��Z��+��rɏ�A8Q{5*D�U9s�IϤ	�ٸ��x�����W�l���A�G��K'@F+C�jf%���9��S]-�p"@��/���Y�L�SI�z���̵K3�I��2mP��8r�����v�C�#R/�;�ew݃h��7��]�P�#左�J�j>1��<֖�6x*F[�:"������h�%k<_�|�]&��$5�=�Vw�IC�h+�AF����џ�yt����|���Gs'a��3,�y���_'-.G�ok�9���9*�T&���e����AH��>�p���"ߑN��uY��'�K�͇�6�6�)/\Y���D�-،Cf��Xê��b���*V^�h(kpũ�LW�z����S$�7h�&(�U�;�	G�M|��`�)v4��.V�{��4�8���O^5DZ���u��f���ީ���F�����'�gH�R6�t���\?](��1�	S�܎~=�A�}�TU��'�b���܄��:a`�Q�v�[�	ò�O�����R	揶����vC�<�1c�}^r�N�xL�V-#�V[8.pS���(W�Z:�����[!�����hj*���������^���jvҧ����\�n��a�מ�l�t�X�;iĔZi�ޡbۧ�I(�Z��b�>G�����;i�1���&8]�Ja���9
�m)���X���i<�&�g�����tb_�����9	/Y�0~���lu��2#�[������M	`:�\�������a=�ԇ�w�%p�l�+V{G��dP���6���>K�W�2�H\u�>
o����?�i	W��5�p<�1�������S�.�]��&�ٔ�{�b�Q�ZV�A�A�vn&uYEd AMi�3k�n$Y;��I9 6mۮ>n&3��|�e�JpY7I	���N�ZIt��3���?b])�h�kJ�p�q���^7<���	��T/=!]�t��8�)O8'�KEG��	ƃ�]�Q�9^�_���I(��g��1m�F����ES����l?r��o�P�S�z�oI��D3k�Q��P��_+"{=����>�٩�Wa���O
1���u[�w�˒_W�m���W������QD��Ҭ���>	�޸���{��,En{�'S�h��"�&����8���|�6���a�S,EK�ߝ��ph>0}Y�j�C�@�"�)��/�_��i0p�hK� ��%�]��+ֿ����n	<%�����&��<}���knE)�{���4��Y�7�Z� ǥ���顥��8K�ѥ!#�+o���?��v��}<�h��aO�dtK��7FX(n�~��1�kD�?r�kh��n��*��L�4)�ؔ��Uc�VPu��� (ZO�Mq9$&X��\��FZ�r��[8���4؃�C89>�b;4��������+	m]87���?��yY��ua�� �#6K�î���۞�{2�?���<��1)W:D�|�b
�/�!zJ�
��`*R�_�0�sd����#�R�� 
Q�7h��X�8���!�J��x��veho��1jr�Em�c�>L??X�����d�c~5�C+����UWUa#�d�ԏW�!5E�Ή�����,�s+�<�Ғ�X>�~H���S�DLi��ں5d�����T+��L����#D��'!������P����v{����w �|����=�"�~�E�=ig[AwXJ#���OBB"fr���R?�d-���P�_�^�>p8m`oi��y��O���6�iy��^0	���Г3@0F�NI��}�	ɷ�j�c��[��$�4��8����Mgd�8�ɜ�y��,�lh�<�h