��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY9?�C�><뮍�l
�j��+&G��)���ꋕ6Д��Jv�ܫ���qn{,=�A���sm��[����?=zC X��r,}����r ���b�p����^s�L����Y�8Ѕ��\##�A���T���B�A��45��S��Q�$i�od�w����Ӊ��V;mV���=��]��{��$���>1�y�A����|�����7�\x��؜���j
JsZ�]¾M*X���sz��o;���69� }��Mn\�O���a`�0�3�������*.7��&)쪓愦��2z���뺩/h�T�+4N�C2�#�f��s^[��P���fE���X:�t�����d^Ĥ�$�ޯ� M�C��,�*��ʏ��IAz��"A*�9��_��1�El�x��b�rY�����UD����x�U��&e�s��-4���a�v��{�#k^B��b�]�J���{k�#��6�f�o����}5����R~x�|�v�핳��W�ȏ��f���g��@XصN�M6� m�@�{k������B!�N�-84 �1?�`�ů
%��le$P�m���a��*��x8XM���9��HU��+��.
�܎�?I��gE}I�x	��O������V���Ȼ$���������9�892mI�FoY����S 8)a$������{����i��9��)���׳K\i���p��vԖ����3�2��C��NL$�H�J�a��� 萂�]X�.��$K�[�ɦ������Ń��n�8���J��I��I�D{.��*0�*�չ���x 3������C$�\�	��e����@<������,��);<�8�j6!߆�A���Ĥ@�Wֿޙ��~����H3E�{L�w��#�J��r��}�'�{��/~�|��{q�iU���KѰ�qۚd�}�`�m�����%�j)%XW�Z�Q!��o9�(�
�KesmZզ���}M"b�/^�T%��X!���:��&��x��%��Y(��dca�A��&����Ռ��+�����#wE���wi�@x��d�wa;�y ��$���2��C��D6�>���-�'`e�=�b�.`&Gވ��u�� v�X/8��ސ3�F����>��1�t[�.#�ct�ۼt��+^U�e�U����^s����5
L�)Z��ĺ.�OY�����F��Y�>��:�Ge,n{5㖹�p�>m�c�A[�t��Ήot��z�E6���RE�w5a�m݇�	hJ�K=��Y�$Oe4# h��4