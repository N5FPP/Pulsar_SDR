��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�۫k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��ע9�!�"��F�Wnb� �i��a��c��v�Ϗo@��Z2�[�Sh�+����,��ơ� ����ޞ|�e�JH��j�3]2�Q�H�a�:8r1��3RSK��i��ʀ��Z�� �@��2���
5J{[y��0�lg_�]rmWa�^��ͅ\���,������z�s�f���D(z�wut�pc��z��g!3�8Ɂ?�?�;�w����Uw����B�4L�˽ِ\��	�|!)4�{�u�W"=(
�lL�����*�<�U �a�����GY,g/��u�$+r,8.凐�/8�\8�}����>�+��L����5B���Yr��Ph��i�I4�__���y鮶u.biԴ���&��$�i- W�y���/C�L!l���&�����.��C:��{rˋ�5Wro؏���N�Q9�N�)�h�3�v"���94.t�}�ubyC��q*��H��&	��Wj���ͣ����[.�r�ה4Yd�1�|=�����l7�6�P�T���:�m����w��I���h��b�A4�=Pܑ�*��k�f�92"��7�6j9-4�Ӌʨ���ˏ_*�x֞J���6{�M��������k����_`Dfr���u��:{�s;ע�I�_�V8��D ��q��d�!Y�J6�]GwV9�%�I��^�|.�-k)!A��M�t����B�r��w��\��Q|��c��M�d�U :w8n�0�_\�yC(��j�^����LA/v�K	�ņ���蜖���B�41|�[���p���*�v!boꂽ9��	_m�^��2�#c#�-G"��i���]��D��w���8���+ߊ��3�+���=u�Y���fF�Y_>'��ӊ���e�L���j��{�pQ��4b��=+_?]�Ot{�8�Ub�r~ĳMK�eG�v�����o��h���J2���+oq�X�������؜�����܍0�T�?1��ߴ��5�p@����K�4��E�J��{I��͌e�&r<֓=�{�gW.G*f}?��m[����U杍̢�a8D����?��S�%��b�
=�P�H �IA.q���{�kDL~Lg���_g��ܧ�g`c�7hn�㨦�l�e��:�,�T��'((C�mDU�`90K� 7>�ׁ���T:���S2�n\DJ����|��8�&Hfd�wѝ�.B7L�_"%瓯�������>��&��<P�Hv4�s/��|��H���5'VH`x���^s���5Bw+#��M9X.�%*#!3�q��3�<&-��ƹغ7&�/�Ԅ���:�-���N}����Yzq�t�,P�lc	����ش�k����ۗxW5L� 3�ͫ���,����)��u�̥N�:O��Mս����0l�9f���е Ğ�T����٪�g@��./���x��,#h�'{Lv���\7�n�/�����)��T�D��X/�K�_9<��TT��d�~.I}�N&v(�9k;J�j1��s�+����
a�o�L�7���aO�S�-٬Mብ8�9c�Nx�Ν$��[jGF��\�O�}��˺@<�P�Yd#.B�?�"FGK����>J^m�ǖ^z7��"?�'@tmΡ6N3��[�2p9橝cPfR��	�l�p�R�L�ȝ��e��z0�M�֐\���$PDA����J�ӏt��q�ڎ؇s���BV��H��y��X�	gF+wh��U�'Ԯ׽,7����%�|~D�K��^�1-���y�`�>ښ;{f8��ǥ'q��Ξ5`���@!,�]e��\T.
Gۻ1���y7K�����ߵ�
�G����
I5m	gr�p�W��\OO$Ќ��< �H�l�1�����f��rl�6�w)���rT%�	����k�|*
���bL�� ���zPN#�2��g��,4��@���%����(��|��<\؆ �r8��!�J7%>�8U;�r�P���f2�d|#��s����'h�:�)�/
�es6K1�/0V����P�}��S`����n�KA�N%"���h�eCL�`\�v6,�æh&�a��J�c۰���,p���ԙ��Ez�!�~��o��03��qe���Y e����2�~���9�--/
�h�[�1܅��)���R�kd�v��`������M4����8II�]I?4o3�_%\����dպ�RȪc_�q<��G���\���~��t>o�W�9ς]���@��?��.V��� ���?��"=hXj(����:T��j�ϟ��'L"�t�A���W��,Я����n9s���@-ǢQ'E&��I&����P{��L,��Z�G-� j��f#$���Z4Q�\b�7�>����*Ttj��Dr�p��B�J��"n]V�NFMy S ��\���S�Pr��֗%�k6�7𣏕�#"�c��V�?�Y��k�jĺ�� nCG��9��_`:]7f��Ӽ.@��5�C�1�ҫ��S` @\(<�:�&�R%m�!NL=�`��7.l�<�k`�c�{9[�����l���T-�b�O��#5`���� o�4��}G�F�I$��e�ؾ�ҏ~�����]=��a!Vvk�g�V�-X�䛒�l ��H_�������z�?��0�,�iiS�j��n���*�A�9ek�XN�Q-��e������ӣi�{�iX8?y��Fc�{�1O�XW#�V|3�Stq�����
$��5�|.W٨鲍�-[�@X4H����F���
�x��^1��{�m$!��{1)Bl��=@�~�q���$�ۺ
kU!�UY�����_��6��O���^����E�u%��0=���~�%p�0@F�%&Ips����_.kξ���������s��JB *����]*������<�v8�J���@�r����-5�B ��
J��=���E6��)����A2g�H�9�u9��'p9=p�� �.��;ݭ���,O���f�y׾o��J�q�o=�=�����S���/�Y��0o���UG ��� ���Ԍ͞O��$��������� ��S������%�cޠ|�q3��c}I;N��m�)^,Ё_�ܗw:cFm6�������o6U���pL^�Z�2}; /�����S%����]ĉꆊɍp�V�����̘N,|�@Ql�!��!�b�Z�-)=��n�X�{ՏހWf���YE��Ĵ��$�k�\LT-���Nw���T��.��i[!����1�'�0���w�k��̭[G�`�W:�[,���i{S�L!!s�����M�����D,��K2E6E��*/��nk��;>�V�q��	��?�X�����v;�);�!�X%-�k�	 ��o��F�ػ���K4������h��uB�AMۋ��=eZc�e�ր�趦��9�d�\���q��>������̚
�WQ�u�8q��/F�UF��f~���x*��a)!�4~�l;�Oy3slk�Z�k��"�i�>7J�S��Տ*���;\�X·��u�[k �F�Bu.�@��B2~�k#O`��fye"�	B���Iペ��(��n`>pcL�}+<�~�sL�2���0}��u\����J\@"���W%}���2��Ն�Nh&��_�Y�o9��V�	R� ͊!;u0�F�y~�3e��"#��Pj����/o|��ͭ��8�B��u�+L1mձ�Ƚh���9_��+X[I��hlpoȯ�Yuoݹ*~4|�V�`��F�i¥�6��ʐlyGf�|X��n�>��F�N��?��/�X���ݝ�!��_@yx #r>�[0�]����;|՚:�ț+�"��/c�v�5>Ez�x�B"�3>�^߂�� �0�����ܝBi<1`��T���FJ�����*�w%�p��b�9U�s'�H^�ڇ�@K��=z���!{��W&,-��u�4_��
#���EO&����K�È^�i&���ܮ���4��o�k0MXpx��J
�k�M��#�f�$�Ky�Ƅ��t�Dg��TY�����,���5S �L��M��