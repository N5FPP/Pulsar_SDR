��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY�5����p}�"�,]��}���YS�6���h#��ɮ����z;U���gu&����Ȁu��D3Aix��`^Q	�$_���!y���ɟ�YyFCғ�e�ihm���<�,�����Zl�b��N{�M4fٱc���&������X>DJ�$��.II=�����-��J�{g�h	t ܥ���Z3i&�H*���.��K�<���g�̗P��RV��R�������w�g�*��=@��������<��EzQF7#|���A��#������YR���讑]���� W�/�R[�T�~��(�unߤ?�V�g��tL3#�{�����q�V8��[G�[��e,�.l�������������B���'9�U����đ�J�.�0���9̤g�k*��K1 �5꬏��1�=�^$bM��+{l���j|�<T�A��6M�f0�m4/�)=��Q���m��q_���:z��nD,�6�MJ-��@Ǚ���t���C�U��dZ�礋�妎+�@�EUE,�`���["��Jp�H�es���+�D�Ey /��_]譵`�W%�T���WG��2��#e-԰ p,��mȹj��g+�+��Y�SǑNF��1��H�TI4A�}�Y���`z�6׾���\�W�H|�]�R��V�|�'1���c+��+ n�F�;�=te�ĕ(d�/�B���i>�_K8NY��,�r"�󎨜dZOҾ�R
;��峗JӭX�Q:1@$_�q%������6�?V�Si�+ZQ����W�)��w�P�ݰ?�r/�^�[��^�����~Ի�<�/���
� ǿX	�+!��~h��0�4�t
�Ӄk("�;�U�=�Jow��Kc2郬�Jm-�&z�7R���^(aLu^�s����
ld�-��E�So_Ÿ~o3�uXǔ�������ٚ1����hOL`��O�y7��1$��4�f����M��'�MҼ�\B<���to�B���T,�yR��V���V	�	������J��i7N�=w����b�L�S�b�E#����3���T�z3�b���B��A�JRsq���6j?N��pgGm����zk�pf�<�9�����{�t�s����b���TĄ��a׽�:�<���+���O�$�>���U�m�=z�.��v�>̇�G������_�tU��<(���`8�����\�:u��\"��!s���Z�>��K�l��.�g��(v �V��i��%�zH.�&��<HSj�r��.lB��Qԫ0�����֨}hV�5S�jX^�"S�G�v�x:>���]��n10�DH���	^�P��VB<Y�����=�(�W���j�t-�#�L�=77�uGT����i5�r6Z�V�1����@j�#J����Smk֘�pPa�Mn��p���X��I�P4�=8H��&/��xT�5�����v����b�H
w����t.�����<��׷x�8��1��ۼg�Q��ġL4����>W���
�!J'd�3��w+z�B,[�i|ϑ֩'!�\�-�Z�l����c���1�ɍL3�=�-������Z�V�bTZ�N���OLpBn��$U���ө�twc$Vfg� c	�8-�z<���2?f�p2~�U���i�b}�ׅ6.����q2!*�o
Ӝ�`��6J��ے���3�4���(����τ]�*��l��#8oK#�U�|Y��m����l���G�����������Ӻu�ǒ�t�lhZ��N|������_���M���fL�Ge�1As�ɯG`j����I�5H��&��)�&��i+�PTͺ�hY��9����������\�A*��"r���/r�n��*Q��0~���è^�K�5=0ۄ�O9q�-$�6��}�$���.�6l�_�ZB�9Ί�w[p���w*�iP%��Wij��-j|{�Q��>#�z��7����m�E�e�#2f�a�fJ���l�P���5vFW;+	|g=�/k��&YM	zV���,�X����ϐè���4V��{�JP��h{U��ݜ%�x��3�s�C$b��)�2<7R&t􌆮<z�-��ݿ�q���3���eo��x�:s�.���cG5����,�!:2���Y�c���.k�<�P��R��H�֗��m�d�u{TS~�@�R �,�\�������h��

B�{R:]s(#��Q:Q��J��4��m����\E��O����=���|6��&��x�0�_*�z�����
́}�(y ��6"����[@oXM�9c�s�pk�-�|'R���������{��C�*O��1�o�7�h�^ajq�ߦN�R5J-����K�/%���-�����s�V��Q�E7Ǥ�Ǖ��~�������O2oNֲ2�m.E�W�a���:4c����
R��BKO���|{�R���S�)�g[���Dk(��ƈ�u�`SDloC?b��?���+�I��2�T�-�-���'�#6��h���]ַykrܿ`1���d)]���C�1��)��y{%��D)2�B����Ha�ĽV� �l�y^t|��l8�� }d����ץk���qKPE{B�Ǒ��@Ff���RQ����w��/�9ほc��
�uq���{"���b�I]�1o��%���X���LC��7��x�t駋T�= yp$)uy*�MPM-�g�!��Фh�m̂PӱCz�P����S���&�ǈ	���Im�˳Wh׵�ѕ{��bpq~���8
c�cqm-�oB���Q�'��a�H�H�Ln/�B�
A �G��41�y�:� �g�A;Lj�p��`,e�9��#������RS��A�(������ANE�b��|(+E7�M��n�6 ?]����X��9-��.?̉��Wa%�Ke��3�:.��r�F����F�sJ�8�V�	:���z� 曭9��`[��{.�R�))޺��{�J&�݃�OD����>`/
�tlq:'�X�	fR�`�W�gG߶��	���ǎĸʀ���i�MQ頼��C��~�+Ws��*�w�%�����+�E� �L���f��I�۫�19oV�C�ߍO��_
!�m(�"�\�۲P�E��}MD[1�k�t���տ�4,�v�5�sM0�zpk7��
NQ@#\]�)�^(@K�Bl��{��Ril\���vY��5h�n���'�޻sGOh��(Å+bL��@C+��ѯ|���8�ho䝓E�x���l`+�9���|�2%֤)�dF
f���i%��	2�ʥ�:�hX3�I�Z��Wz�R#�1��+���ϵP���쁣O3�@�B�ć�F)�=�kDv��A�(�<{���6k���m:*x���7c����˲f��ڗ7��!@=E__������5���>� ң�m��tT)���l�>�Ce�(��+�r�`���.�G�TH�Y@�����Ժ�a��Ջ����#D�Ժұ�)�uO���@Ô��,�C|�r�
%�c�B]�l��g��o�0`q�[�`�W��Ŋ�@=e�$���$6�Tcv��F��}��;�8���S�;��ϐͻ�ŵX�1߽;`������� N�N���0V���;�r_�5sv<u��r]X�� 6?wۗ�LL㜨�+\7�5fv��~jCP$��A)�2���'82Ԝ V2�3�V����r�%/�f'��w�I.�۸PQ	5�
�����赼�}�Z���B��Y��9mB���O�f��% wd��j���\, Dw�*��dt��$�T6�/�d2L��?y\�F��.j��_�F<
������"���<�+Z��B����(@R�}�a�o�2=�=�	�:����3��f&z{�o��c�&&6v��+�E���m�Y��0ɼ�+$rU��<c|V��Sl^�+���^.�/@��P[��hg»,*�}5s�3�q���=���J�6��"�v��Ej�4@���Q���Ń/��X\0"��$�X�& ���,Oj��SR�@��o�e�*�Z�B�݀�۽� mZ�>IT���W��y����@p�'�����4�#$�7�X�Sܢ�r0�Ea�!;�0Nڿ�&
�z9�Jp2Uu��y
�'�2���q��@���J�;&�vzY�4��6G`Ob[�+ɢ��w���O�����|��]��0okG]�����*dw��)|�5wr���o��- ��(f�?Ji����޺�[`��59ɦi���W�������fנ�5��ɨ�p-�����N�Z�=�
dD@e�;����`9��ش���Q"��_᷌��a�u��S��8S*��U2�%�Sb( r�G�S�)�����N�jy������dV��\\-��JR&ʀ(��������a���N} �T�/���[����PÞe
iuݯ`��sc�٧1���Uϳ�����@	�
hث�`��+
�`l=J�q��FE�����;�C�5@�M�4;2�bE0Uϻ׀��^���;O���&����܍J�P/g�"�5"(�<����߆G\�m>��!l��I��<�����q����v�W]�	@��Cnx�N�n�����D�l�a�9�)�<r��ׁ+����������L�;���>�0��������ԏ���ˮf��	.��j����G�!����W�z9ZZLlj�#0̴�X��.U���~g��6��Q��i