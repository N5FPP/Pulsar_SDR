��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY����B|uz_���	SD�2SY�mv�7*	.;*���hR}Ğ:�	���ˠTK�zv���Oy*b���cbE�����F�~���NX҈�
N\�@����a���ȷ�P��XĂľ�����myҾ�TA�mΔ?E7�ɳ�0����s�����8f�n�h	�x�[v����@�6��d!�Ɣ'6���W�#��F�g�}5G�/<H�'v��i)�Bƥ��ⵝ����!��!�W�K�·x�M�z��.�}�6�`�#�+�hL�s9(��"�k�@Џ�x��U�_=1E��l���iʕ������d��,�߳���2�/��x>N�go���wZ��p����5��l�>k����I�i�X3��AQ�}�nz7��ByF\�2�hr�*�ڢ$� -�L�Qu;$ǋ�B�M_cC	m0����e,g"/�ǚU{;KTh�a�6	"��ĩ�����O)�B_�p{���c��M����sK��@�Ł�~������S�9Ɯ�K�|�g�yXֽ��dld�����y(��~J�)�� L���b�t3���˱2�|�`��T�P�J=I,9$�3�HmAn���~����~��
�蕗�������5߈����1ܨA�a���I<�D*�`��XS�R�p�u63G���zrQ#� R{�t�C2��ϳ�ꍺ;-���4��m^�/q
�Ď�P�w��r��;r�%���?7e�hP�y�����:�%�y�u�_�^�U	U�0�W�լ��߾��'vS]>լ%�8�� ~�p�*+3�{Gj��qe��|F�u4�a�,��#�Qyn��gZRb�ڄ���b64��[˷b6arNj/��
')�v���5�Z���9X��Ѣ��U�OO<�AƮV��Ñi�H��f2����+- ZN�_�;b>�i%}�H���V��I#��Y@����z@����Q�꣉��#�꿨B��DE;�^�6n��S���VEɃ��e>%�ߧ3�:!z�ȗ��(8j��)�q��@z�?S��pQ�2��� �����w#�:"Wg���6�Ƚꕳܭc�&6��Y�����UPҨT׳����q6@��翏��/��/Xy�l����V5Ѿ-x�v�[`����\�p�o�l;��m��\����.�܅K)Z�O8 �z��,��bb�3�	�Ч(�p=r�6�v�j�ſ��[Jk"\�g��x}rd�8������־+�����0b?>w$f�����cl�J���+<����+��l4M�X%d�ӝ܏aݴ��-�s�O{w�0�m�*M��g{.{�`���K9)/A�� ��P"����c���y�Ƈ~��D;���Q43�Eg�tn��X}��uG������4q=�����YWly~��W���P�w\�m�hJ�lzd��b��s�v#pL�~�_�p�`��`j�NR�i	 ��r�^̄�O�P�1�F!����u�� k���I��sk��5�׷y� ��ҋ���Ѝ��ьLCN�DzStet5�B(�}����8�P��#COq�+g�Q-�a�yDi5l��X��^%�B��(1/^I|86�N�>�bq��5��[�KHK�-���
�F�1���*�NaCQ�����2�Q�H7����¬;��=RHO�� �i��~�����ɵ��.H1j��0L毋���)w|��v��c[�����/p��U�m,�m$��Ksu8P���Bft�1�����&#�8�o�s�˕$�{�ݽ�3$$X#���B�IZ�?{��*��8�����O��欏CނXUu;x����Ġ��c�5P)`�ԡ�WP6� uF�K:p:��#/�:Y�/�#��A�W��m�,S~�X��E0��4�ZOd1�{��iԶҀ��ft9����ߑ�l�u��K?}_�`P�Id�P��<>Hs��ϝ]�]��PɚG��}�àc�-ގT�8D�� �0N����а���C5���#�c� �%�¶�5yX�3�Ti�,��e<+��,7���]7�z���v�uع��=Kk�O�f8mk}�W�y���̂-����%��94qbѡ}��O�K:�s�C�b0FId&ck��0o�jq �J5����GZ6p"��v77�5P���ᦩSb^c�`-���n;%�G�g��!��e��+I�~Y_Z����)��D�VAR���9!�R�b����Jd�k�,���1&��Q��gD�H+����*HbD6N��V�O�?^f��Ftmp�y�K�����5��z➙3���Ҷ�a:��Z�}��EO�	w���oo�t�E�F3Yr��On}��<�#3�)���D���-{����e �c��L��>�|��'rU�!N&�׏�b�J5��&�_��jKa��Z��zd儇��(���4.0$ѝ���������P�ziUi������3ݫv��з^�98���"�o^Wd�	cmOǦ�_�F�r�9��PKb��W��ip�<y�7s��CD�?��|�:bԫ�;b;�h���&����=@̘�=�o�U�2zn}/�,[6����J���/]�?�?���[e�$ƹ�(S�������@l���ۦS�(�t^�ij��\���������zX��I����V�����*�����ߝ^�4�C�:���P}ԲTdB�	�QpE�ۥ5� �^�!8�T#��@�Բ.f�(W��G�ry�R<MV�0N2j��:�ngA�9��7��~'?G��!��[ 0W߁���˻y,�S����A=�//��]`�?nu��1!![�O�n9�K�&�8X� ���
��^�������Le��-
 ��{q��P�7$�`%��H�M������~6�}UO�����h�ܜ�s,��f�*���W�yH�@���6:C�BP礏��c�h���OAD�/���D�ę3�U@uPv����5����f.5w��d�L͕�ʏ�[��!��~� �n,KR]���HIQ�^Ф�0�Ԧ��z�&�w�~��2i��I6epT�F�J2�h�Tܯ�n����"�	�^�x2�J/ϟ�А)��7\�S������W��9 V�yȼ�� *~)���}��z��<#'_����(\���ZX��ĳ�AY���2�Ok�l_�h�WR�p �	y�ᢇ��ԉ[��A����|�:�=��s�������Rh^�)`E_۷�`�6�塚��:�"l[�j�d�_��Ɣ�pB(�~�eӬN���J�{�C7K�G@4/�������5�����Us���K�"U�B�\]��|f�`iU9DЯuJL��8�Z7z�J�v�'�~�o�O�[X� �b$�H�������Z������#���?�TC{�O6��G�Mq	�N�#�W�=`m��H��י�����T�κ� b�K3`��ͣ��D�ڗ�,f1��f˛��Q���Fa���LP�i���p�����b?�NM�L�ӺuY������v��v�Mo�4�>%&�t%��s��z%�[�䦦�Y�8q
�H����䐴A����S��ʑ����e�ʠV,�i�jm�N����+d���;K<8w�� �v��#8�.��2�s�?bT�E4k_kc�����>-�a�=�_`*"��x�nJ5R8��A��QZ�D�V'ʴF��{PY�^~���W	^���A=�r����P�G8<�~�����<�X��[Ҕ��`l5���ˣ���j���bTl*8g7jS����l�&#���G�o<�@*���A# �����G{�0�:}Z��g�y�K�=�"ڥ�^9F�g��"ö�����X�3Z�It�3����vj�"6�2�	<E,� o�Iw�7�#Sm��/'�k
[�=��%*��W���(����G. TL�/j�-��8ؼ��%�1�B1J���\�Ɔ>����d��h�l��C)�J�+.����!e�ZkJVAG������Ă';��h��iR��pVtE��������9���1-��b��������,X�QCo��e��-�<��# cG�0������f*B�[�u~���:gD�r#��K�.<�w�ϳ���UMX �VK�+�L<B�h�a�����?}q��(�fb�v�3�N�<?gc�p�?�����,�qE޺�����G8�%�R];AO��U��]:�r��]o0�����"M%��nŨH	4���GwP3\:eIB�mJ���M��Q��Xs�%;��Rq!˙��^�ϣ���\�DZc�t���m�X��s1Z@�.���L�;(����w��"U,�q(������Ɲ�U�ռ#��k�i�ϥ2�j�F����%n]U��E*�����ɡ�I˔;JP�������~��!���I2|�]O�Zҳ�;��������L��*Zl���j�:��u�V:�G�52U��P�����#��7���'�.iJRK�����1����^<`MCiM|up�1)(�?�їb����NjPn���hB���00�m�c�e�F"�����9�)_Srk��w�9��4"�@$b��F`	�򃇈���V�KڞB���Y0��{Z,�c&b�7ɴ���	�)_�qk@���û�s9��<�j�V-w��	����P�����<b��,y