��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�۫k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��5K�z��!��[��S}Σ{$Gx^����c��ƀPfƆ���|mU��_yr�m���#����}upb�ٻ�-�O��z��¼��%��c�@��p�2O�*6�1#�+^���>�
9���Dm���w7��P�^�1`KH�Z���&���8>b� �9�&�� �z���޿J�5�vѧޤ�b��e�>A���{p�D,��mEe����@04�k���J�� �,Y�n�p���㩛۱�d�#�A��:�?��xk�.P�13�o���Ǫ�CM��K�K)2��e�Q++�Y���;ܣ �^�I����V>hx�**.��SS�y�,0�QY���Z���� �H��S@$�y˷z���C&1P�g>o����0�L�e�#���Lм��m�z��w��}���a�mX�g'��JuUʲ|�Q�-p5$����"BS�<M����ez;�X���o|0�v%|��(�d�����y������'��kB��� ���h��s��l�&�,��љ���4�`a}�g��0�K�[��y�v3϶����qw�3Cw���7�ҕ�����Y$X������瘗" �>9^`�΍�4mܘqG�����}�\^!U��2���&�*�9���Fb��у��H�7������w�w�}`dd�����h{���"���ܭ~��*����}�N���殺8ڪ��a�9�HS��'�#l(v�����kP��˗HqZ�8�c����n�qf{
��ri����6������}�x�P�<=��{N�4�_rN>h��~.(�!�u�+qeߑ��Oڲ�aE�É��2o�X/$5��s�E�mL�:I���м1Ȅ���3�,��4v�yQCzD��쁧q���q��y��􈸄�CB3_X~)|�h�*�\�������L�T0~eY��hD�]p���t�Z�����0��t�'H)��rO�F���w��_�]g݀O������3O�6�0���@�)�`�bg<$���"�Ϲ��Ơ%l���9Fi:&�7��GY�5:6�I����D}؃>[�%q�����K�����x��M��e��c����eY����%-Q�x-��f����z�1�)��7K�.J���tJ���w�������@޹<Q�$U�Ab�ͨ��߄!9���͹�,�[k�X �c�W�A~*Um&�Ғ���鴉"v����O2�6�Ɓ�	��L����Gtj'��P袔�'�G2/yD^�|%�_;B_k��1��pԼ��O�"
w��"�Y�3JtS�t����m7ȇR�\fZ]p�;��{��mb ��]������r�5*Hr����hy�,�^;HՑ��!���.w;O��7��gz�E��_�(�*T ��wbKWFC���qy�`��/Ew��1]����+b���U�F��5W}�5�Wv����6�{�U���J�ؑ���ӷ�`�_��r/�Nߒd��3i]|o���Ɂ�\B�Y,���÷{��F6W�M*��2v|&Uʱz�y�-w��8Pbt�eIe�D/�b2f�nm���e�S�p�rMC��N������&��m��n�U%�d��b���'�@������~1,SNB��ĩ�` ��\y$�V�~��l�05��)}@���	<�-1��]k
Ω1�u�|m��u�� ��E@^&���ُ�J�a�X�(�1/͖�(�But����Q4�Z��)��X��֊����}�գ�Zt�[$3b,��c�4ɭ�߂W62� s�*��)��  �t�*d�u�@���&�Y]Z�
H�H��{;��B.�T�Cc�!>X�I�e��m��n��!j]�rPq��x���tE�0�u��K���t3���J�U5����K�:����p�l���U|����M�E�����b���=*�������z���7N���=��1�d�l��,8T�"���zb�֭N`��D��~颬7���Z\2�_x��4U'�O�<*0t,�WpU>r�#J?��"Ԫ6� +Sy���2ա�����r�(=�VjN��� �_6�9�>4�W�>�Gj��w����G<>cl"�2������VJ��4~�����l������]ύO�*�9�%h��7��+�Qr��e}Ʋϫ�~"�!W-m�g�EP2u�[����=�r%�O�K� �on�`Fԋ���*(�F�6a��)u� ��fכ���.�����*JB3�ö}���^,z��w��%�����L�%kA;���z-IJ,.�k &­����@�M�����9"z��q�)D,i5s�'��e)DG��Hmv�b�sJ���B�i#u`���͢����C�BT�t����b�b�$h�/�Ubw�� �+���	�U���Ƴ�F���A�Y�Ϫ�Ч�q
����
3����vNAj��{~J9ڥz^�����"���em!��Eu�y
$�"�7�쫥��9��!:S��?�w���.���O���63���]��)ѓ���$l�E����5��G�vi=5�!�7zAj<��~�a��}�Q�cSVO����j^��^�r?���r\�����h�6���.���i�R�I��<8�H1;��=�	�6v�;��d�jvc���#�y'J<��	�*��F�f8k��q�y��i�N�b�*��c�!�]^
Դ��_%�s��`����iE�۰��n����:o��x7��\��0wO<
�K��?Tj`����jgGqi»O���n��[2�#f10�hu�m���	�]�9��u��y��Ѫ��^�a�ƴ�p_�ٙ���*��sxXG?A��o�33���L=�1��E#�����(,1r�qG����P