��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���2�U�z�[B`�#�� 3�����E��R�=R��1��TH�G��N�����` �۠���<q��c}�޼Y%�(�"�sڙ�AӛXG�{|��AT��x�PL(�]������r�@�h=n�O�^����	�{K�*�q�a�T�FV���:`��Q�օ�H�m�Z<A�=p�/R�ؙ��a8E?	[��C��|_EM!���MP��� �R.Cw�j-1�,?���Mׄ��E��T��� IZ$\��h��I�d���cL�mG }������3���@T�G*C��'���"t�a�3kM�����p�s��7�Q�0�[0�yS-*e��۞�`4�,u H��{�k�p	O-O���I\��vC&�] �oV�T"f��.�=�-ԙ�v��vd��__)��#� !�zL^�Z{������ۍn7�y%��O� ���?jr��+i/�Ϸ�:���H|^?����]
��ѩiYm�y^�%�rZ�jJi��d]ɞ��al�L{����٫��V�L�c�g���|�m�7Wbͯ;��o���X�$j�O%����5��4������X�N�����w}~�-�P���^_�w���a�H��&-�_�}�(Ji9������U�c`;s5�2R��p�l��d��<��z�2P�\�0�C&�DZӲ���f���+�^l΂R�o�*m��b�px}N�|8�6�Hy���U��S�=W8���5@�?���gt!"E8�.{֤�8��R�᝜F���������l�|+,�?��tD���DY%�mx_�����-�_�Տ�^�W�$f`a~'�
w۪�2]v0'�Q���r]e�?�#��&�,.�`�R!a�F��)��x�ӱ���sq�}��yM���$UK,H�j^�E �F����`�%����z�n�8&��w6[ǂic��
F;�v��KL��sCˁ�>Bċ���o�fwLu'��v�n��tꁡ�"W;�K���z�W������1�:�1&g�E�G^�	_J���U��y����zE7L��s��I��yi�����E{��KbK�50��E8Ɨ����v��I�Ͳ[tF{T�G����lvb]��Ң�Pn�D.�3�V��FV<u�e�����	������ӞD�Υ�g�cPjJ�.�Dk���y�N�	���Db!��F�Sa�@�Q��)�H�r��@������`������b���nh��l�
KK�K@`{������@��̱��rU���������,��G?�z��-�Z3���Ɨ�V�A�.oߙ3I�η�쑌�����|��P��WbB���%��:�S�h���kR!H�_��W�ti=Nz̼���Έn��;�n_�u�t�sV�h��(�I��MJR�B��o*��qeLs2�2�@5�B@dB���Q�`�Px��:�p-qF5��.}�g>M�ln5~�t1f~��&K�k�Itv�<G��8�L�m�"�~��0T�Î#���.�NQ�9p4S@�7JTF�F�?
���c�?��*��q,S�C��x<D�s� L��2�PM��a�l�g��!K�Af�^tl�))��A�Ȏ��_$E�����2�i�lk1����@�3rt�v	8�R����vi�G}#=ց!��r���K�@�-g4t�	)Ou�&�����
�$��Bȹξ�A)T�	NJ�xo1�)+�a�������ַ�s_�9��	��J�B���ƌ>�dߥ\��|,�H?d���!�G�hIY��� �\c����F�ԛ�w\�ť7�ܔҁ�Q#m�@;�*�W�_K�m�{�̓�N��ڀK�G�ʹ�)��&��Cxr�]eh�mpƢI��G�N&��ӉR�d3r��$T؛�ң�T�bh��DsN�����(Ov���$�.MU8I׭�D��d1"n�{�]ö�ƈ1�O�y
����>�Q���By�V��5 _�|f	�l�
��Ӫ�]Tgi~�T��Ԕ:�]h�'GMnsK��(d���H��z}~�T��VR<�Y=��ODZ;$�~L(�_ơB.i�8�*�}e0�Rt1�J~��
������"`�[Fb�<܍�x� �� �%��Ե׭<��Ua�tO#ǋg�{�	�+j�g`�e#{�̏���'ݗ�>
!{���R���ޤ�䛈��	�� &�Oz�h�}��	��+c2�Ř�e� m?���CÅ���d�ۊG/�!_l�?i�dl��C,���tj���Y}�v�m�AJ�����<T�w�gG�c�ɏ'$w���o�&��.B�B\s(�?i;XzOLiB+�cT����z��)�%�"s�f.�Џ�ﺝ2Q؍�/ɔ������l{���67)�k��'�F�����i�jq[ٻ�pq�O�[��6���S��ʏ��S4D����o�h�RxP�؆�(%��I�+��;�zU��&V7uI�]i�4?����Q�> �=���U��֢l�"ǰ ��,�{�vV?u�h�Q����i�����x"�5�ek&��QQ��`}���8�-�Y2�����"JEjړ���0�㟊8�I�y�j�H�j�������{��)����T�)��*M��>"��Z���ܦL��U��8�k#{�%/��}�F�8�K��\��] q��ѳܪoB����ɦ��\��\	��h�!,�^�$>٩ ��u���zl�M��}�A�^��������/V�ͺ�|�f����՘>�7����k}h= m���6O���3����d�u�����.M�^���׸����PK7G���>�Ef������}O�E���9��B��8aMJ�&��o�Ȝa�6������s��VA��nT�\�������7��&�TWR�&S�����'Ͱ�UBm�B(�<qm�]����"�V�%U��=�/Jm�!�z��֯��^�d�11������J��( �n!H4Ló���j�M �w�<8�� �6u�Zv����i�V����	@��&�ޘ�T����r\�'�(�Qq[Z�=�5.K݅�nw�d���dF�7����^��J��;�ۄ��^1�&Vz��K��NI� /hg��-���*�zE�J���T�-U��V"=���)���!�ZuY�9�Ɯ�=��.T$&M)�i���]�	[�æ\2{�	����L��=
8w	��x��}�`����9۟�Y��8�ďHc%�2�禶����1!���h�RC���wj�&u�����s��W�H��!I�jB���P�7��S��e	m0��
�'����A�S��կ�5��4A}��ZJ��ٜ&�X���]�>�N�J�\Y��u���6��{}N���-�Cj˫�Z���t�����H�x�^�D=_1�r5��	�F�]��Nl�>�U鴭z����C��(�\��Ñ����汏�5Ai���]Y�D�,�4�ǾF]C�<��� ����#B�:�'0"�j!6G�1��M���l�}ܟ��M|��0&/��=���Ro�e�x���9��No�����(6�0$5Ǿ��c��#�U�s����G�'��}��I|�~J,k� �!�Bb���|;�4H�t��gC�>���}i��-�E-l�g�l(�ԓh��c�+%�Q�x��YG�}�}�� "ʞRk !K��9~f�Ō{iv�)_W	Pk U#[	��_)�N>G����<:��׺��]:�g�ya��$��oޤ��u�m�eY����t�u�N�9�lK�ʩ�Ci�a��d��x(�E���2嶳;q�!�I�1�W�nG�zĆ�U��Ĥy�S�-�3�b�D���W�3\��DY.6���N��͓=�M�G���M?Vj�Hj�=ו�L�ʚ�BEOH�cE�����:g� s8�P�K���q��3� S#A��5�`�F�O,�4RQ.H�ܟ��=�4�EАú��˵.�TQ�րPnJ��{�!�.P�{�E�)����l�x�,��7�����:�RL�\I��;5 �%9g`�W7 -��O�����b�R�A6��rɔ5K�z��ҹ��EYߑ�P�z4tT1uLW J���(���_D>�m|�݃}�1�L)�]�kd+[�9|�*��L�i5f���{m8�(�Ŕܝ��%F �uP�w�A�'��+��=��1"fc�5%��u�����<a��_�6zU`�\������i�Z1����dk�w�\�N�n�f��` �lt�K�|��Ab�p�!b�q��)��!�e]9z���o?��j��_�v_�!�N��Y�Q�t�Vg"8o{�~a���	��({���ǩ𨾪p�q�V��>���7ś�̽1�K�&[f.V�8S#�y�&�)v% �H��k�e{���ɷ9>��!Î�GD��u����4��:��I���8���>��br�z�� 
�½��Z�gaݺ���]�TPd�b���fKK�:��� a����]Vr�!�.C*�P<_��ƭ�H��o���C����Pw~�"�y�a֯݄z�����VP;�`�M��������ДA�"�H�[��ҽ���4��ЄrAl[W�F��a��-�u��3"
T<]]�]���SJ�I��*<��O�
A>h��~��BOP�N ��6?�bdG�w���2��|�G*�.\�y�&�+��d{^F?0��8�Q������jI/r6~vd#�j��I�z�-��t�1v�7Z�1����o�
���6��O+� �=�!�r®{����o��Y* �	?o�rUk���V3�j�&����!���S22O)H���Њ�J_G�^��h��Q�;[]�R�c���%�'���$�����0�Pe2[|�M	�o�+�
�����fIT�U��Ӣ������^���I"����4:Ƹh��^�`�����=�]��I�cC�-I��3��ɢ@k`������"�C3�&��gkR|��挎ؘ}������4���)�v�.���((}T�;�c c�5t���(Ƭ��~�3tL�1S��Q|��趪y�$v�(������c(��4������|2��t/�𒈹F1��f���������ʰ$��_.��cI�DBJ�!�$>�:��l�C0t<��
1%��8!@Ť"��C�fW#������~r�md��nPhi��0�).�r&�뢯R��z_��;��'D�m8ҵ	W�5ڳ���ա
Q�)]���f���Z�x&�cP��L������FB���UV�r�WTKm>d �J��0Bwu�5���I��_V�{�qs, .�R�"_ԣ�I?­4=G&�e�䭩P����j�[B̀�4�D��X������Y��X�A1��?��:���4���mU^��TS�|��z����V(A���9Kb��e�$���f����W��4�ʩ�^C3B4�i[��L<,�ﱸ�H��bOUa����@�Tap�d2�ꥸ���?i���]։oIӜi�j���0Ė�&G
���u��	��\��;�o\���	�7��aR�K�L�M�`#Jp@M��ǉ�����w�㌈P%v0��)�_�ů�%�=[܍�}��x�{֊�������ܷ���`~���/�Ɨ�&D�1�xmٴ���pv�I�Ż`����7U�5B��J�&��t�2r'�b�r�j7�l�jxX�f^�������:��D:*�Ľ����`���/��?|��W_���!�g~Ba� ���/�ȮI��^�&Ѿ=���(:u�V��r�.���:��Ƈ$��2�P��5��҉�o�?_�RRI���PY�]W�'�� ���-`�M©"ؼ:����1m�vN��Wg:��q�&1ܳ���:�6������`��͆N��Z���O�4�2����pS���0��M��4�z��.`����3�}@�K�5�J�|4�_;�פ�	�S{���ck+�D�8� ��C��(�y�	�j�lƨ]!���%��A"�����:|h4��cf�/���<�֫f����V����b����h�Υ�E�i84q��Idph��L]+��I}%B7��l mB:���/)��A���Ys�8�ak=}��v?�c�"��0H`���������ra�	���ES�sD�&G�cQ0P��	��[�����Sr�By_�\�6�Ӱ��ЫG���eeH<�W[y��^�
��{W[M��\K�	r�bB���]Wั������˲:T�}�n�]���^x1e��r��|6��y���X~�P!�'�o�
��ۢ�{�$E�yq��+�Bqx[j�Zߑ�^�cy�LUX�f+�x�~�f��f���]|\_"slA�`�Y�Us��}��,�`�g+D�t%�F��2��Q�k	h�B��t^��r��a�WO�13�o_ѪY���vؐ+��������%>�4]��KޗSX��͎�p����=*f8	Btv�9����y���+���~l�uK.|�E���.��9LEx��)��F5�h-%Y�T$x�jnz�@��9���׭}�����K�ۏ:��5 Q��3���ۭ,P�[w&(Z]���<u S��/��H�2� rd����;�T�{�n3��y� ؊n,_(���c)1N7(��\�3}��zVA��8^w�U�\���m,W�"�pD0h6O*�R�fT�SY��7��;CY3]�y	��8� �E�$��$�Uî�`�h�=8T�� ��y/�o������ABMn�&�z�Y�b����@��K7OG���܎a��i����4�b뻊R�\���l�m����~rB,z����g���Di>�*_*8NP������G+cF��-J1�%.	ש0ȹ}˜VÔ} �e�Zo%B�����4�)��yA�<<E�Ьk���a�7����"ک�&.G䦐~ݱ���"{�[:����9,��_ϐ�2L[�p�WL���P:^���1T�\��N���+=B0U�̪Yu=sBI͠��V�f���������w9�)X�.�sA	a���<N�|���3)<3�<j���v�/����_��~`h����	�Am�"�4b\;x$�J��q+.�h��_bگ?��j�դv��U�cK^�)��y��9��ga]PImH(>��0W�댘;�����$u��@?�k�]�%���E���xلt�z�4��Sd7+��speě�8㊶�("�k�7���ۋ����f�*���
��~{�L]���4f'	��Z������4i����Y*j���Q@�u��n5�k fy�K�ϑ�ځ�Y2y �:Np�����a�5�#�,����&�h0;óǥ��%҄��^>�|U�������ѵ�U���ӊD�����%���l�ӗ����:\���?�b`���g�F>�����m��[��_��TL��
��g��Ɋ[�����&�R�3Kc<Ӱhh�2�K����@zdX�u��t�>�	h�K�"����h}>�ˏ�0�M��`o�8�V2�\8w�Qo O�M�p^)�������n!����E�W�����,�I���9�!���i�^���t��&k����Z�zю>�
%��®+�h�\�S"$Q0���Zs柱8�n���w֨�݀���Ea,���I��J��Cc[9h�iۭC��1�B��.��Ns���W�N~#_g�66�{�H=yR�T�W!��e7En�9{��k{Q5OR@ݾrX��j7r
�aK��	F��,v�E�`c�\�Bc νu�9G!i�A��a9c�5E��HB@3r���e:2a�BZ,uҒ��ʥ�>�
�J���q���U�P9�xX�L����Q�.p���D�;[\澃��8N��`�a������U.�����+ġ(φRc��.�W�G��*�$��V�Hړ�7[��έ��j��/Vx�㊰�̈́G;��&�[�Ĕ�;әu�����{a��yyh�_�_��	�A�'�/Lg��z�i��/ӔEW fssjP1��+5|%��O`�<Lm���o��4�X���[`z���ە4^�ݼ�Z5!���(��+qy��3�s�RN�=ӓU. ;�� �u+8�d�d�=�
8;�Id�B�}ߋ!�U?�^�b�'DB!����I%NאL�ҷ���v�n��CfP�N��ٮw �s]���p����l?c>�̍׳��RlѢ�k�ƿ��n|0�?k��UX4�K���a�����E�G���9(�3���K~��,�������Y)$��T,�_w�B��s⼓A޷�]���9D���nB&�#���6�Q�����P��i�����H�U��Yj�,�;�o���=���4g9����i��+��O�.f��ꎤ�i_q 5�h�A�}c6=SoZ�&M{�1Vn�2�2^���R���֣�ot��f(����m���w�~�
@6�{��J7�x]���ǅf|V�QF���:ފ�#�=�CEck]
6����NmF��nS:��������e�����.DI��*ځ���¹�L�j��c�����T��\�C�����r����e��D���I��{k�'u�����<q�5��F{h��-��_����f3���HV?�2�F�M��EÊw��\�I��Vj�vRbי͈�潺Gem�������������"ccĘp�d��%��R�ԃ�+�e��+�"_ֻDt!]�yw#i��֩����M]�(akv�m�LXt�����a��C��,��7��C�_���jH\�h�\���d����"U���Bm�2���@�Ž|����Q���3>Pc�t^�IP5��぀~1��^x���!ԯj�y���Ke��h*�n�6��W��( ��̻c����A�X���	��q���̋#�����:Ib���¥��>=ʐ�����H�A ��mE,n�C�<�y����:f�v�,��EYZ
3&9�=ٕ3Cj*1bU>,�	��;lp���2�M}�3]�x0��:�t�/�Sh���HeC ���P�u��wr&��/��'1�B
�I+*�D�w��Ȅ����	�<��jr����޾�o^��》�t`�|yrJ
I8�H*L�-̓CT u�׋V�)�t�ZWx���|d�_�n�\n�46$D� ok�de��1 ��|�F1���,$#]~�٦�M�Xs.�>�b��O�UB�%��5����Ϡ���O��,�y<�6NʪO�W��W�)��ꂅc�?��5&�6�e�G�Y�`�k�U��e���\K-G�w6%�~�ۨT�f)�_#�h��Vn5�	l���SA���5���!��{R��O�:I�ˤ}9d �.�����{(!��0�/�$Vo]n�fPL�%Ӗ̮��조Ed�]�����Y-^���v��E�:�KA5�����v+��K�?�D����߆@�Drʆ������!X�×X���q���?�6p��N2m��8L�Z�d�u�k.߻��8��:�~F+��G��x"#����d�U�C����.��_����L�p󒃫�G���p�7��a��%28�,���H�q;!�LC��@]*��I�fo�*�J��ۜ�^�"d�[���.��W�5?4twW	�+W����ע�4���w�+�Ȋ԰��eũ�K�����:p�rh��&Mw̫�?�@��/)���Vǳ��
9�sj�b���<��ҜM��R�>��jz�gtr.�5\�� ?R�P�"Z�a�k�����b8��'��=q9g4X��"�XO���:�S.��G�ߛ�m�Qί!�0y�!������ z�i�Z^�s�wR�AD�Y4�m�vruk��~Ԟ�LP���7S�F�&���s���(|g��f��ëʢ�b8���0�l�U�u]6�s��:s!%�ec�����l����[�!��]ő}8�Ѱ/sJ��͈�Pu�Î�O9=GN�=�4	�g�yZssZv�C�t���;h|�Humx9���\�� }ϊ��pė�G�Ek����&ݢd�bv..�0��G>݄l��0��k�k��d9�f��v�?QV~/�e穵�����^�k��Hlh�����l)̇�8�:SiR�&!H	ԓ2V���T%���e�߈��+[f"@���	�,�`.��>�7�G}�2����`��h¶�8��y��n>�K%aM�Ϟsk��<�f�Z<����	�'�������HZ������b�#BP��AwY�ę[�T��rސ}��+��铡?��{�-��#�)��"����}V�6į�QG����[���dC�\��<�P��b�m�F�����ِ���f8Ȣ02 �5�c���8����6ZƵ��]�D�p�s�=H+<?�1��Rh= ]�r����S���=��=��j���D(e�DBLǩ*�!�7�/JOW�IIep�ǀ�=�]wܰ�鯬F�����J���9Ee���ء�C�-�I��i���V��C�W~���yWIU����s�d��M4D�౲�[:�&�E�'s(�#�df܆�\P�h�l���c�JGX�) NB�6w�����8m�&���8Y��X�G�Ą[��r��hW�%.�{s�pCj�'8ro"bY���t���g$�׷ʝ��H�(kE��k6�Υ��+Z�2Q
fF���<�V���@eTi�W��~`��5���:��m=(�_N�R�;��`ʘJ4|��Qʘݙ��p���Ԣ~��_�jK�]�|yg�G��O���B�(�]���|��;����H�����:�6��ߓ�j  R�������++�VW�R��z-�m��QF����S��C25��c4ʒ�<G��"�`�¶�{���t�;R��Y1d��h����7�ő�$)Uw�C�&�T5!�_��f���Ξz���I^�48u�K��Z��(�q�oŦ4k�h��x�VN�(S�6���#E�| ��_9��X��3�\l3K*��Y���V\�����n\��R�f%J�D�(%�Ş�B�0���a�x�5i�h��|)�<N�����ϲB�&���s"���`�I�����B\�|�ƨ"���+S�n�m���r���j�v��nV��wʅ�}9��jO�|ɼ�ϢC�aLv�J�ˢq#ԍ��w��u*f)�ymT��N��a���x��@f���n��[+`\j��Ɨ g����jz.z�S���â�~W��6^նx�yLk1ꦪ�g ;]C�	�"����?�;C!���}��.^2�V����Р��B֨��W!'Y�s�Ύ<NT�i�'&�>6�<'i���[�5tԹ���[�����rpL��_|��'������(��t�s�+��0�7�a`3�P�X�a�����Z㒫�\`���ӝZFb�oi��ߔ �H�*��@���Q�$�H�s[̽�0G��Z�ɳNQ�$V.l?U��a�ʅ�YȈ_:5������������D���X�&ME�z��BT�$���aGĽyP�4�z���̮}�v��[����6�34�/f�|�>�$�l��)8����\un�o	�S=줰XCY�V��*�#Ԕ�C�z�ua	h :���?󾳥�����K@{�����5m���oS~bנe�����j_k�B�.k����t�X��0�s�&���q���#����	v��	�ۻ�����I�s�9ZG��2�Ƒ��BX�>؍�
� ���<��������7����W��0��Ё�x�\T�
�	�	U��O���V�j
�k�R�g�L��.�S����H��+�i'jځ{�]邑��� ���A����׺ ���`��� {��D�pB�!�$�H�u��9��v&$�J|��Xb�Ҭ�H��ޜ8&7z_0��� �(D�.@:M�e��E�49Ty���ۏas��A�[�� �#jIY�}��c�#�{¤r�?	��"�'�� �0=/r����Vފ�w3�*�ru�Ψ$���-#�v�Hc/�Nb7�4,t��X����7��\(|Pmac�_�3&c'ժ�=�i]���>a:5>�� I"#�	���0v�'i�y��)��	(Y��7��.8�ř�}���b�S�yQ��#+mV1��6�_��@�6ɷ�*-���z�@�P*��-*��E<�G��bϬ�j�w+.ѥ��|]��2?�	g!Qi���=��#lV_����=r����[L\I�Wk��_krh��NG�?Q���Jm&�����cP�_]���Se���5ull�X��ⲏG����顒������p
D;��GJS"�D��k�+F��4�2�\���;����@��CM����9���ka�j\h0��{:y}��`�D1�ǫ�c��W"$4��,T�b�����x|�iw6�y�BZ�[��;�pޢ+6oK����(s��Ŗ[��x\@y��~��?޻�^v��^�ɩ)>>�jQ��I�:��v���4�Dܸ�@�\��+U"$�s��_~G~�C��M�K�*�z�G��k.N���������S�Eӻ�HC�ZHX�w�zq���X���<�����}9�[�X%�dn!x,b5������nE��T(I{�<s�V���(�28�)�秤�{��b������C*�ϓ9��M$٢�oW��('�TĲ�O �o�#;{- ��2K��F�'���ι%�e�V����T�?g�_�e�'���Jy���w��Z��֫�о����(컘n��jґ�ԑ[���I�Sp��c�3��'p��'.�M��lk��������`;����D�O�cQ� <	U��t�\��(Ab��2�r�L�*X(}�_AqD�A�h����@�K�˕�xIEf1F�PtST�H�k� �yE�gbA�G-�=<P9�2A̅q�)#����B���ogx��Xn�y[
����|~�]�\�)��-����Y���L�Gl�1!�n�D���j��e0��P�W��տ�3ebV�
"<2N�]���$�ws�a���NH��X2�F*
�K���!�iP�gB�n�{r��f�p�u�OK����[��2�uצ�
��z�W(Xz8�����~c��8Jg?�R���
%w���T|��ٜ��b���+IA�>��Q�C�(����|@��&���"���Y}9h`{
`����ϐ���p���&�S��S��]���±D�����8�Ǚ��T�='vL�K>��L}x)��N�������;%/�NX�G�u��2g���r��4���ԇjwE�-+	�"�j�W���>��
,��w٦{��by�p�vɍ�gm���c=�l�?췑d�U>�E�������-�j�S�9���}���gJ�t�����;7�z��n�t&���U0G�k[����$P.\b"pn�7�-|J��Aޭ���Ho������a51lts��\�Y2~��LU�Ӽ"㭙��uZ��غ�@5�,�}�S���f l_§�ek���K���2@�Ɵ���G*zT�����T2�(ޢ�C��;ڴ���Jk���Ė�0A��<�1}��z�V��s�|�ے�Mid<EO���v�(�p�Rtǜi��u��.IKR�l��_=`ir��;��+���۷�.�RX�����_����f@�+T�u�+��\w��o��K������#�FpõQq���5J�E�_�5�-�n�W��Z�^:x/3%�pBƓcJ�?��CMU+�x������<{(��
��+�֐@K�m�q���CDW	l��.�"�4�S�7M���r;p>̽� ���6�g�A~����+�����\�;廨hU3����iM_����ʰ�d.c�6V%���Z���!��VQ�+�D�<��h3R��7>=�)N��r�G���"~$����%�2�{#ͽ��9)��	�7D,(gB��.��.q��&�6��>������u�I���f݊��%��Ң���Igy��Z�+tZՉ�aT���CF�3��'�KC����1����e�Q��FҜ=�+-�t?Ǫ¿)B&;�I~~����(�_�b.���+�>"_�s�dPj]WZ@՘|ì�D'������A�>Rg�O�n�R�f��|r�W1��������������}}ω���߅�_�w��?*�ՙ�H���|9`�M�|%�ʲ��q۳L+�����F�yò�������ۼ2�xp�l���e���!"C<;�Ψ�Ùt����Ȭimd.����规�1o�?);C�|�_��	F@x�^�1%�C)_�b���`��	q�%�����$'��Љ�pU��Y��W&�����4-D5+����c�����Hd��ʘ�>�y�
C��GW�WÞ�xϪqG�:���1�ԋ���a��a�m�-�����N�dY�FQ����g��A�VB���[��r�'����?����E�??J�IȀXU-uz��)�hķ����p3�X����H˽��P@��dI��$#�V%intKy|��3\B��1�� R�3㿆[l��{2��Ȭ��/;
��V�f8���>O#G�w�P��%h�[{�\�!���	h���Io�,U�����,l��/�ɽ��U���>�a.3=jZ��6����pZA]F������m�)�{��#D�EнG�����*_zm��j��T�d���i�T��SU�sh�?�!�zU<Y�`�s֟�c�٦�ٌ���u&�){��I� �O3$��0��QSR*k�����ư��dM��Ѝ$b�O��^��g��q�ң�a�e�"��^����\Z��<*�UD9J�] ��v������<��!�3��P���t��K�(���-'�6���hH�vT�⎙���>a�E/�\�`�	~@	Y{c�]�1	��8�8�֢o���):���u'��B�{�V�����v�/�1V�Ka�&����f7�/E:�4�kڒ�XJ���"��}�\ˑ��4������i 
x���4��;<Ea��mv�H%~lf��,���&�;�"�B��m�){d��T���vrS�����Jfv��W�����*�u�@`�?�H��Ys��#u~��5��/�l|kQZ]��u;��R��a����Bv.����Pt�ܴ��?�a��w	�1��kA^�|�!��Fr��z�|}]�|������A�9�t���đ��4�[e���ICt��[��jW�xDJt��6	�\v�$��<L���'�����-��:ڭ��s��N&Y"���9h�GJ��y�q��R>svn�Iɵo�jqU0���LLq����U����}�1��D�I&]K���N��HfD��jF�z�����5���H�B�a�i)z�<����l�9]�/����WA�m%���~t�qQ;���e�םf�kM�G������_���/.�l���SR���п�ؠ��E��!^W-���/o�u]��Z/.g��,2�o��Ze��L���.��=��o�$ʟ�p���vKH���JF5��f�^�bk�<���q�=s2Z���v�����}�.i��0ȉ��E��9d�e�NV=�{��y�[�^!*?x����Ů�K䄞���4P��H3&:ד`_qf06��|VD�QZâ8+�x��>-��V�$����T&�ϔ�?7]�f-Qo#���>9�6�̐ �Hc0k�6H��P�[�ii���s.�>|T�g��Gt�[��T��>!>_���Y�
�����Q�[�B_��*n�7,W��ܲ���'���XaL�alT
�j��ڏ!9����wHk��`~>��8�c���|��� �M���y���;��۔b��F�m�[Y��T)#����⨟�}T���������޸�O�t8bi���ɥ�ђ������� �"�ǣ(4��WB�,SJ�"�o�qi츂��]�@�ߙ��b&�Ř�1��Q����Q-��u+�c��[��I�#�7 s�0����#���ڤl揃L��#	Ҽ!��`�˽LؑA��� /s� �C 6e�aߥJך=f�k�BFJ=��i�cO�������n#"�mԴgF�?M�����u+I;�M3'�2uX�觎��L77�-�����3l����Q�`���vp������Dd|�TGIX���u.ثW��BPj9eV�[�ɵ�df��x?�	����΁�l��$<Y��R�_a��;���?]Б����/"��m���!�U�����?�6�a#.~�إ���� �I9�ژ�y,E�XoM�Q��V@�����'6i� �$	��)L��1��{���L�E]��������V�9��}�NCʐ��J4~���lN��]xI�M��ޥ3�6��4O�E0�4�[��i��O�	��! ��=텊p��%�7?BNO�MM��xF�� =�ܔ�qM�Ђ7�)�������])�"���/<+U���ܞ���u�8����R���|�.H�n�'=OJv��%�O�7�̰��_���yq<r��b�F����v�-� Ct�(�3YAZ�"��ZG�>2q`PV��U�s��)A�X���XH�W��e��#_^ߢ'�1A_�Ԯj8��RYL��C���� ��^,�L��O��d�{��HVMǆ�hi��_,��]���ΜD��M���L�����l�к! ���}M��1���5G(��H��^��n�5/L���B��ckȨ��Vl���ՃX�ߐ��z��Ᶎ?u�L�
Ui���r�ѩVAb��Z%���Dt���D��ElN[W���`pdSeYV�k�Äl�˖�`�"��  �a�hy�>`�Ջ����3TvR$P����g=�յ/,�Z4���/Xٜ�T��P��-2g�p�ߑ����َ�y8���ի�K{�����̋�F��Ӯ�j�:�3T�*2M��*t�Z��߆][{ң@�a#TPs�D?�����@�2�4\��+����h)���o9c\:��V:�g��ſ#�͈�Y�+�?cu���v�2��<�;c��@��K�p�`q��)r�.W�{�V�(��tkQk&Qۮ&��[�:VƤ!�[Ǫpؚ�)o��{e[��ͤ�3r��9���O�\G�/'������L_Q����OGŪ��|�*|���S��[*8�#��Pb��ƀ��	������b`0	u�Z�|y�T�ѣ�͹Y����s(������b�,;x��y�o�LR؂Z�ߋ�/M�ɬ�ُ����+k�s����c��Q��Bu%{�R��}�y��z�%���`��޸|�p�s�n����n�ra�U�~��j�91�ޚ���(����֖�EA�y�Pfa�n������5]a8���&�b��6I�ʟ�jt�﹑�����}���B���g�Iؓ'Q�e����xs���6��؝�1mgS8/\�*8~z^T�qfqG��g��v�S��f����e2�M���COmh���'`�0�y=v>�>Ix������I�y��ay�JZ�(@�I�I�Dl�Zo~6G����ŦȪ�Bg})�@��Hb���8AcY�:��jTk!e�F�@�^�_��yI�չ4׍@����-&��1��1cK�{(H2�����S����N�;�/;���I�I]g�D9���{�AAa��Pq��l��+�O�(Ѯ�Ib��Xm�K���p�1��=B�~����S������ �+QN���V� �ԣ����,gr����bF�Q������D���r˺_#�/�y` �Ci��-�JX�差s��ă��cȈEl�M9���������-JK��◛ƧR�Lq��ng�*6%wב)������D�w�����A�_��L|:�:�e�j�Ա�뉍���bq�=�)�_��
���.���!���@mb�2UL��t��=�c���ϳ,�#��EAWG+ł���'�G|��$4���V���GފD�Ȳ�i�V"-�;
�Xc/?
���i�t%���� ��O�g�8�Z�;�\��K�:�#2�J˼��^8�4�z`T1J�z�h6�Wa�ګ,Qm[+�ஶE��xȺ������Td��@?`�X,�R��8=堾1`�'��g��R �d[�5�i����'�yz�)�q�'���R�]�3�N��BZc�a�݊�K�v�L���U�	4�|Y�.�τkZn|�$ho�i7���K�(!T�l��1[����ip�����JF5��Cs^z�B���E��}i�Pi>�P�or�!��`~�<jv�}�����^&�>bOS&���X�_�p�E\)�"��Vm� ��p���-.Z��/6}�-���4��G��/��*Y��s���S׾�Gu�X�M�\���r�]j�1tf	g?����/_������kf���ב'�Gi��B�}�^hE�5�P�ѹ(yj�* ML���4�� ���M\���)4�hQkd^�{��k8\��4�|q�n��C��#���}���[�6vߎ�:*�:�ZX�dWz���q*�I�>Ho��׎yr��M���v��*3=�'����-�hj���Rѿ\�"�4r;jx�'��Fν�v!��f("c!�\_cJ��y��:M�%0�"WO�����l;{�l��m�YR�`>����7��a4���Ę��4.�l�����샛Ө/п��[r9����y�2�^���'��_� y����D�0�̷\*���aW��K0'�@��y_jL��]�r��4�8���S�Mi^�ʭ��VL�����T�jY�|)P]��!����57x��*n���(]P�X��n�����y��@�m�:2��t7�t�ͷ^�9�;ۮ R�$�;��6K�j�LX�����ܐ5	�41q�r�H��S(�!a���V�mP_艑���\�*�!|��kvM� @�wRT�]>y�k���#f~<�>���~Fqέŋ��y8��a�F�3����y�k3�q=�!��1l;C�����D| ��Q�ij�o�'Q���������3A�J�I/�V�W�I'�>��T�x>GOF�A�Td���[�ݠ�J{eG�(cg	H#�5�!!�jr�.ya�o;g0	-�|����"� �b�B�/��t�d�3ϗ�Դ}���,?������/h�U�ϕ��!O����C�]�e3��Q\*��4)!�c�b_#@����^EQ#�M�	I� tAot�aj/4ggis���+[�_>���:֚Cb}y�����XM' -gNL���8���x�)��.鹚���h �q=�.���?�q{���?A]�h����g���� �e_v�Ά�b�G^���LJ�G�`��&>4<rZ���+H�VsM� ҃����7��V_F ]_s���Ī�~�h�!��a���i�lU��~���)߸���юTKp-J0/�VX��]F�������+�5#�q��ҥv�~3���7�\5q�(&yC��
������{^dF�|��?�0F��U;�4��O��:�����❒�ʩ5*oh���B�_v��Z,�� ـt_e?b�h7��,��M�R�x/�B9"�;��<��ݩȴ�q5��c�pǌ�q�Lo�yR�O��(�^h����G������<K�5�DX���3���~���A�
�-`����9>���z٢���1{[��)c�h6���$�K�C眐�f��=��3�i�NI�zmM=@�~O�խ�!�U2�C���k��ޡ_�X�Ҿ�I������sU.}��ziÖ6L���q�9bA$V��N 6�ܻqt�	�B�k�y`F�BI��Z��%j�A�K�9I�zmt|(_��y�v1[��/t�/زH��6Ze^I}c�C��)��/^1�9�_�
2��]ɒRfV5����7Vޱ0�k\���&X�a����<̒'��]�&'��Mcu|��L�e�Sl�g�_&<,x�Qs-	n@�ʜ�ᯎ�'I���;W�xˈ� Vrƭ���:ˬL�ɔ+�nR��yx'��u[ٷt\Z���
3K{��:NF|�=oh�	dN�;�����)
eCL>�"F���s+�eX9I�`�Nj��\�Kؾ��K�%*���$�к�\I��Wj�����̳����m�t����4�Z���P�N0І117���3���tx��ޘ�M��Vǜe�����(�Y�r4/��'�Ȅ0��޹��%O)H���Iu�&p7E�@������?Y����MTo	�:dA��f�ǹ�)�Ɇ��3Y��d�):5�-9"�HƲ���+�c�c�Z0.�"w���lq}=��+�v��'$�S�r�j<�g����P��ƻ�M���͸#fT�:�Э�E��˥ �o6��;��u��ԡ[xE�Im���
m��|�cȶ���7�	������������z�1^����R �ʚ�NM�*1'��ށ��צH����9�i��}K$�����G�6,���4'����@o��ZC��p��a�5�Kb(ܔ�g��<xV�'O{�{Pw�q�G��4^?�w��wr�Tc6�^���3��3�k�C���R9[1�*�LTk�����縻���r��Q
�X�����h�2����$>���'�I�ݳL?���<�+��k��?�,�174o�On��ٌ8�CUZ���P'����m��l� O��)�#�����-Ciߠ8A�z"<�=��~�|�� �����K��Y�4�,���nH�Z.����_��^H�o`��� 6�z+�I:���`٬���M��余��\�zϧ���`�ʕ5���}��b�W��/-5��Ns�=h�Ny�,� 48�
�+j��#q��H^��su���ýo��d0�cj@-�����>���rf��ʍG���I�ԇaϯw����*��	[�s�¬Q�M^r<2�],���Ɛ�����zJ��:�=EK(�T1��3x�§D�@��ݝg�U^�Z}��h@k�dw�%����7��(��hZ6���uO�Ӭ\�}*�(;˲��M�_6|�=ġxi�n�L%nD��C������K�����k���	�,d���E:L[&�ښT�H���=O�A��	R�k�z�=�'�Jk.*��:{:�sDx��Q����/g,�呺�H#�6��3=dm�����r�_��K�u���0QP�	�z� ��.�w����P9��5�b���w��J����ٟ$j�팴7'O0�@�:��Ө�Aqw��H]�)ZN���	��۾���Jy��e���5ׂ`�ш����'JM�| ��.�r�9]O�zm��� �L� 53l*��J��V�v\�ē
��C5z/\e�c�Ϥ��N�Ʋޛ�oy���g�eg�E������	�W�Itu+��3�gW���J���_K�>,V�y�ʄ�EO�rZ4܀W伅�|r����첦lH{�v&ej�z��8ˇG��WG��o��n�O@hd�P���&�5�g��*Vc��(�;^H���z�`.�J{�3n�b:X�������lCwU{��{Ӯ�8<Ө�ؒ{퓫�+�7�3.�^j�t�����h/�{�.??V}FS���s���
S�.vq�A�������r��z�t�0s���K�T�M"<_����:�k�#H�mL���Q�:�'%#�J·E��\�i>��kH3�D�ݏS�.��1�Gl�sZ`��L�5��h��K}���G�E
��-�&�=�X�W����=Ͼ�X��ʨ�a��c��O�_�NH���>#'�!�:�y�|������(��K�M$ۘ]̼#�r�u� ��S�],R����ӈ��2_�O�'�>��4~����>j�t��Q="���cw4�� u|磌��N��?Yl[h6��N��U����d�xiN�ܨy�!955� ��Hܝ.��j�~�s�_`��"���4Y����u<.����V�d�js�Z���UH`c���qJc��T�#�H �.�=Z�=��]��ZJ�N���c��A��ld7S��B�8���bқD�έ����/��5���W�FU5��.�A��8Hh ̀ov��ԕ� ���0 /�o�$��d��Υڻ�rYh�!I�@�hu{s�z\$m��]��i��$QB,o~b� T��q���B� YK0���U��k�����֠�]�͍H�9<�I��φ�=^��^����b ��J�T`:Dqz��YqR��lQ�D`�a�:s@E��r�[n���v��u���d��b�v4b	��T�G��;��Oi��[X*b#��#v���^��j�l��cH�>�O(�Q���I����O�"�Fy��nq���7rcS�"��G�9��zNWTa�Z���y�͍T�<�٠\C)u���(؍eS�0b�s�!%]h%f�bt����W&�n�?��U�0װ�o�^
'��M_I|�R�MUlq���&�{��y;��-y:%6��q���(;��	����X�X�o[̠9�1Y����n��S��uP��nA�Ew��\?�~��wh�f�ڣ�uUi@�AK�8'���u�i���3�/�)��u����� �vu��a��L���HB��v�`��ZB��r��b�O�+Xe����)��Z"���4� +�����_��da6�JaݗN���)�̠��s�W����?�,���R��&d��aX��P̻��@!��U�˝mH _n��8�[r��,�r�=��q���^�ݽ�F'�A�[6�\�*f0�g[?�Ŵ5xL�kȏ�)�_n�i��0?�P����dA�3�˙hX�ŕ��ޞ�4���Q�� .��̬ܽ�P:N��s�{�6j�q�S��AS�!V��M�i�T��{Ѷ�8\����@.�o�0��^y�m:m|���b��`k.�kj�k;n��Z
���#�׸����}�>�(v���F�^���C��9ЁK�G�X������
��	���������<;�@�^d�'*��G�ڣ�{��O}_A`o!4�����t��4���WNG�\~!��!^c��P �4QEIS�B�.��"���/�=���hH��z�Ʃ����iS�Ƀnӽ�,��^��a��l1���ޣ2��M��ra��<�:�X�@�a;	���B	���kx?B�_W8�%��˿
W���^F�mS�VH���$�p�p'�DWt`������A.S:�u�v�C�I�)��wB�S)O'�����C*-�v�^K����fA͕����:x�G�|6�j��ݬ�J�rbm�s���8Iw��h+��v&��R�Rz��`��S�R鈰�F����d>E�ARKuۼ;Ld�z��Y�ZJ���˟x/˾Q�|)�1}MOdJC�Q_Wݏ7fǷ0�A("��C��$��x�d/'	�Gyj��~P�"{��&�SQ��g�[�&L>:����3���2�A-^\�
��/�f薨y��a��gb�m�Lr�v3�=�c���?9�n}�����,~���m#t�~�
wL�PLOO�+���<RH&rd-)�G����ڊ�J��xC�w��Z)Ķɋ�O�H�J���𡤸�F��W�޼�)t��r����|�|Tu�y��Zp�6og��Ǌߺ�	+�p�}(:�9�F���
_f��Ts�1\D�u��~�WTߨ�+`��Bj�.f���pGP�e��2*e�1���u�,oʪ� U��Yg2MgXRIJ|)��O�_ωYD@ky���4#ZfO��\����f�\��ۂS _������R��h�;�izن8��r�����%@� I]͎�TH���F�΂*ɩ�^٣(���~	�R�S��^�c��h���!B��W� χ��bK������TqQS?���p����~a����νW�Ӿ|�a�ue�?6�7�Dy���n1���D�م6�<BĜ}�:����b(�K���	?oq�NC���\|�&��v�z�C�>�+Z^�r��0!/����//����u���?�hġ(��
���y�
�nj'+\��X�e�~`M��#����G�����n�(X_'���M�������ݫ�Ĳ�w�ߏ��B�)�/��)�dZ}<
��{[1�a�+W�|��m6��$�>������%�'�I�^�wM7��]O�Kq}�k�3��D�R��\�:��f����c3WGy��["6*�ji�����(W]h\57�io�&a����[�h�IhvE�ѹ����L^9i$!�}wf��X��s�.4sP��N?B�Oa ��OIV���B��׏rmPtX;;L�L�����]P	�r�*�tQB�)i�,�y�Q$�������`4't.��;Y��n�-����4XL�Bu{t�d"��R����ע�TV�� 	��^�U��f������%��xZ��`�?yL5m�/�K �_/Ɔ����PH�}D��g���c��� '���x�PR�-�Ks_��^�G�Uz���X��q$�&�.Ӏ*�LP������vP����}HU�t�1U��<��lQp���uH�q���Q@�v�U���W��f���|5&(Z�Sq����l�x�?��=��(�J(�U<�=���evG�]C�g��̷t"��}��Ŋ�_���%�W 3�6�Zh���������%�ct���[�^2x���,�晶%{Rj<��2�qo�TM������|"��N�-��^lD/����>uE䫳A�]kqC�)���]�quuj�9�S��P�zU!�[��<��`�l����5���S�,��&�նK�X����}��_L����^��Q6�!���3E��E�\oWq~�̢��f��X��JW���o��W�C%�U �y&d��d�`5~�cK���0)}#Jt��������&��;�0��z�p��aV-��M��·F�@���^�Բ�.+����L�*���L��ı����*QG��0~��h���>,���+]+*L[�b�0%����%�"�������t���+��gOU^sKv������A���B��"<��d�^y�8k����V���9W�}���"�@/���bi(@8<��~a�R.��Q��]�6�N;c"��k%2f�h(�"<LŠU�,��#.8��E�D̋/&H����lK�%��.N���������r�� �@|��??��U�3n��w��Բ���ta<���/�*c�q�ff˷���zѝ����m"�>�׆h�$�H����fwN�G�s�j��s �G:b�]�'0~������:珶$��O�\��%m ��%�K��koy�Px��ɓ����P�~�7[����:6��/�d��D���эN�'C��W��MSf���'��<T��h�gߵ������C�R2g����{�Nk��Za�_=~�-��x�W���O(��m�E2��Qu�s�"�P��4�Lwa˚�"�� 熴m�Y��[댦	�]��;]����7�ڷ�0���V��a�-/���R��K/�p�c׈��HZ�_[U�-L<�Ny�Dr���?�"���\�[v�a�ж�݂��x�4�`�c�.s5G�P��`��$����CK����ܾq��#�p��y�� !t-;���6G���O���Du���r%K6���5�8iJ��-�
WL����(�:"ؓ��d��,�@|��^*�NN�@�t(��,��Y�"l__Y��%́� �)��s=�VYy�g�߈����!�y�CNa��υ�;�\F&�A(���g�JְȖq�UJ�l��d�ڭ��:[�9>�����ZG.�_�m�~�k�U�5Ж�~E�sO-,N ���M���5�$o����'��m�4�2�d~���n�M+O�@�3��z�y�I)�y�䮚|҄{K�p�+����:cҤL�˔�1���{�y��õ"��!�U]�{�����,�h2VKQV�_BUhF�v)ی�xe	�IH��� W.u��{d}D�������\�Fx�ʼ!;�-�Aа��Z����V+�H�#c�\��� �)�!��7/��Sr�U1��$)w'9a�2`������5680_B��5\T +{��^���_8�s�s&���jD�x^�;D�-�l-C/T+�G�v�"�D�B�i�״fI7,���k����u%R�{��-L����f��d_6���7pӣyJ��[HC^'S��/�$f�["�
�=+]V��=��i*ro�3�ۡu�rے���?�H�MMKE6�^f�"��#JGReNs�DgO \#$��H�L���|���C�i����Z|m��
�u�H��Ɉ0]�)��q�j�M�p:Z8�<�������'�H}��l��3D�O����7�v� �1�'��HI�ޡN������R!�y�X�^�=��kl��~��©���^䯉! �l�IQ�K!�F���.�"lh�jA�qz�� ���f��R�5QCRY-��W�{ob󛐟��k��0^!��_L�s"+	����{B���Ȋ���:���f�Q�����oa:q��c�W�%������s-��[EV����06�$�O��^x�2��Lq�i��P$�O��D��'0�U���)��~��p�W�ۣ�ҿm;GVTVFS���q�o��c�f��	P�~"� 4(TQ�9���3�h�h��x�]ݮ��P���a��ɬ��}У���Q����`0�����l �J�ty��N��[u�0��L�O�L^��(eu�z�"ԁ?��qzxK	(�  ��;n(l����9���O3�5���*�,��������7l8dWd��V��BMR�+	t?�7�or�?�E��'�3�4ɰ�K]���V4�n��d9 @	/�e���b޹��b��#X��?��1��cr��iD�Sk��N;���a]X�=sIv�{�F�Db'�3���G��g�>��g�{y�f����q����3j�T�#����Ѡ���%�/��|`.�~X�3.=D�*����=�e�if�v"����0�L��񁣾=��;�O"(�#���y]�6�3(�%�<�P��X֧��dv��`�uP�1I\�`�=����d�E��uwO�^4!4�!���ʀ�X
��4Gu����_��NTJ�G����s6P�#vq�J$�^fx�!BX�&�@.�d�Bq��Ě���l���(���Q�ʋIR7��F����7^�fS��;3e�_Q�1LK��7D�A��$����!`��,�%ⷫiui��LR������Z{s[̳���h�͒��$��-��"������f.;}8�{]%��sn*����]���~����
y�\W�@1I��7�3y`�j�@�*޺)]�g���&�5[5!a��6� ���=cc����e�yS�tx��*Z��5�BF�a���5�Zs�~�p��K�Xw�Z��
JVA���y�H��W��f�F0�Q���8_���0ݑ���>^d�c��f�f�IV)%���nL��*�窈��?�3��!$,j��j��C�E!��q��R(t�<�����|"ԭ���O��aᰒ1���瘃�7����i�����0��6j��,�6�$�艧h��8�B��E��nPU�f��.�d0D�F6�8�{U���a�����ǒ(|���,�*-�U��]Q.�4�O`A����|��\DTzoވ|J7y�W�7��@��:/��{�{����w���􀩤��pe�# �>�=*��R��~+�x����M�t��m��� ���:�Ӹ�g=ǘPV6����|�Rsz-��ŏ)���N>�ɞ�d�*W����g��t(����3�(x����a�2��4[%�aX����x�Q���$�(X���9U�������>/�"�M�9$>��"�:�(;��{c���ݐ��*z��F�NPK&�H��![ˆ;4m����ew��P)u�ϭ}�c
P~�>P���,����n�"�[]V��;�J`Y��a�0a�>�:�����I�⌖m�9��H%���B����huM.i���Υ��s�i H���@��%�Y\���,� ���-w��������{\�9=�7h���k�9%��[�/2w�Й��Z*�I�L�хen����_������s׵�����,�3܀Սu9OR?\R��B,X���6���fl<e�[���7eNG&���3�x̝[��7��������Ԯ�� ���p�2;+b
3u*����D\�P���Lت:X
�N{923֍��#������0��f�� a%��8r��k��AM_�]9*A����t��m-�+�d��޸��a�0�ݮ�π?�!�>��P���N?4��T�ΰG��fHu�1��1T���~�v��*g���i-$��a�	�<O� Vj1�M��
l.�w����xze�p��(F~�2�(z�TdM���� �N/��f��>Ӧ�����rB��C"��a�/����C33�9R/{;^r�ȃ\��Kw��2^k�;j&͚�pL���%tq�5�
�0�^a��x	$E���h���_��Y�vg��~�[
�v<9ǹ��2��pZ*