��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VYjf�>ρ�f��W�&��$�B�9q�!|n߈/&�4�پ+��sU�9��p]�H�ޏI�(`�R��a��핢�L��4b��Ҝ������د�C��y�h�g�2e]"�;��͘G��9d�������Pw� ��:B�xM|҆�L�����~]��-G�,�Jk���71e�|�z=�}�J3��.��.����Q�MF@�T��Mτ|Q�8>mX�.��͇CgA����E�L����L�Y�9�Ů��S݄�����TG 2��H��+�H�����x��5/y�1�Vld� T�(��ٵ
Zt���$�.�ɸV�,��wpV�Zʽ����#;C%qMf?��Y�@b��3�)C�a��M��~�����X��M+=��A��j����L�+~�AV��f�T�Tۑ�DI��Y��96J�}��;��푾���f�Ѳ�A����������2!f�s�4�b��I��g�/"�	8�I5wG6���n!����!
1����%۔��˝��%�Ti�]F������1�>X|R��]{��`��o	A⎹�Z��B����c�[�k,ַ�za-�P%����7�x۶_{*>`;�9���]R�Êg(ШR��3d|f�#%
���iV��S�۝�SXg	���į���{�[�(W�=���5{�u�񝲬�H_�oU���� �㌶��ި{���	
����J��?�}$-�S���2�#L��\rj>��7țwX��]�����f�������)'h�j�~��&��b�2���.p�
\h�-�Ժ�-T+k�<wkj? ��(&+T|�FƉ����{F-�o�(��q�����f���'`x'�������s�cM/p5����ex��G��<��6��q��S�q�B�v��#�c=�LU�MZ!W��M�����Yy��Ϩ8A��߳ň$�\*�w����˞�Q����腫���DP_�t�r����o��8���ф�����T"6E!k��c	-��|�ٖp}8ɵM�4"]�9���@7T��>�:q�̕ɴ�����.���ַ�d���C�������f�S�UMj@m��G=y=�L�Blc��<�qR+wJB�K�ud,��e�nq����jl��~�W�-� a��o�0��L����p�>��o=M�3~צ����0K?y�s�16�w���Q<�.us�_ ;���ނ�`s:7�U�U�<zq��(2���J>nr�@X��婆ohui%�I�
���$�(�ɍ�p�J%7-+rlv��v�Qݛjr��2�k(�#nJY�!���ҷli�[������3G����`��1I�Q���:��eG�ą�j���g��J�)����9�z�Z\f���]��x@Y�=����t�(�or�}@,kmp}��oCePn�{yĮ��_�h'i-'w���::L�=}���>�Y�w��z�\j�4YH��O�[#�Z�#i���h��^�C�P���-����:Nܳ`\��86�ER�a�(Dc?��$=٦�E!6,$u��N�`���,O1[���>bp��z��/vo���}�_mF؝F[����|��������⛍#�v[I�r|��l�"M�q�C�S�|U��.�6���Z9!?���%��t��Ug}�+� D�y���,�s�C�vs��u<�*S���QŃ���b(N���y9�%O�d��G�7���v��y� ��[���x�� 2�$��g�w|�w��^Jnn�K���n7�N!�?YRF�(���z��<��;��=��ި�����-����0À�Z*�/!�wec}�P"h�d�ɮ�7��'�����҆:�z�jZڐw��<h�<���E�ۇ*��W����XA�}u�K��q[P��M��_|����7��N��F�F��.�3��Rܳ�7,<��k<�Q��p�`Ĥm� a��rCk��?������h���:/�V<:>��#+����$b)�h �t#̪3u�ԗP��!��Ph�&2~�Fx���U���Z6]`�J�A�HX��-a,�k�x� k~w1���X2�v���j|��us��fڢO��2�u}�ҧ���!!O�{kKv� ���{x\j'Qd�K��h��G=j��l*��E��?;
�	}"(c@���������b8Kׄ4�P�6���p�ןk�/^�쩄�'�e\����>d�9"_��z�.L�
��3�)Dn��������a+
o�28������j(H�:E����r�u��BF��JC~
�L��uћL6��Q7���"!�FF�d�=M9�&�[$0��
�����0��N}���ૺ�Bo�$�4��o�a]� ą+W����;��jvIXfq���B��s]�3py�%08?LwҶ3]�l�ְ;�͆ �w�����-�鵮��{'Fi�:�ޅ���5bā<�:s��Í��b)�M&'��T�~�tE�8�~>��b�r8/�;h��ET)��`E&!������3`�sy�+�X�����ָ��T�iW���e�M�)��w���j	#��g�0a8�����-8B3s&� ,_I�	���E��.Gmq��~%�-���2)�Oi���6B8���a�{dÓ�N�4�V��@�5Um�q���I�:�v!���7�*�X,�[`��E?���9�gj������_�e�~�ɞ8krdp�	C�G<�[vV ���������g�W�$�a]�E�[����˦��vVњ6�o^�P���B>É���jE!젍}�0�_���3U�܊L���$68~���q
H4���%�J��0�-�8�0N�-|�3��9&!���>�U�⻛/�WT��,���h3+2t?t�/�2.���?����V��7m�\)�E<ᓰW���=r��C
���-^�c�"�:`N$o8H��/T3��)��z8Uj�<�t{��Q����R��`5q(+������w*��.b��O�ԁD��T��	��r|=Z�c�t�� ���1��=��;�&��5���2�~cב���A
,���ٲi�0� C�28��1�9q;�ijd|,w�a�[�J΂�J��MRX;5c�47�Syq�C�:K|8ۃ:�	���{�D����0({��+��H��Z|.5�N��`�>��V��n����p�fG��V/��GgU,J8�)�sR|m����Κ�|mut�'�����&�})R�Y2�zt_�v�S1�<��={I#r��q/ax�:w�/��1�e��1�4�Vx�nt��a�vڱ�6�P�@¼��VZ����~d�2y�Cx��>�/�u�O�0�sjC�(R�L�~.UZ9
A�䀆�E���A�.��Q��$��"�gC>2�Ē���Kk������|�)�<ɮ����W��*Ȑ�_s�r�5���M�>^�׋Q�J�°��DHP�h��g�����4s�]g�"��q*�����@�죧W�N��f�ɴ�x��i�wȞ(�u�IL ��!7Y�Ď`{������hN�z�����\"�	�z��:�o�k<Ľ�;ԇ��ʒ�b�w��4��S���|'A#�I��_bQ�qQ�L��I����	]�k����_<�wdS�۰Oo���b �����gϤ�j��/��T��$� %�C3TG�6��^Ȓ��V���w���~	����t��Fp$=������uz����|��|�}�����N9+H����l�å��"5!c$)��xa�6~�B�����j��i
;�Z�����>�Xٷ�ȏ����B�{��UZ
k��Ps�`�a�v�ё�lǮ3���p�n��,)yI�����Lٯ?W_PP�fٝevҲu�Ʌe����4QP,!�X��ZH��ЬA���F�@';���X���)��&Ob��=Slvi;����;.ز\ �����T`�2�������������j���-V4�8�GF]���/p��S1 �0���H��Qt���d���?���?!+���&�+>��ܖ�5�bҢ�q���<�լ�����;j܄�"\�ܺ�;�7��ȓz��R���ㅵp�@%K�L���E8�p~HvS��t��Ll�.�#����0��e�ю�l O,��J渁ɋ�S0��6Q�]3�������\��/�s�>ɵ��w�p�1םy���E�p��&��ڀkG��	�ڶj�g�!1�H��ݏ�cj�Kv�o�`��"eQ�X�N��u5��?���e!�EWt�?t���$
-[��u���#�A�I�����l�e��y��'�����x'R�D-u����t�����n����՞�����|�<���Cׇ�Q�<2[���W���	2ֿQ���:�ʍʡ�g�Lۈ�	�"$���S�5p�j���$��ڲ�M�fAf�öw�ǌ�3G��"��<���N���7�����@����iY+]#�>��H{�/&W���6�z�V!Da�՟0^9i�'Pݭ��P���;��}�3)��� �_
�F#r�^Ctw�$a���H��r�[�V��;b��=� u2��M.F�?<UT�e3/���K�+)�x�]+<P��0@N���S���,y�v��^���M��(���8��%���t��l
�K��5&[�ب>�hT���t�����(�C~�̘9�#��� bZ8=�r�����\]��w
W�+�+ϯ:vdpX&�ix���d��p犙>Enj�2 vS`���C������0��/���(7ێF�x8�J,C��W'�����m�k|���Qi��z�4׭͒(&�-�.ZZgk�Bbȫ{�rV�X��`@w����ݷĢ9i�:�}�b8���:�M�SF�	���=��UA�T��L4Ƣ�.��2ukU�d�MC���TO"�|x1[=)�����쓫�h���]ZV�2��w�H�"��cm	�N�0H�=�,x�h�~�Q�:Kw%�Ó;=�5F����`.ˤ'��/��^�9��B�.�����p�p6�l�/�p����WE��Uu��{A���bS�֛�(����Df�J�hӜ�OW�=�]'�N�n����Gpk��$]6��}m�>��)�� �9�~r8�O�R�h��o�T%T^�a���0V�5�=�7��y�F�KΨtv��CY���5^Cn��{_:��{sgŁ(���3�}=�b���ܸQG� p����UҤ��>�ExG���Û��a@�n�l��Jv'�8ȿ ]����rUc��坯�|��ZI�-ŋ��JRz|�yiGk�*��.��+��a<�XL���-����h�����w���?�O|.�,M�F�o�D�����Da.rwcn�� ㇠ir���`�2$�,�Y�R��oO���)G����m�c�j�9�DJ���6[���������)�"�d�5E:�߬�p��Jʪ^�;��BJ��A�k��nܵ��1��0g�ɀ��o�P"���ڷw0�,t�2���5Дɲ�g�r�����?�奇:ג�!�9k��Z�P�ig�C��1.!,���O�7L��x�Dnug��η`6��E�G ��������<c�~�QEM�P�ǐ1X�p8ye�.xʎ�����Ҫ�]�)t�ͮokf�ޟ����5w�����e�MR8`�0\d�~>�1A��Q�Ӏ��p������+>J����k��l��
P���I���TUT�/w���7F�QjY2��y�>"(�8M��kK�i&ꂌ-�pd�8:<#�<?�(���!g���;�%�uO�56�Qj<��i��Y}��ޕWd*S7�A�{GXX�-l�Њ�3:�ݹ�(�V����r�A��O�Od�����ٿ;�'
̪�B�U-����vUMjÁ�T�s^/� �~��y�CFh����x\��(!��D�/Wef��$�k��c�H���������">؉�W^-����r�^�k����J�����D�#P��^�ľH�^B�M+/��W��x?�D�;�.�`]b�"!)�"Kg~U\�������}��>"A�YډU]凯/SD�1��B*�ǪEd��6?�J����� �L?�Q��h��#^�E�C�_���ި���d�r��W�'��5��7�>��]�\3:�f:��4Wҷ�6��)������γq,�sļI�6`Dk��B&�ʡ�3�g������?��)m��W43� *�~,�ax�y�`&eUŞqjH�����]cw� ��[���E�l퉝�6{�����"�z���C�$����&z�/E���Ϟ)C�US�,���^�S�A��Z ���-���z��X�%�Hܷ��_105����q�ef�/�̭/����c11���NZ��#1�$��Ej^��G;����1ہ��WnF_�?Sf��=c�I�6�@���h\��ILOEL���燠^�ye'>?�uč��B��7i����������1�.���ᶭ�*%��h��j��-���]� E�<�pD�ml����DUU��؂ޝ	ȸu?g��W�8��0G��$�i��gV7� �s��uĪ%&2�ڡ��콳�ie�4(�����zá4#�-[L�*�%��2	�i�yk�Q��Kc��W�z��l�O���UpR	�9����\��^��fkhu�4�EA�� ��w�Ԙ��4?���>l���p<+c�!��S]��CM$Q*�P^��ɥ���r�ڑ�Qʪ��bІ�H ��!.��l��)��ߑqp~�:�U�F�@�g*)�I�j	�g��sܡ,z�.���6�БCE�[���ޠTT�g �K������}[7GI�W�y� z)���Fو�2X�mrDh��/ǃxE�~(�����f3^ �c̮STbN�W�����{4��"�n+�zJ�lmKa�;C�`z�Ү|�I��Â�v�;�}um��h�[�X����(̛zp����t�ћ
tCo]��>08����I��;.��VW�hN�=NEp,�<�iٌ w$+�w���}���p���i�$�O���{M̬��_L���ם�4�QD�x@+jF��n�L^)�����  o1��ʍZ��7n$n�m�_~fc3���=���2�>�����m�U�c�W�,��W��Pf�o/֞7��غ VB�ܟ_	�7#gYY�t��[)}�.�ƎmA��I�$ɏ�oۑ�u-��-$�w��T��˂^k#���mff����F��>� ��i������x���*��G��f!=���כ��\�� ��(�7 f� ��/)� ���?k� f���?��%�('��º��"0�1�VG���3yH;RE�`�MqN>����;۝�[TZL60s8���h��q �C����ծ���q���~ce�
���>j�wE3��ԃ���]x�=�]��3�Vw�h����o��RJ�����^&s�K|���l!�y�g���b��������"p�ȧZ��~$A2�|Q#�Qx�7�����@���S(|�dI�-�ē�i��$�W]x(�iJ�����F�ʟ�)n��-���I,yP�%�"�o�[��"���(Nv��^%3��N�����8�h�n��=�
T)�I�"�K����H���d������nîD�e�vH���ߌ'v��~�����<hk�l��x��Puc<�`r)�z¼z��^�pz#�bi��6��r�t� l{zX�;~3В%4b�򓩌��-����㲟tW��2V�o��|Mx��Q�j��	:+@e*`X�ę^TH���U*���s��p���>LrS!�ҕICs�I�[������F���G��AE��3��`J)2��T܎TC��?;���(ɫ�@D��@K)��vY��(����g�Dvc^©K3�m�#���[�\����Ku,?��b�o2@No�c̮.�s�`<�˷Z�����k|�� ��DS�Py��A/��#ˑ��:�/���B�ņǠ'u�Up@U0����X�9Nba3��m�i��N��Z3h��)Y���w�����ҙ	v���G���O�@��k\JIQ~��1��Y��h����;*��҄W�+�&=2�5��I ���Z�8�� �����Ɇ�R	oգM�i����0�^�L��&T�a�h�W�8\"�h�K�p(Ӊ�v�S9u3�qa9�Ҭ*ɕ����O���K��Nl�[d�1<�:\��&�'�#g<�[�@��������lb����ڊ8a���Z/��w�~��V7��h�������n�F����`�� eɀ,}A옥Q	��D/�|�(�9��H߼(�A?�"d�Y�}ay%�5��%�뙧BoT����g�"hI��G��>�54|Zr	i����FT�[�)lX	���Y�9�u/��d,��}WЌ��Ŗ`*��8��<L�yBnJ��Ғ���C(��)NGi�Ө�?���,P�>�HN��<�Y�xT�iި^S>�+hҭ�nn+�����n ����v햭��6�Dm���~�r�U,8
���5$~�*dZ�eߑ�����XҐ�E_'d�ϖjv
r7�z"�$ol0.r_3G��ᰧ�u� ��#Y=#�)��fykt\]τҾ���mv��,�r�n��t�^�s?64�a�Ԗ~y^3�[���9�^)�apb�g������J�ܑ;��֭bŊ-�L� �����;���yT�$��Ԍ��0�88�j�]Bz�8>���&4�� s�2�`�Ҋ�ݓ���6"��O���E���9�l���U�.B�F��8��v�M��%�J��.Ӯ׆���Qk�f�����a����h���Ts�V�be6*�Tu��O�$�
A�B%9U��U>��-DhU�O˥S2@v��V�\�	�Y���{V7I����>]{e��1^�2�:|e�[�9��	��Zz�36LA�q�K��)�(4RLǦ���B���ysC��k&�.�Dz���7p�����{I$J��ލ�ӓ ��4?�j'����
du����Hg�-]��	�8K�5эS��<zYop�n�-]"��;��4c�S�T�0o�wX)
�ِ��)`\B��d�U����ZR����u�j��2¹�����s����e�@S�ѯ��_�f�1	�o���c��|�} P���Rd��Mζ��ۺ�k,6Μ�K��m����ߕ��k}<��l�b�!/)]`�ɒ�������C9L/\B"#(�!��!���p�p�A�c�OLl8�1�}���T���u����L�>����yk�5�j@��!_	k�Bl�Ϊ��h{�p� @��o�.f}��Ր{����1�7*���96X��ꂊL�)p
vI���4j��z�p=v���/����2v
@�Y��C�ߥ6�9��x��C"���Q��PWۻ�|T���q�J���ɵ�@ �H~�B�UUjz��]�T�M���`��H�x�٫��J���S����mk�jTTk�"�X��K�����1dmC+Z�,����'�.Ku&j�`[a��p��iV
��� !	�:$�jD �,�'N��	5E��Z�`+8Pgs4~���\S�l`�ך����E�=�A��nr?3wZ�"dʮ����$��4�j�{M�w[ �x~;�`�K����DP���[�x�'�(�"�6U1�@��ur瓄��.9�gJ{����)�,U���⽉�G�=+�4��-h`ै2������2"�bJ�ߊ@��EF�����.ڋ=R:3H��Y�7��C�_5�`���;�Y�Ah�͠N�gVW�r5Fq�5i9��1�?��P���.ʶ�2v.p:��֘-�9؂����^>�L0�0���i���癚�w�=f����]���%T	���R���Ƅe׺ٚ��@��$kZpv�:�s��q����p�q_S�l�����J)�N>�`�Sn��d�/bi���x.�ۛ%{�/��1bK��9^��5�^�=����1$#`H�1��WY��'B�ɠ���Rp��O��<?�3���/K�5�'�o����UT�+}�����b�|^xh5qo>�������-�I�ơ&��{I�"!����v8�j��`+�A���hm��)B�"�:'���yې�6����Z�}sE�Db�nw�8D�2�C��lo竢�@=u�[Y�:1�_��C��HA#.�oc��Q�.g��^�gh:y���5�JPU����/��o����벊��X%��U�I¶�t�9��"1�l���.�9u�+�����=7���c��d��y0�`{���NR�=�����6�4 ��w���%�%��A��a�B��U��y����-B�\�Y�G���E�ٞ���7�<��\�|r�#5 ?�c�����
`�a�v��|^�$�f7���^I�:$���uɻ��1Yq+%��X���קäߍfQ���8D�)��~�L��UL2T��Z�J
l����]@P�,+�> �ئ�����Б\إ���˙��l��X��gue�=0nN��)�Є��qK���ZQKM�]�`Ws��i�	3���\G�{}Pe�����!�ʚ��G�boS(�-A��R`T2���V/ Ԇ�C`��c+_Ԁ�St�G�Nr�$C�`���7޺�:�<ar+y�F2!�KGT�����tU��g����~<.z����D$C������m�?��_ެ�8�'X�W{c��۲�2�Wˠ�b����CA��������dF���qZW���'��Ŕ��������?�!G�ڛ$P��y��9�}!#��
�A���^1�B8����W<�5��)�ӏܫ^��B�Dt;�N*���Y��/�ՠ%�,Y�
T���K�P��z���c<��j��t���9Fjʔd��0lR�� �A�hٗPxi�D��*���Z�F�gםQF�	c��ԝK̹`z��sf�]ί��|��Tn��n�9b�4����N�٪eE�J���Y�d݆����u=6��Td��>ڧ.����k�:#�hιbsg�qs�R����?1��d����P���3�|V�I a�Q���Js=S����nYS�mj�>��n� �*b��>�>�Hj̉5͐�]��{���Q�4=��d�A��<�~�"�,�%� 8칁xp���s7��fd �yN�tg��Hyγ���Y �@qwq�i�(Щ�������@'�t� �l.і�������:t�D���Y[/Go*^&yMN�[!z����2�|1�q�m�r"\~���ˡ" �ډ>�'|�X7�1��J���q�� P|"��������j�Yj-�F���c&,9��l��[,�8�2���\���o�޶�g�Ŋ��HVg}��8Y�O�2{H�(B��Q��;p�]����*��}�����:%#��Q�A��HCM�� �<'ݶ����\��T�-aa�x�F��6��j.�9��솚��
�z-T�6ͼ�4l�Ŷ���_�FD��j��`Ws��� �7�8�9D/1=/kj�`�YK��%Ru��3��J�huk-)Ovʁ��������%���h�Lp��j;f�"�^C�QXc�w?[��'�^�NK#<��>i���,H�a��&����5*�m�!|�˹f��ێ�}-�w�C\[�{�*<P�>�
���Z���W�+:��t|b:�����]�^Lh`��՚1��/��Z�SX���,��x.J���uݨ��y���p�-j����I�����8�h*m�!���6�B���`�{I5��fy���ع5x&�,�j�����^E���s���S�p�]�^�)(s�Uk��V5�����I#E��o��rh^7C�sa�]]�y�>�.��y�@��@�¤�@)�|���=�ܘ�C`���߯e��s����^�?i�0��jʷމ�[��>��������qo�Z�n�h�̪�E�јy�l�������N~�9�߄�"e��eT�9��s������앴ۜXG��Y��<�U�?�~�M�>`���Im,}���0��bq�i7?E<�TXM+vKE� +�X�F�F>�� ��{t��e��[_�K�u �{��퉪�0{�Z�<m�f�Y�-e����V�ݏ���ğ�ڜ ����ʌd_j�I}*̗��<����,�i��k_F�gG[19�*i}�ց�# ���áȷ��e�\���"��V�ӯ��)9�:h,�"��~ׂ�f��+p�o"��H��T������
_�}�[^�NF �0�It�@T�<��gQAn�����/��
�P����y�0th�|�0������YĠvy����\�����R����Fݔ��(3����l9�̺|�ˤ��
n/ȍ��A�2�}ױ�N)� ����՞������PE��*>����s,6��e��u�Z���б��������)��!?��2�ǵ�@�%�SwoS��Pu��WIy��Or6���Y+�1���K
�H�N5i1�4^��M�����_GT>�ǈ@�/���
 ClRx�HMA�F���g�D���F�����&[3���\��^Q/ �b�>�vF�����=���Ntf�}�I^��]���A����垄�i*����=�Nr9��ۘu.]{[��41����������yꂽs��^�����ױ"ע��f�+<w�� ���3UpO21
��?���?�(9�{?��1��Gg��)r)�?�
�6�O97�^����T�Ș�!ѹWRY�kǷ�ޟ:i���'Ѭ��{v#��/�fF�a�N�x?��2}X K~*ۻw�(vQԮk?k��
H�SSe2#�qe0d��'˴B�Ge��D��f��nw_��ͨ�|���6h��	wP`���߻���	�/_��z�%l}."��d��T��<Jͻ^�󯥤x�&��1%#�Ի$�ɣh��ʫ��2p�U�Q�sD�%;�+/,�/Y�ҏ���������]�\���M���F����/f�$���Ĺ ��k�����t������U@�8lK�r(wD4�:dpC��\�8�T���@�%���ڨ�Ԑ�5�e�н���nE�
0���Y�r$�VP@�[�i�b�\�{`υ���6�� �c/��u�������p?о��X��C��-DL�����SU"������w/Z�(���"�b�$��I��Z�w7h��u\�05�i)Z&*�������'�E�=߱������&��YU �ؾ <�Q#F(pZ�h�e�K:΁�9^��_����j<=��Uw���X�V�A���f�On0襐���O�I-Cb���b��[�0��"<b�VK���mu�M������-|||�!���$�m�"� ��&�󡔠\.f������WJ��뎂���=e�`�(�� ����bو�iZ�Z��ѧ�u t�*��ƯdgQ�(e�����\��˷�E�nC��>�4������B6��.>���8�;�wL��]t��FH+��<��5�ஃ��S�q�V+Uf�|�4�U�Zwu�|�
W�/Nb���M���	F�b��<5�n'�����@����p�2�^z��Y���ĥ[Vj��ؽ��+��t-���Q���6�u'���V��+�Bf�,RM�paT{��0��I�G�v�j4�p�26�Zҗ�'ȴ�s_�����6qos��ˠn.�H1J�$�fC�s�1�W�����>m�x��/�f�_b���3�.ე菱r�u1�� ��Xv��.աb��J6�����8�P�YL��1v���:��-�u��Kk���lE��)EOV6h�*�!���X+�}�p�z��j�(���#sl�"1eIgkb�8893Pϡ)vk�D�_+�T�F]��V2tVg$�&r�)?5<����H4>�]V31��T�Y��`����n��� '��8Kx�}��U}������d:Rɞ��Nʚ(�G4��^-�߻1��et�MN��P�^9�J]�����U�"k�v���
�S�D�P���Y�rMe^���4���:Z
'�&ߥZ"�+�/:��F��m@����B%b�^O@��h�0���t�5��+F��O�ɠ�!�yI�;��������-"�^������������(����6�H�5�/��m�)B^���<�X��T���T��NS��7���'�E�x�#j�Q��8h@�tkH�;�}§]U����`�#�(�K�1aK�?�i�˭'����XP �5�A'H�<`�D�����<C����ŗ��MQ����P@�ѓ$�2E1��ܥ�����ECZ��OlH���Q���@(W/"����>|�����Z�='����\�m`�'�h5S�}��1�WT����\�xR��� ��=���T��M�f���Ϣ�����?�M��v��h����h`��n^:����l�Y�={���Ub�+n?��	��y���ۧ�A�q)��n�\z��j��H�����M��wH��_p�?���cx��^�#�;\�������H@�ڽi2��-�ecz������ {F�2����Y�e��&��|,����mg��V��彇s��}�� �z�.��C#��ғ˺�q�:�M�	ǧ��[�[�pl1:�M N�%(���h�h�$u�����@�&-����}b=+1A=����|�^�
_�%:u����G��>X�:�� T-��s�#!ʨ�tGAIZ��9���ˣ_`��q�u�����	�M�&$�$�Ť�W��c�z���y��Wq1���SD a��{��.m�0����l�w�U#�Ωk��A�������-��|�i^A'e��n8QvU�Ix-���F�Ձa�0��H�70����N�:��/�TH�`�y3Lh�+�����(����r�����L*�(�*�����c�B��:�c"�R�H����X�V�����h�K/#>۬�)�J�(��Z�"8�2�����Y&qx)�1��~�;L8����9�BE�+K�����iv���@g�˵I?k������b�`��g,,���󝿆Ox���5[^!}�� Lv1�Έ^�(~�'��Rѓtm�n�Gl\�V����!���7:c�O���i]Ƌ�U��v䩀%��oh����U�b��2�
9��A��v��C�#?���1�W��=��< �7���`st���~����MCT�[�!�/Hǋ�%�4W3�v���|U�#�_�ŕ.p[��d�D�UHr o~nn1�e�{O#���+O0u�M�̿����-��~�x2R}=fø�	�&bnT<���p:`��_f������\�[����J�a��g�]�m� l7m}�$��J������u�
&C�tW�d+��q�T�H���$}����[ئ��.�]�Qm����ϡ~lp���F��<m)}+��vLr�c��]��P7ȑ&$1�}��Č��n5DZ�qd��D�{���M/E�nP��"a�VJ6@Ĭn'2֚��T�.��5 �z�����=L�4j�l�����r#/-o
�Y ���_�>2،�x��,ڻzfqB?p��l12�ݞ�@��wm��b�q��m'�����Q1��{�B�x ���Nv~]Fh= Ss�?�6qo�����5�F��(�;El{�}D���ې>�]"A��P7`��=Nm
󥃈ÖC�]E< XI�� ��������]��Q,D1�%���3�?�Ĳ��!26�=��J�O�%��+݇��a�C��'@��i�m;0�������b.YW�"�Kޓ)o��V�(�Ú��(���)�c��N�S��[���U�.�� m��Y?G@a��Y'��%>��?CC�HgH"q'Ԍ�8q8� >��'�oQ� 
S�r��F�2զ�?�m�g
;���2�dy�3�\��V%ɜ�Ӈ�%�1� =�^ CL��W�v�-n�j��Cq�վ�AD���id50��I�:�v�������j�Z�"�]�?���O��hB�� ���uY���1��g2��.�^��#�/Coy��+tWl���d	�NS��D^�jA��Q��^��;���({G,3
qe N�����ӭ�5��G�T��2�|t��:=y�G-#���w���$�g�]��05�l:-@��*��R�jam��EN����~������8��-�����ͺ|��T���Ck9�<.����t,i��򎫠2�ppT@����u�G��.��FE@��g9��&KĵJ�=V��4ڜ�!8@��,Z�����+;<?�^���:珱�6�����^��R���J�5�*��.����-��E͋ 6�|sY���mt�b������E#?��Mj�h��yUV+�����Jk���@}�t�YÛ�+�
V�s�-���S�{yv�p��)�J�j�s\(�mA4"�s����;�i#��`ͫc���#�Ejus�	��]в��������;��/\=���D�-�9̴Л?'��\Y3z���s�L�] /�iVu���KU�F|>�j�p��d�
��l��~m�Ĕf�U?Qu=݉�u��nB�*!�3���66S#���*��+S7O!��xY�y6��O�0�L1]��*�(����c���R���]If��!ހ�	u���*���c���=�'���^�%����5��?�jU踎��QGL���?�O��E��0j����χ1Hŗ�ߥ�#-�x~����Snc+�c���}��Â��E0X�ڪ�Fr��j�`�,�ĥFX1h��x�p*'(aRޭ1�z�-4�0�����@ѡ�o>:zڸs�%�?y��Vez[�\�a���@\�׾J���Z�D��E�X�"-�=æ�1#\RMC���v0p�rv��H93Gw�8!���y��~�C���ʉլ�aS楝�*� ҄��c�����!��y�` +���Fz��$��K�.V�Jh�r��%V�@�c��X�!��>z���R�_7��}��+k
���3�.�{�;��=,vh�A4u@a1���6���x�		��+�k�I �H6X�й�����~59>���fWUg0����
��
��� �{��jS�p�?��u����sP��r
]��o�;�?�R�Z�v�?9�w��W���½uh�֐�<���s��U��a��z6�S�����,t��D}I�䙷ň����Z�6�۵����bŌ�<7 ���7t�:�&=��-@�����d����B�j��M>�"�D6j<Ӟ�^B�,�#[���]��`���VL�����^��ڜ0)z�\�a����&�Vi�
��8�sCHik���=}��� ����˔;k�N7P�r[����W�B-<a�Ew̧�1��i��&LVm����R�`;ʚ�6׾k0R�=�sR�\#�8�op,@��8�(i�����9"lվ3w�`�A�-��a\ �aGiGh�@� b9�B�l���/Puqe�g�������QRT_�xl���N\2 ���p8�_�;�5lB�Vl4�1{o�� �q��o͚4l���}�3�f�Թ|W"]Sw��u��/i�Q������@:p<MM�%,�a0@|���O|F�����Ρ{l��g��e���뒆��8s��z�_(f��@�H�+ß���Kօ�4�ّ�t>��N >�_�h�Ə�y����9��P@k�|K�[��f���I$B���BbT7��,S�y̤3-:�HaV���VB�2R�\�(
oR�#�O)�{��s�}�e��[���Z��H܏2��������~	�u>���$���A�>�8:g�����%���ژ��&����h��$W(�!��fJc���2QqA��c�~�[��Υ�L�/_�줍�5W=�/�b��vg]��ޔ:���5�Z��(�E*iN��/F@`_����W�� ����!�H��0^]���\vL�b���O/܎�*�ݑk���.O�/ZWCp˞��1[��-}_7�֑6����&r��e5�E�2�hn��������ϱXI��Bv�b^���xl��}|-�k��#��k!P���b�5w��(;S�`��(�;O�5�P��'&g����I6}D��㢋W)�J�N�@��~3?�r���oA=`�/�����ϩ,�8���G�� x?�0o��N(�b�i���龔	��^s���¸�DϹg�}�0��Y���O���^V 6��O�V�+7���I}�I�ٌ���j�r���3�86��ʻ}ۨ0����'�mv��#o>B���2��4����/�].a~�T��?��YR�9�)7���I�"3�H�)��C�W)|��G��ʄ����r�^��r-3�G�ܤ{z�hW�m)��ς�x�C8�\Y�1���ٳJ��6���g�qo7R��#
���b�+`B�Y2U��'*-Z)�����f;�P���΢�:��- ���u��E�����^S�W詇$O-)�ŉ"	���h���o�|
B%�;�'��"Wv*vR��>.ɑ�+���a3�f6��y)=,V����/ʤxRHޝ�L֜�����?�h�N��;$&��JH<>��:f�=�!3�~�V��Nhq����9�+�o]��R���'|&�ci�}�*�����Nc!0�4Ԍ�%��H<��r����$���E&����W�뎱���V��u�H(�����	3�{ޚ�B�w�2�KHȶe]UQ���<�A��6�BRH�B���#���%O�L���a�����m��i"�'��a�'x���=#���!s\��	/M퀚��Bs�.Њ&f�i0���ϰ�P��=�b[�g�v�Lo��7���^��JΫq�o��}i5F�����sy!_O�C�����3*?`z�wL�Tyȭ��9μ}�9a�*��X�}g,�}��*�yZ7��GT��Th0�>E�>0��_9#E�(	�;WF3S]$V'�������9a%$�M���oa�s��Df�z���F�9L�=������kQ��!���l�vS����,d�~���\������̀�`nd>I,�M,�w�%¼(��̾�]6��g���<�-���|#xf���ģ��u�QO�G��Y>���]������4qd�.Q�b���<&g��._���jgo��p%x�;z���������y�cx����i�2J[��d���{����� �P�F��x�Cw�L�^�O�f��M�A�f
A�$5z�x)KV����(?�`c��F@I��pjO��4�����0����	DX�WyD3�ۺ _�s�V��a��f/�~�A��p�%]z3;�������X�
�IH+��CF�Kg���|�ϳ���)8}��D?�\�	��������b9�(�J:��ZY���M�+�v�{�A�z��D���v�7��#[=�;���&	��ԣ�_Ua�GO(2�����','jF�S�_?%`�ڣ����ur�c�7��g��Y�������Y��S������I.A�"�4�I+"ު�t�h��SyP��
�cAt��Y#�^���j���_�#��),%#p6~%t���������&�]¾K�n�_E��|�ܖ����^��3�L���������Q�<ͻϺ-Ѷ�B��ir2��<�Z1yOD\pwlFS7�����\�S����/'�(�Xh ��0re9���1����v��������GT�?L����O	�*��/;�U=~�\\�$$̸�n"��p@��3�j�kW|�GOѫ�EY�@>���x�/�;
X�P^8y�u}�>$?�$d��A�^o�\��I�-0|9��ک}�SK$��/3�Q��ʑ�Yn��:٭��9�?ʿuܬ,�[�x��Q�'=w�=\�k;t��/;e�3�s�睦������*�6�|�̉h���م�a��z��
�{#j/R�~5��>�'M��!�΁�_��E���u�}�������֟�{�|┉�&��#z�����Qw��7��s�L��Q!xgG�y����zuu6R,���\������ؤKx���u�dȝ�|��LL瀃Y�T����b"��6O�̔~�1��wf���J��c�+�=>��e
�����ll��A��Ttv�~{
����>s,i(�z������ٛ#Z����Hl�N��Dk6G-�~AV��ڹ턙�S�Ŋ/��F�8��Za���h"�|�2A�ʣ`B�:��`\C�}��������  s���v�����#cU7�o�WOCW���ӥ��	�f������d��,��A���@���ߍ��a
 �_� ��'ԏ���26h�Ź��˲穹�P�G'���L�Tš�����U��.�G[�y�θEk���R��З���]Ce��#oĩoӆ*%����ܽ7���\橐����a�Kʅ�d8~7N�E8�)�=�s{'{�R1��@�	��^j��-/Xܾx�[��+�~�-ɞ��꥕x�Y7��R����B]�/4�"�K �t9@~���^A��6��k �#B���%���؇흆�/�h��)|�̟�\Ȧ���	
��)�J�/���	3ʃ}a�[P�y�!{0�q�!4�	|'�n�����YY+70��z'�1�p^3M���b ����0t�O�k^6�"`�;O���)VU֧{�V|�גJ$�
�Vxx����@ǽ�U��@r�
��m��5,��XC{ʩ��@*aQi`�0�Z*վ�~�Qw�I�9.k�s����������#���pΧd`+%�S��ϡ(n����K`	B��>���lϝD@4:�e�y��+���ui}eP��U�kz�E
YMW���p�}!�=�C~޿�t,�?9�i��>���.]����xUp��Ep{ڃ ��h�إs*:DI��*9�������ڬ6~)���D��,��(-���D�m��M���6!Ռ �|<^��|*/�<��M�
n]o���W�%[�mq �����ݢ:Z������2�K�]z)4$��	�?�~��
F�}��aDKuDw+��;�o���s���m���!`��H�pc�n���=.�dJ���kw��˳-��ۓ|X�`���up�r��Qc�d$����v�!,�����"���[�
I��ZǓۉ���U�+�0e�8O2�I[�?����g�ڳ���>�ZQI�D��4D\�\/���h�}WfK�ܿ{cK�?*�BnNi:v~�:$�e�E�~��A��oS��ws]��_�g���S�HG��.�p�Q�5������A�����K0`����Oa|��>uhl������#nT1�!|"��fl��K^I��K��.+*h�]�Էm_�HS�<6��$X%Є�f�s%���@�ǈ�BC[����Yg���t�'�qǡ��	�yb�8z���l�<>Xj^�ė��Ř�\�b�r�M����m��惴9��<b{�B[O�apu���^�{�ػwѩ{S�������nV����u��I|N�e1T�ƠC�	�i�t���5m�o��~L��RFp��N�P662pؤ�is��k�Ԃ��_f&�sk����5���������%�i*S�\�-�&~k�K2����Kn�N0�pA�S�t��w��^_@6z�s,�zK��`Q��,��-�f}a�B�<_EE:��!S�f+!rO.�<��ۖ��>t^f�%�RU�P �C�����'<4�d�^��d�����¹�PZ�on�5�XY�`�zlJϿ7p�z�E�XR+�
�hte)0�j����P]el+���bF�C¥����c���EK�����rs}��8��m㫚�[��aYN��c��/�;p���<�l4��@_�4И����\(Z��t
Y�K�-��ȃ��E:e��
T=�?��ڼ���G�UG��>;�Xc"�fU��E]�`�_��G�,ty���C���!Q�%��A��4����3i�"�]f\��%�!=*A:/�%��V*0PF�O��u�!+���L�V�h���Q��0�յ�9l�S��/ʷ��D�g鈳�	�R��mZ�3	Ε��`P��!@�n��vf~�cq��&��}p�������pE�5�$���(ē}̆��Vz�xY�	}ٲE0���2 ǡEV��S��L�/�����Y�a0�^���^�.�ǙE)�8��nG�X⚭���\�\2 �y-���)�3�P��4G�J��ǻ[DU��~p�\�\6⏷8��.�\Z��7�����ZCPԆ ���K����i	z���Q�0+2n� ��b>���JݲD:��A�
��d��t�9b㵆�4gt�oںS��j�I-�}��ttȷ�Xd�an�[�/�����%��_'����*�[�� t�,[6}�y" i�l�������)�m*���#�N+�C9�F�1q<���,���.n���-/s�K;�l`ѯb��Ͱi@M�����:R�X�YZY3oOl4�[��4��S��7��`��&���x��;_{�z�u�GX�9�1�4����^�-�����8��T�~42���!/ʞt����*Em�ZN(ӓ�I���=�Se�T4��SɩxeA�K�Є����/�M�$�>P?.�! Lp<���.z��'�-�z�i����.	Ѕ#d�˫���f%�g����w��1����#�S@� 70,�B�y���@����@~߁=�e[���%Ү�!��\�>��8�]OP<�����&��m��l��78�ݴ�R��R���'JׅO�����K���w��6Xf��Fnܨm�Z&mU� ބa��� �E�[��dY��Q�۵3�v#�I�`b��R\hMU20S�O����)�mKWO��O�������ն%EX�{e��M�z������'E@q������}�ݷ���Os\�2tn_Ff���.���?������f�_��e�0�q�{�2l>�!.��QQ��̙��UT%¥Uy.N,����/6�Y7�I:,1E4)Q5i^�zE�z*��:w2<��0�Ȯ�y\Q-��e06�q*���u4��t\f�A���=rE=p~���i�5���u�'xX�����eY��R�"��_j�J����0�|��H;��M�}�"}�F�9�r��	����2�����fgJ ����W�V��G��#��r��ή���
�q@ʁoB�^գRA�@(���pM��)�iUY��z���s�4Q�o���3߳�|&�~�t��0Dc0����hA��S����hcR�>"���q��kc�#�x5�NS�y����9���riL�4#�x�57�ET��Y>Ók�~�|�>3�e���
�)���l���G�@9��щ1�2F�,d��\���ߎd[s�e >�n�9�3�ߤZ�(�Y����3�����^!�5�x����N˺�>xI{�ATK�f�3��
���0k�?����U�#�~���`P��k�y3���jǝ^���W`m�n�|��o���a:������E�q\���-9_MS��gP��}_�%Q�XыC\p�$�E"Uu�m=��z��ɾ�����ħc!�~=k���t�ٱadJ�ϭ��fk�i��:ٗA$�Qy���}k�d��9�� f�	gB������_�m����l���U#d�s{XiO��_���b�go9[�,�)��Cn��Vt`�m_ mк�X�|>3��a�E��f	�2�p�Z9��w��0f���#+ �<��0=G�k8�rK����M���^�~�p��e�O�'���g�`�hɗFݯ����|���WE��Xnz�v�7�� ��j{�we5{Ӓ��28`C�@�#��D��U�pcR��l[�R�� Ģ��nZ5F����h��[��<��L	���������WT���Fa�n�W	Y��M��.e���5(���K��U�(�[��7����*����e6�����?�����{X����Y��*r�Ә�.~�=�E�5Vn����݁i e����F�5qĝ��0MQ���;`t�,$�p�/��Ɵvg�nv���v����E����8�t���� �O6_�D��8�f��z��H��Ѥ�	���3)�0J��.�����b��m�����
�}�$�I�AؔZ�b��,�al��|�x�d1U��ι0�I��`�M1!/�AP$� *�X[�-M,P�3�sv�wE����G�V;�C�d_R��>�T���;��g����Y}En����S[��wD%�Mw#��N%���9~?�54����?*��� 唷�_�ݳ�V�MFv�ً(<#���k��s�V�+=v�Mk�����yI��C^ws���@>�f��'}w�I��)�g �����rv��؁�#'�k���]c+G��{)�lG�Ksu��-9���"�.���L����L��$wg&�
�}��R9#�O��J��ۊ�\E_�ڼ���8�*NKm��N���?tq� ˭i9�~�y~ܱ�����BvpU�(�믋��`��?�c9���k�Q��
}����CpW��]�nIG;��W��M��F+&l��>� �#(Shjn��ˑ��ࡺ��&��Of��g��P{2nnO3�G������O�s�G65@E����'h���E%O��\ 7��h���}MY�V]e��fd��)j�O�آ��ݛ�{�n,֎���~�[Z��9M��- 3��jl	�aVR�^�N�μǁ�y��2�����I�K��4� ;ٻ���?PWb�AKbX����4����[�����Vb.2|�\Q�����(�8`ՔQ�^>��`�n�E�)�Esj(A�
f^к�y�4�&��E?R_�a5�%�E�ɿt���"<���-�Y0Ӌ�X��+^2�"�gL�q�)C�)��Bf����q4��]�CѦ����9�f��9�&��ƌD�@�2"!mR���F���{�Y��1��M�ھ�f�r�I\Wխ�D�?XM�=/c��B$�+=H����,�=����4"ҏӢ�i��;X:Ȗ��cj��;���6]։>�(Y��P@�����W~?yΉ��hx�T�~�Rm�ˁ?�c��Z��:�U��یD��b5K�dL[hJFw�y_(N}�Qf}*ijr}��;hH�C�l\/��'K��N|��\�2<��f9U�X����<�+����4�D�ZP���;�tZ|y�%X�"�恍=r�:�T�_������ W�ճ�e	+�H������{b	l��kF+��ء��z7:���������ب�)v�S�A�y�4CǦjHE����ҍ<�&�=��E?ss�v-q�i��/�
�SZ���1e�>���5�q������|Q�#Ű���5�| jCo �8&w>}Sg�_���&3Q�����g;��c^RF�~v��SǤ�--�:pX�)�eg�	F$�|�;�ɴ,^4��Ĝ��Y[����a�+���T�ᗚ�X�95�$�N��%�[`��N��kd�����I��I���"����;�Wy08|���������CChmk{�l0�A����$d�Y���t�<ٽ6��=�s�M�0�D�0�T�f-,�W��䞼+�^��JM��ΰ��7��uխo9ǋ��� ���3Hb�&%�hnr��u���F� Xl.�u���$�A덯�n��8)�_�N}�4q�5�{�-iG��[��i����ˉ��<sF�-������~ަ�$Q��C�O���U(��Qv	��:O�A;�f8�Ts2�1�Ei#�w-s9YD9&�;��KH�2w6N��}�b^[JTg/b��5� wa\��&�F��� r���z��	�^{�f��pij|�w�}E:���8��g����ћ�2"(`�a�?Fa��Iq�� V	��<~
��׀�C��`���W�nt�$nm����|��
T/�i�Wy�4Cy1�����P �}�߳H_l�M�n���sn-,�9{�9` ��LƏ,��P���|�����,�t���~�V�˲��@w7MGU��Q�_����w��A��\i�b�#�ݰtɓs�%�I����m�� Txf׈�����S�,H��f4\��nv�nu@��Ac��u����wG�/�mȎ�M
�O�^�~q�v��=�?��">��?�/_c>V~���2���;�bݥ6:�Ҕ+�� U�����]���&� �Oo����l9���)A�Ё�_������eէtcd�T0���X���QԹ�����ğ �ʮ	�N�b��u��)#u�H���7����?�#p�.������`��%���4��4�����-��� j���կoVy��a
���G.�8�~|]��ڎF�F��o;���`�	TJ���v��v:��P1����p�.�fa!RR�[�	$�Zq�����P��ֹ8/X���^�қ�4[�h��f6l饊����&�mF�z��KT����N�1SH���������L,��P�N����A|�C�5����`C����4�ȋ|qtdZ���Dԙ�O��O^��weU�K��m�3�7�9��������ÏQ�Pi���Ԇdڌ����y����9=m��v?R�z���9��6p�V���l����{�2_E�Uʚ�K��wR�'<��n���ǀGkE�W����T�z�ŝ(W�Hߒ-~Op��- �Jj�ZY�[m�_��H�l��}��X���_�n�ŉfh[Ql�|U�ZAp�=f��q���5O�އ@Cҟ'T���,yBq���I%���޸�J����X�[�.Yç(6�3�A�$EG[����D��c��n��8m���/���Ҧ���$�q&�K�ƒ�J&� �4����Gz�T
gՏ���hUw�L�մ�frqG�z�ooB�Jz9�!�r*�s3����
����
��>P!����}��h��=V^��BWM�]��U~R�>w1/�f���M��@��p1$M�ŝ�J=�����B�]Kf����ʒ�U��?~JO����ԯd!`�M��\��g�P��F���&n��|fG��8�(�r�O����s̅1��x
�k�2���m��_Aۻ#���W��ϳ��D�b���`��N�����U���#�-��u�J[���s�n�K�_zLM=sH��Oa��ZP^F�?@�\�~��:�#Y�gʲ�/��/�$"tW�/�*�����?�b&1Ǣ]�m��j��!̪�j-A��� �0��mp�w��<��]�	�\�� �t��Vb�:L���;w;�2�5��lMOs���e���O��)!T�����e
���r	�?( ?8�ԇ&�� 
��1����� ����CIV�����L�Y%�?�'�qKFo�
�r����SbK�I��q��,�-UݰV�T5�q��ᦟ��3 |�?�PW#�s��^�p�ʇ�m3 2�6A%���\�WC�O������	��Çh�8�w� �OC�%c��$b�:�,qZh3����� RW=��l�`�"�����ANq�/\�i�7�0��4q��v+I�Q��(�[z��u�������ZF��p��/����_r �Q�S�v]���J��C60XaK�u�0Nȇ)<�!l�����O�Nf,Y$Ay�9�w6(M��?e���w%'�|U5*F�����3�i�vTk�Poa/�o������t$1�^�<�=b;��;(ϗ����q�|���$\�-,�Y�b�9�pB��ƈ|p�����\�Nk�Z>|����������-�����h�O��ˏ:/� �'+K��b�U�x�t����Q�����D`��^Cp;?-���WE1�[�ge4�Ӓ!=,�9b�m�+4��D_��=ck�nbh24^���~��kS	�;S�λ5 �����#�_��أ�5��a����<��f,��VF<~��ge1��7m��^N66�z3+�A�H�{I[�X ��iF<{Rͯ�8:�[�<�������5��ke9�(�A1n
FH2��?S���B�J6ּP�/�2������i+��У�P����t`��fZK��M^�^��SM$OZ3�u����brߨ[Q"��6}5��Ag�c��'�;3m�\��ַ@#��)7O$#���`���I�#��
�I�>3>�Ũ��i?b@Vw�,C���@2��㹍��+��8���8� �r�O9�V�`�x�[F���!@�;M�1Y�y�/����5A���z{�r=�i�E����"E �>?`簈9�+��"Z�0J:r��5�F��Wx�J��Be�Jv�ܰ��p3����;0d�`��?�w8u	�'��}����4}����ҵ[�Y�7���N� �>kcn�Ё�-)`}�R]��l�m�����\�S	5jĝe�f�a�w�5Tؓ�ɸ�=C��
����V�u�swBn0����]����f��,<vVL�����h�x�uY����i�?c���[�\KmV4�>���RjpηG�N�)臝��3c갱v,��}[C\|X����#���[7��.���]��l�pzuv��d2< TJ��q��,���ŗkj39���8�g���-� (P�<nA���>���{��f��=�h	�?�a���v�t�5�[ ��d��o�?#�T����0A@�����G���� ��YO�\R����{K�)����b&���A5ծ���l"��ia��S�z�W��A��͓��0_���� ��&�ܫ��
�y7��sPX���l�w���%@���@1���Pn�i������,�"�1�fի�)�a�U�ҨH5�& �j�@ @�4-vh!��P�N�KF��z<,R��徎���W�MZ𯰱4>�`(do@_K�L�������Ƭ���"�z����M،Z��ט>$]o�gR�	de_$���ZYb_�Զ����M�����p�����Xز�lm',_>e�#v��k�W��9�\�:>84�����Ù��Y�,�S��.0�h�q���2���ॊ�j�x6X�SQ�����f#�*�|��E������:�('и�%������c�y���ކ{�G��mܿ#M��Q:>c��m�E�	uwz����4%+.`�Y�g�¢���Ϣ�����9����D��;R=.���⏇���B:E���)�ϔ� �ܶ��� 5`���0i/ �����NޒKƘ���*'���I(�\�l����&,Ҹ��~�K�,u�y�k�ԧ?��!����tA7��ë�|��U!��]�����'�Ì��P��84-q$1��z�)к*M^2�^4!�2\=�����J�9��ɾ!�o����yn���������rY 
���.�ߪ�y$���':]�U<h�{-�o��yy	�Az���0~���B̴8t�#Y�=H�=�O�X�\h��=��N�1q�@ʀ�~hF��twGy+׽�����p�J}�6�z+?h����v�Ӗ cf�����{��D�^�ݘH�_�e@տ�֣cI�Z�_zdC>�b��j���#�DP7����d�O����WcO@Vܨ2���pt�	꩟��C�S)�l^-�G%]�I�p���n�W��_z�DY����� v�F����@�����;a���JtE��� "�8�}�����x[Z.|��q6Ƹ�ʔ��J�B�- ����O$0'�T�m�x�TB�1L��խݴc8LbcM^}Lv����O��7�!���\dEB�����"�|��r�~Z���q�y;��e �殏�.�}��}��'-�]��Y>�(�.�H��ƣ�����hy�#�/5�����~2dϬ�,�He�;x��FVCv#H_��:Tn]Y�y��Uy�m;�� +�_����}�	F`�y{��W_�S{���6Jæ��2y�$4v�
I�4��B%���⽢
���]���K�n��P>�f:e3��K�[�W�?7v�� �$HN��˾&s>"t��n*�\��"4�G[$(3��<�a�|� ?�v�m��&cЦ{V�`�a����� �!X$ѽ�<��
�|YnS�!>��$*%�~�t��������}<Y� .1�Y<5ű4��ݐ���{�hm	���\@��-$Q4�0�]�e��5Ԣ�Pְ\��[1�j/�}�Ӽ8)���"30� �,;~��3PFt�>^��
A�_���)+Xр���պ�����6i�vq�E!����H���V^�9�ZlS�'
���V��2��Х��=y�14�֓UP^R�����+�D+>�u�l�ĥd�:�f��J!zЛ����@�E��BGC����X�j~�t�Sp��X�6�����Q���M�%�O7�R�m "�VJoc-�ugݾ,��8r�	���P�������	'K�7]%U k`>�a6��i�Ф�b�� �!��z�VZ5�����r�� ��u^"�*䇣��&>��Q��1jg�7�kR��[E�E�a���/9�E��wX�?���l�ւ����T��"�=�~�ۮ��>�id�|Tj��%���)v�?$ד�,>*A7j���ә T�ߔ:~/����!$�= #/�T�:̶Z�d������?�R�hC���d�#^G ь ��ь��ܟ���(�ɳ�@a�������s&`Le�-�_�Ψ�A،-�5�-��I	CWs���¯�3�Ha�WǐԵ�����j�������W^䃰���lstj��nD�[���5�c�����Y�?s��3�2A�dZN��/s�	��zO3:I�¡�"U�*���I�:aE��8�:���\�?]��M�L.�$�.�?����|��}�w���Y�k����Y\�	��1������`�y$Z�L�!��4.��9q_̝�Y���U��e�� �L~,�M/C`¶\)[1�.��Y��BJ��n�x>�/�����I^~���>zπHy�!w���Ϳ
6b+]z�5��j{)$�9��8S~�:����1nOi�w���yDg�"��3���y�s�ݴ8��[y�{`}��m�\�ޕ��S��6�]�,�v��-ك�_qY^�L��=�a���5ꊯ�J␜u��S���jV[��bc��1�Y�x<v��e9���{��:I�ݢ1�2Q��Ӏe�$hߚ�E2�/ζ7[6���W��=�ь�p1%��Z\_d̪ƻ�2� 1�|ա]8���'lv�������Y�sؖq��
�a�����# 6��E�螵��`q�h�jD����ߌ3.ޝ�� ���?�1���*�Dp����\I�-D/�.K-����_���*֙���+E+V�2��Yw&-���;�J�/�ě�*�	�g�x�䭹����<X�_����J����י�p�/�Q�s�;�_��)7Eb���OQj����)e�z�uZ�3SM���B���Y7�_�_t�儚�II�V5Ɯ\}�cmO*���;�<�����1d&ctq}J�?'$�`�Pyp�\��^���c����� ���$�n��Re�������"GOeO����2k�ሎ��rm�h�y�� ��>Y��T
U�A:��8Gt���&1�����Tl�����@�S_%5���A�"�n'�e��d
��+X-#WIPx�Ec���i��~�D1����@h�����b3�v%�59����Z\`0�ZG���\��&=��rT�[�֐�p�iQ*��!ô��Qg;K�a��\�/����H�=����ߝ��"ǐ�~�9�nw!����
a��D�~�rNgl�*+韫�>�D���jF^G؃� 㖋1G�"��3���|�ɣڞ��C��!�J��S���P�gB �'��g9}�v'|I�|ڪ\ޖ/��;Llu�47vbh^`.�
�/�k=�tΗ�?�E{�i�@�s����[�X�=��w�_vD�h�Kj��-���:9��v��P��~b�H������?�z#�����20�[�V~D��r?��{��;|���UH�$�`�%}H�O�m��1JP��l;�~�0����V�uע���i���xanZ���z���&��E��pj�×L��vj�@�˚�hn��j{c�f��+� tk�WS1'�����!Ѳ�z�T�b���%����<B8i}�5��G��\�<sn]�lX���MʵE7~[��|͉�ôNGʩ�ST��hdR�,�7x��i� 2�2p\�8��(Ф�&�o��5MΚ�Ҙ��Q�`ӾX�ִ˽��C�iQ����Hk������{��2�o���9��^ow�ҠH��)Y�
�ce�
[Rl��U�V\���Y���O[���j��ڙ����:��_F.����G$Z� v���� ��W�Q֤�D����)>���!n�|�C�s��'.�;d�4-䣃
��}"�<c��8C�57��ƣ�U��E��S� �Z�ݔe�~{��0�LM�˨��wd�ao�S�0����έ�N���,�S�"�΁'��	�w ��*J��=cƪ��R��	�pKm&Ф�O���ke�_����fJ�yLZL��O�WEN��]r���k���gw˱? �j1Y#�d�6�B�\h�0��9�B���>|�+�u��T��Q�N��S	q>����bJSb݄m��n?�΂@�7^�S����LxZ�[[�T�L˴N�U@9��c�o���q���L�A	a!�h��Y��U��vL�`H]�x�w/�d��/ռ���,󎈕�~�̲�+�J�XИ�ߓյl�?ڌQ�:�Qa]+lg﬿%ȃ-�����
���
o�c}"�H}L��p6���9̝x�Xr,��I=CX2�P�/�h� ���FA��I��)��9�<p��0�+�[J� ��|�q��ł�f����"����5��NS[����h�۽�q�^?��x��q?r���?������$\�'�NG>��iȇJ�Ąh��#n���������G���;�qw��(y�b*�8�;%i�2�소�)�U����T��f��'��}@�R� v��j֟����l!!+?�0����ӿ�}��fE�&a�\"�T���W�5|
�d��ѻ%6�Ш
_:�s�ۘ)�L!v� #�(� G���s����?�o����F5�2+W��IF3�EXm�o{G�=�w'�aT��]X 7��Z�tB	J�(��ΐ�5��P)�Rޯ�^"��$*�����iM7D�V���g��r*�r��+��q��샙;+<m\֏	���8����� �t5�A�Ĝ�����܅���� ��6��{a*tz��w�,Q'q��h���3�N����z�X�o~�px�ß�ӧ������:"`.i6d8VC��{C�#�[L'��b�s�-�˓��5���y�[x�=*��n��ȉզ$� I�ۛ�{�,lh�k�z��I�:(��֣�*����.�(S�|r2{H�7@<mi(V}�	<e�N:�!�$v�������>H�*-�u���~�GgJ��\j�`��Z�є[/�$�aj���A���Cf���Z=AdX�U�&�����O����8v�'�~!�To�]j7�l�:z��O�[�=~"65wa��F\�w�\����q���vw ��DѺ��֏'�5MK>S�zZ��X%��Q������������R{L�MV�����B��Ţ�K�GON�T�8���]�]{���5�k�^����g׻���Ps���A�W!�;������)������>�z%C��*�5��6�m�4�Gu� �x>�Ё�߬H�����2Lx�)�%W�d���ƨ��{�;;�����":x��Y�s��!�+ W<0� ��f�a�|ٶ��i{g�x�~v�}���U�n�ֵ��\�hF���sj�L/��*2��a���%��jQ|jC��Ju�<�,�9'���¢�9( '��_Me��.�zd�N7���lP/���S!�A)?$Rf�1���������0wcF�	�|h�:�f-���j�S,�e%�k������i��}�V�2��ń�қ�GY����B֋�R���q4��y,%�:��x�=iѳ$*k�WC���w^y�$�y�M�)��j�����q��W��mu�����<X=���0��:q�k#&�^���HI��qY&~YF�Q����4�i����F��&Z���07�f������9��h���}~���v���<�g��r7}p\���O��_��J��%�7�� <l��a#c�F���74�2+hqN������gk`��@�m����+�Å�Pb�V˰x�U1xYɷ�xLk���~�k�M��p�bgS�{*1W��'3�.����];2�B��S! ��f�xCaQ�����V�ͩ�8G�����>�I;�;25r#�\zM�^#v|o��@x/��L�2Ϙ����ۭ�=���eo�^�"�k����\�D�zir�������Grwh8�NI�X�!U��X�'lO�5f�o*UJ�u�huke SR���K�.�4���#}$���]=�X��ܻy-�؋�id,�\`�> ���6L�a7���1�D3�1s�a[ދ�|k�.�D�Ǔ�i#�I�ݩO��7q�L*2���N{���Q*�*N��W�H��ZX�R
Cc�?ߝ#��<�Y�@��	�,�1X�	��hA@���6g��;���q��������}(�n�r0�a嬷E�+QRU&�!F�m���|�Q4($g�W�#j�ߋ�Vq�V����pӝ0��X�����t��<�0�����s�+���� ��@�IsBz%�a�L$,�=!B>��J��O(�_M���L�*�7@���;��w>T�{�J�}�$ah.6k��k�D���k�|ZΦ�'Ӻ���}ӛ^�@"����#�Jjv;(C	�T���}�M���WD~;�#3��~�_9LCh3'��������/�����P�%��t��e��/~����s?��X��5�q�[�9�Q���I�å���`�Lb�~c^�£��U��BB����ز��ן���	α���']E��xH��f�׃�	@S��\
��������i��d�Xɥ\�����e��|�)w�{^%M$ f�Ţt��nc!��5���Ȯ�b,BO��=������(��č�
�� Ɣ�YP�f�c� �buP�!�T��
1?�=4����B��WB�C�*�}ӒΧ�tp/���~vH_��g¶����:wz�Ó�^<���p0���n�g��,S���[d�g�G_�{O�Q��@p�H�_�)k� {'h�*j��P��boú�|_�ccÛ*��N�	�-vɍ�^T;D�I���5����XY�<! jgУʦj�-�4�7�9��Ms6�=P�S���
��У<c0	V<�I!�q�)�|�����9�
��]Ή�v�EFS��`�L�K9-�0���M�u�,${��aE2|W�[���a���:�g��v�����0��T�zZf�^��X{ s��j���&�i���6�Z���^HB�M�|:,�	�}a�U?��i�h�S�B93!/�w�k>�9�^H"��+E�A�{��4�Ms���R�j���l]�T�
E�9NH�N��l�zk�D�	ܽ��L�s>�T��ST�5baz�N{�AAכŅ�&��?!gN�:k��|�y���L)���۶tG�O�ʯ�e�����?ϯ��U��=I���cI�>-�Ƃ�!��-JU��R�j���5<�M9�>�M�?
5���kڡ$8�B��>�uo�{wI�uw����b,#�o�F{A��4��T��(�>QZBv"f�e�N1#?Ya�O}���k�x98��b�p�gD�.`���P~�UdԜ��!F>�h_�!`��v��X�j�>��Λ�i�!��l��QG�$ڷx�׺NB����]l�H6���*����W�%�A��[��{GDi�%�?�Y��8������ڜ����v�c8�"2ߐ�,�)R�c�L6J�=PW����s�[X��
��)�/�l��+"��t_���7�ʅ��ə��3|on��Pp�3����c��'S�y02��'��5i��lI,E�[���!��hOC���}oV�^żE]��\��+��EH���w�ݻ J�Oِ���t?��Fu��N�}�ܭ����A�1UuRZ��`J����^������pj���$2��A Daldg}o��!����DI���*�ݱ�A��0L��<�w*C��%Wd�Wj)w���@Ь;�y��yh#S@B@�*�KX A�:A���`v��w�hen��旅g;r
#7�'��0/�צ	�D��a�p�so�ͧ>�h���]KGW�Īi��4��Y��X�<�i�[J��*j�+�ft�B��wz2�~�K�ڭ:���?���:q@b����׈	x)�+�_�j�`��t�}io}Gy)���:߱L��Hyż��"7U(��Lx�n�w`�[=�q�?�XH��)Z32
����9;���b�44%�1(��#��:Z��o|UF5���z{��R.l���7	wmc�k�7��(��}��C��$�J.�,?�����g��5������9��e��ݎ�����N�����>%�	�0�q���NZ����<e���6�uM��i���Xjiԙ9���������vy]!$0j���;�{K�=��`�X��:,�Vh�/�M������¤�\�"T�.���U�;LEǮ��|�d��$I!Zd4��*��zxWvJj�D@Ey��ﺖ*]�Mb��P&�G'NB���ޢ8k�zfz�l�B��I��Ow���	�YP����5#�4_W9��b�Tm2I�_��(��8}��"hoD(�]��.�_�3��E�Џ�:���P*�1����e��XD�r��x��m��-�DT�ai��^��&|�0�NA-lA��YbZO�m.���Oj\a?\�2��oM'~�R�`6Rx�k �"^˲[/Y�X�ʊ��* �˚�^���qr����uN��Ɂ�(I��R?"�I|� ˈjVY���s�5�b�Vc�0�����E�YTT����]���V��i�/Q3�^��A��X���^�t��_ ����]R�"�[d�;nNM} 4�S��m_�Y����MWv�i�6j�(�6��LB6u8�X�H�L.�aV��ĸ.ӍC��~�HX�abs
�U��!�y���V�N��7;֩_����Y��Ń�5�@�F�Ӏ:3
c��`!������ӯ)�+ X\�At��7���ߙ~�����}B$O8i�Bp
�Pӳ"�E�u��@u5�g�;̬��R��g�b����+�'���3Xl=\�����g��)r��CR<����Qރ���e������#�M�Ւ�K3�ξ��;�F�o���r��9�;Zi6�p}ڇ����ų�A@N��D����|ɖMw	+�IR�ƭ�A�PK��{e�$gYfS�����NP�W���N�5@�I_�O����PC��|�����!���S�M�~]L6�ʳZ(��	��˛��q��y�L�ZͰ���I��	�Ȕꀭ	{D�9�d�P��r��]ο3)�|b[�����nT���"�X!v��Xx�(���"ȴ���LZ�"'�Z�����,'�<����/rBsJ�dx(H^�$�l!��j�����#�	<33_���A?p��;G'tEQ���� �6O^YO���_���H%��1�(����_&��]����A�������Ii�@�D��TÔ�琂�2"zuh�'��b�U�n�^F&��O��y�w��
��G*���_�Tx�)�z����#u]?±#��-o����C#.f����K�~�. ����qkEB$9C��T<�p�#��)��1\0!u8Qo̔Jf�u��SMZ�ӿr�ʂa��ӫ���7�:^?=aWB���B.Y=SU_�GK�d|:�gU���b�rǥ[�\ ����������Α:�̏�G�Ưs�0K9�Ğ�/Wt���1<L�Jn�=�������4^���U�z�pt.������x��B�p��"��oM�*��
���R���Il_� <ZM��C{s����j��N���X>omy�^�!�	9z���r7�8��dk���C�>OR�p7���J_�����"����mE<
��^=k��0�\�h#�����On�{˞$ 3�(�`UfB��p�����kP�I/���I�3�b��#n�2��>_�[�e��֖�ZF���5!��{O����V]�Z��,�8�(!N[9��O��j]J��Z���E�
����l��[HC0�J����[f����NO��~�~�CY�W����4'\۲�r���EHP*Vf��D`��a��Lr�
�i�[�)�M��7�ډ����;�>w	�6��S�^A��������t`���|��@ǵ0�F���F���,O�mė.��|�h,�`X��|{�a�+�~�a��T����qDE���R���.���t�������M�^�j��8�prU�U���H��"���	�����r����0P|�"��g�@����D����>p.�Z+ߕ7�Z�L��l��z]����
#���j�,�+�A�A�90���8V�j �t���s7��-ʜaI7�p	�8@�1�M6��ob�
p:�����hP��R��c#;���U���,*>���<�s$ՈmyU)o:*`�m�6��l{�LS����Q�W�����=r�c?k!s	�0́l�J���C���ڬ�<\�0p�LO�v�͎9t�)3�Y\��(��"c�0��{T���
�\9���mB4�����Ҿ�geo,cbG>�NDLN��X�5�r�V@�<O���?Yկ��>8�Gt1�^��9������w��w'�$���v-�Y}�qː�� o/��݇����nP�����a��Գ���Õj̋xi�[��e@�,�z$��|�k��L���&.jw{�j�Ҁ�sl��|V&��� � #�V��@m���h�Y ��|����MS�'�`��7�ȁ���f�%��C�:Z�<��ҹlcpρ��L�~&&�]�3G�*�I!�Dl�z[�it�ӣ�!���"a���Ć���n�aU0��j��MD,G�֢�L+��Qk/����������6�7�Vs4��x���������i��$F�Z�a7F�.@u=��}c�N(�9��6Ю<aBD�`�̹�K�`q1UX���򯰽�C�^iأ<�!�J�wBO�J�BA�Ra�;��/I��!ا�h/*^*���� <����6�1��W�qbXoB�,	�F; ���*�NM����m��&�P�؀·U���i�&S�u]�ݪD�/�2��`_pE�z3N(��h4�.��'v���X�*9�9�D+@)��)++�!�H7�i0�]<�̈́�!���Q��_�R:��@r9M`��9�z����a(�|Qog�s"�r�F�6&��\#�ʈ��GB�F3���Q7]u��z�`<f0Z�<�+�l�e��o�w�q��`��4�d�/H&)��S>�p��)�fF2N
o2"�ń�j�s�n�>��������_8es�L����%Q葇%)pm���<(���8n ʊe���R���/��c+oZ�������a�ʎQj���إÙ9Y�Ρ��������Pz���]��,#3�`�o���Mj��nn!�5X��C[��i�!�с�����&i�2VL�V�	�]IU�:dg�����)�$`����p��@7�u�}�1G-G$&	�tG�<�I�æ�Ν��B��V�kP�ve,�ky67bVcAJ�|B"�ℝHT�dS�h_�*6��Y��B�������~3����;<VfS\+�r8�����-]0����%���s3^f)���_V2W��h��Y0&�/��
���%�夎��E�?�Sw+�M�
W�}|"\ ���&տ��*mT�A��`��D�0O��lߺ�|;�X�[��1�0����^��u�K�������)���y҈�Q����� ���q�� p�Y^��B���Î�מ�f�ˑ�ŻA�'1쁐�=S��5�ˬ���'���ʠވx)��ɐ(+^O�F�W�M��L$5	���6�=�2�\�����r�4�� 2$���[���@��AVy�u��dJ�ݾ�G
7�wp
%����B��3��#�����`^�K)�bH�V����OrL<d?��,�
C�/$h��͒5�,By'n��
O�m�T�K��u'�n  `�`�Ǩ�����8�Rd��bj�Vp��δ�+&����\4��M�Jyw�В;�[�Q鳮:���<��[�Ұ�/���S��N.��<=� �`t4�otJk3��f��ǰ�q;���%��<O�|���wS�7.��b�����6"A���%>�W:��!�)K��s��N�zdDu2�f�H�$�EA�%s1 t&��I����O��t��-������}���#���UH�-���&�s ����C��-����ę��?;�n��
J�22A� [r�CE�XAA������W��"U!�_�ܦ$WB�@w�����".���pn�s��s�-���2�k���|`�C�:=������!|�A�ϔ�F��(�����u��=�.�}Uې��͞��/OՁ�����e��B\����6�I��CT�#.�ؒ׷M�l�s�LOv�ʮL;�B$ݞ �4����vf�E�\@�����p �~$`�x�v6a�!jF	X�7��O��I1��}(8Zp+k*�;Z�e��9�=P��tVG�Ly�b/$��Sq�p�v���n��&������8O}s�=��ѝt�@Ȼz�)�v���O��}*�|*@�]�>�B.�mpid�dF��n��ƻ�w4��iQwZ ������2y��L�o�!���.<�OH���	T��j��X��o���2�{U~���M{�)�R�@��f�;X�Ȱ��87����J���K!��礋�8W�Bq�
����j��:�L�?hLȋ��L��"д�	��p6��Ҕԅ	���io(e���h�I�6����f��y�������pu�J�Qy�k�SH9�y���۶:�B���Е,C�n4O�;��k��-�/�?h׀�q�^Eb���4���F��ӗ3�H�����ۊ��~��S@mوH� BU6�"ӹ�L�2�M�b*�M�L��:�H5N�G��h�	~D�_q��2B�F�RU��z:��i�ƹ2��#�6k����������DF�.4v\�*�Dǲ�#�-�O�-�r,�o��0h���N��������wه=�ş��n���F����_���(�4�To����",y�!u���=��=�;���qܑN���7>�d���?�%��10d|������@^�٩'D#2R�=�)��E4��ǖ��--�U��]T����p ��CO� -i���'��}+✇u·kE�W���L��S�Δ� �Dm�f�C������� ���̧��x&��u�$8	�o#� $���$���˖�H�r�����9�2�1�����} t ����g���K�X�^�f����О  �q����l �t]"P�J��W�*A|�w�����a=��W*�JZdlzq�Q�E���nWz�0	�,��#����n?�U�W�a�A!;�/G�r*����F��Ѵ����_�*Ne�	Mw�P��;�z�������m�P|@�����)��UJ���i"�BRY��]m�Ƅ��-<Ár�����msH]��٠�|���2*U���0�9E����U�+(��5F�q� ��M���́���iM\�:G�R��_PvE������!�O��"�7����d���ݩX靹n:X�a°���IjVZ��Y����՘����H4}|6+�ZT$\=�+<w��Lq��Z�#X|d�3�_w#�@;Ig���8�A*#��<~���`@�q��W�C(�˘{���c1�l�v��|�&8����Su���V�����f9�W�[����)�giټ���j��X��-!k���U��8�犵�Fa�i]op\���\6�&7�gó��PJ�${'G�L�É���N���nX3)����
������/���a�w���D,��Q��N?�4����xS�7� y�G/gR��q��|F��Y&.+MͨT��>Z#�n�ѯ���Kj���ڔ*p�����'�jU>繤�3,�Q�ڰ?#ڣ���Ӄ�gI�����z/~��ي-84`c=aۧD��QrYU��N���%�we��٬��dBx�/�.q2��d|'th�.�/�$���ׯVώ�aI 1�Vs��~�e 	�%Ev�+.	\qwVyM����t�,��� !_>S���\_���ANt��&ψ�T*c��O�2�`T6�
d�j4]}~(�Ҭ�5���1"ksZ4s{ �
��3r�YǮ��BQ���:�R�mj^�V�0��f�9�aYH�^�Ȉ!��h��ݠ4��3����*D��Q��	~��@�W��O��p7�m�S�~E� ���7;���0�K�_�Ɲ�kI��BD�Wt)�˰��`>ڦGj�T���fB���:R��b�����AC�(%i��yr|j��_�^���k+�2���t��e����wų�>��d�\��N��(�rIb�iF4pS֯k��L�Bc��j�;����w��(���}ѕ�k)�^���x�0���n�# 	�{.��ZJW����}��������M�^+o%v�N����##���B����w��+����mŐ�� ��>xY��S�z5��$�'ۘ'T�uظ7��H�$����r�}��n�}����y��hO�N~;s��	�p�c��ģ�6��e�S�����#�_�<ka۩�]��8�qv���̙�^�Z�u{�_�6��R��>��U�b�u�����R��^�sxOv K]�cw�7>5�Su�C��A)g'�`�q��73T��h��3�G5�T���c�3��#�W6m��z��؋�w�Y�4�w�'V@�cR����52U�`��2m��G+�0�9.�(��u���|�Z�!4{�*���3v�rO�O�Z�Ll��<r��i-X�������a�X���h�2�d�i>a�2pzA�<~A-)J�Bl�(�x�b��g�aM����Aq��>������f��<!'�7��D�Q�8��:y�2�#/�v;�c�h=��yT��8��D̗�@��᫮o�"�����"%8q=U�ϖ9��JЉ�
��oҁ�*���n �K�)��VFV"GsXCg�4�!U?��dY!�_���p7hsw�2�$�s�^`�nR/bm_�o��2��g���g0��f{�4
c	�k�j�>����o���:е:U�����H���߂D�yd��U��`7к0�ʍ�� �-��QV��z1�
�7�ע�pV7 T]\@���q9�i�Ɗ���GT�z{,�58�-���>����렶 t`�D&Ʒ��t�Z�xl�vz�LC���39hn���Iwn����x>_7I��WlHL��J4_~�y�8�=��X޻�e�D���H�jAj9�H�?�L�:��~m�u�/�-tޔY87)���h:��D]��䫨s�k>�54���ц��&E���L�"���$L.�P���Q7Z��_5o��$e��eL�H蚷ކ�m88 K�'���Ѿ+"��7B�& w��7F��2�0�x1;ة���2Fw%��f�`h b��P��*���gWh�g�u��䮎3��uc���vI= �e�:��nu��5K�f�u�O\�]�Ҍ���[��=��w#�v�(���,,��׸13K/�OtW	c1�,�;���aSa��*w��O�����s+^%��#�{+ua2�v2�R�D���u�'�~��g��k�+r�&Umr�E;�����z�'\��.�t������LF�Y���2#
�_�O���Z��/t/�)ˠ3�{-�3Rf��7���>T�:��aa@϶DN�4L��c�s^�i0�W^��x�?�r�)��R+���[�Bpkc0��0:�,���'�[�⽜�z6F�>�3̺�=���R:gA*�g��ﾸk��#ހ�����2���(:v��h�%�4��M�����4�kf���5̶w�
�#[;�%c&5E�g�s-q�D��GyL]�Saf_�����
8��g$�*S�2�OKi����3Fwq��3���1�nar-������� �B����S���n)=?a^b�b3�M�20㢜#�.��=��s��y�3��hE��Jˁ��x�ȅ��&� ^������p�����Sm� �����:)�6��;X9Ors�����PV�@�8��1��Ǩ�acSZ����4����W�
lf��n���4/Ii��4۞�1H��4�#1��>J[E���ʷlU�5����U�7)&}W8f���_�N
���3�*���sU�3���u�s%E�o#��j��耜�Ng�l���9���Lg�W����n?��!������6�RqS,�!�^�9�/QX�0$�^KpF�ڷ1��|�1Wz�`�7���L�6�
��Jq:��	�2�� Z��;K� ^1��-��?ɔl=����F�>�_��\�Ԯ�3�����xR�c
���GK���!�u�Pu���QLB�5�Hq��S�^��3�J�Ո�X���(��PAE�b�>�ƽ�f0(�V��6=_��'|�cE7պ�J�`�Qn]:o�q	_X>Wڱ�f�:d��}������9>�~���G<0��}`	 �@YP��"���
���}�����)�C���!���9�1P���K��U�6�)�;���wTù~(�e�"�T<ދ���(6,�-��w"���X���h�hvT�1��փ�,,61��{��'d�jh�SP��|�cQ���,���/�i�<8�mUQpJ�_�ā��l����h�,�6��=��7ĪxJ�ԗHIϐ�`=�N��(PʿG0���al=��Qh����Û��!�e>G����R�ǐ�����;Z��&�I#��;��R��5ztː{�!�^�5��O#��BQ\��[����`�@��@	2�>I="H��	Y.Ҁ��q#`�O ��wkp��6y{~��v��|L��;�ͨ��*T�A��~�;�³��/�D����Tg���Q��[������4Z+��r"c( �D<[�ּii��m�P��	�,<��Jz㓧��\�s%*��ñ+���~�*���{x���h��y��"w{zk\9|5��.M^6D�6����3���ꊛ�Itg���[19R>�W��x�|��r�'�(�io�r �-�=M����|�9HlD�����6�� �ڸ��g- 	Y���\��Rx��4t�m�7}c �0��A�#�9���='꽉��Ǉ��B�,���5���'k!�ǚ��H��j���
.f�ڊ��rF>��u��#8���'��;�Xz�����w;?�a�l)n��+�� ��o����R5*)_�J
��E�'�7n�)�����
s��
r��7�0-�`9��ϐ����?<��j:J4N�Y�B:�����N"��(Z�4���+�W�;� yF�J�1/]���4j��yiC1S'_�at�������$ �{�~N�W�L�wm���Sĝ_�~�Y�J����aRb��t)���(�+��5���ˊ�~�`3%� �`��Z��Գ�Y�(0���,�ۗR��%M��;j�σ7d�y���}�џ�4��-Ҏ�l~q>*��	���lw���� y8�ÿ����f��M %�ʋ�2�`�O�R��F��ޜ�2w�4�"�|��Mߝ?(�����ty�w����$����',qD�[�y��5E��ql�:^���~�:����=�@KR��V�M�ҙ�:Ke;"#A��˵���.)y4�����֍� q�����k����skT�l��[�����>�V�T�R"Z>�{G�]_=b�M*�c��MRݶ85C��﷪a�ڗz!�J}��p��#9^���xl�t"��0dPK���H��ɔ� Mf@)��2h�cc��!y7�i�4a,L"+�g
�}��r���H{�b��q���D`�;�.�T���C��B?�@{�`��C���L�Xx�z`��^���G;���AR��~t�nLJ��b��x�l
Q~�Ԋ����W~¶��+��y���P�E�5�9�Pe�p� �M,nXB`�V�RP��*j{�ѫ���((oE��/%��)����ʩ`�#͸�A"��B3���k����ۺ7��t��J�������@��`vaT���  w���S���Z~�`��@^ā�=�_��0D"$�-�<b.�2Q�O�|���x�Z^GV`�̰���Δ�����fdŌВ�el�=��a�h����?� �h<�=`����5�ܒi=e�&
�d��^��� 7i}�ࡺ�!���Ϝ�I��<�^ �Z�%+6<y lҺx��0a
�hG�g���g�蠴��M��RS���Wΰl���k�H��y߀I姈�۷���Uhi<�4A4|6��`Pv���p��uQm��c� ��嚑�hH�v�,3���e�l��m��Vr��2[�j�����0Z��10I���?F���R[�����Q�Q�Ko�+��BՑ���3�o�"#Db G6�a[����s�?a�0e�Ua�d��!��@t�݃�ő9Y��d%�)�{�� ����|�D���<�.�av�Y�)Hs��<�$�Y����e>�t��O��@�����YT��d�Ӂ�N��l�A�hRyÁr�e����.���:��Wp�)�y��wIG�~4;L^��;��H3��
��b��Fqy�H1S��/��4��(����v��y2:��J ���ifTPE�5��Whk9lT�b���*ˊ�RQAhN�3�b0({-y#͢ǺIB����f���bT��V~D�,X��ԪҘ��lK��|Ȗ����@��sW)�_Y�	�2ь/GDb�8�րX��q�"���*˂pkI�l���&�i��$�ڕ��*��-�"̦��U'v\�r�3��oX���g�	�6Cvm �t\�̚����*�)���V��˥���O��x���i������/b�e���<ȕ�����H�Sͪ���afX�hJ�!jDm6I�k�bs�x�h��㖙�{�u�n0�/c&�K@��IdӇDl�M��7�Bl��
E�̺���8B5_Q;R'Fi�.��[�|K�����Ã�t����xH�r6��������
��q�j�/I�C�+�X�^�&M6��Q�>��Ŷ!sh�yAT���[��3�_ s.�"L3�C�qX������/��lɳ��Tk��xf�\�Q���Qo��� �sN�%��e-ލ����X�}|��/C����I�4�8���B�z�r'_>S��Ղ�
�5�lC�Q7q}���`z��7�?�`�"�>�X�7-�2V[S��ey4��Ѫ� Z�(ھ�=�K��Z��Kv�n+�ѵ��J0�p��w�<TZ�\��X��"��)��sO�W�׉���&��ѽc���AaI9	Y�t�q��P�,.C�}}%�Pb7b�C�Q�����O֌�9�b��X���l��2���Nz��Q�p���#��v�<s���M�oP27����P���~�J�f9o�������L>*�F����Np�D)��Z59ܰOG3��9ͬ(���^>٭p:]������6)u�_/�Ϥ����_e��'�)	&Y�h@�W��Ĺ��$�Q���k�y��E�i��ņ��j(9f�t)C�h��m���sQ����8M恮I�;�������z�7&�5���6u`q�E�7�!�۾Q�s��>�iM�Gp�(��5�O�WU�:~����/e����-����P�Pi�
�(zT���O�����R��S�22o8$цj�}���sB���E�:����A�,ԣ��͊���>��r�u���cIT����h]�%��0��䪰QFq�mjCD�ٷ#��2R
.�+7�ݱ��d7Ht=�U1��
�/��sDy(f��Ī�ž*�)�5ծ�f�!�UN�F������5�1h*f.hF�_L0-�VS��/���}lP�b&��i����U̈�Y�A��)Rm��.�qYu��4
���u��u�S�E�#�Xտ'�2?0]�}��9:�/~�I����#w��'�Gf���eD��©Y���gq�5*��l������m�J�vɑ����9��p� �i.�H�Wb8�I��
n��@�,�C�E%Ri��ܝ�bl}Ί��y�%��V�V��]�d6f���F@=EŻ1�K������»ژS��/1��a0�V�q�{��o�|�cll�d"u����~A(Hrh��O��Ƀ9J�B��e5��XQ���_�!�!����oR{s�,���V�F6l�.���r���9�e�Fi�B�\}܍C�$���N	�Y�����6�o��zB���Ppā�Tv�đs^)z�M�����ܕ1����c�Sx��a!+|&��]��G�L�#��^��c��k��J� �z��|ث��xƢu��*���}�C�{eFtǲr�XYJ��'�Y�튉e���}4S��nqò�K�wT�:��P"��R�>˕��֦� ����;G!N�ޓ�#)�=�M���iӿ�E+>q�8���g�
X������_����-��	T~H�_&�����tA7�$0��1ąBD���_҂����=��&Q�δ�{���8"�+����(���
��3�2��	��<�u��߇��_��Sps�=�brf��x�����M@�q"?+N(�Zp��<[R��A��Z)U�=P���a^���U��xD���4y�"<m���ac�i����S�aƀ�Y"ƻ%݋���:�L$i����6��'QTZ�b�5��9�V
��ח���!�����o�( ��z�^ʋ�������.eA�A��8z�\�[N��2�G荔[�^b�mK��N�`�L�Dz~	�x����E�ot�h�Z�6ur+�(Q�?������Yؽ�#p��� ������S���*�����L]�\�_q/�D}(N��;�V��,n|���w�HUT�m7~"g}������0�����B���z`K͞!7����N�-��ǂ��sfU 6�ѭ�=���n�U��3h�bΔr�B�϶;�NX�`#��K"
R���|�s�N�"���l��7K�n�i�:]gD� 	�QB�\�8��?��u;bդJ�ր���K��9g4��yYA���a�ο��P������v�1�x����������m{ ��B9=��gU��s������zwU��X�9�.��a��j�����B��o���Gem7�3�[y�yѕLU;�-��K�d�Bd�2�Fq��%c��Ep!`�9d.W��c�M���Т�!�-���#�&'�I��Q�k����\�~/a9��e��4�`�?^f�T�<i���}�8a]�V�Ky�&9]b�8u�_VRWDL��P��_n3�R��Z{P ���#����t��l5v��C{Ab��R{����q���S�~h���W*ƙn��F�Y���]Y�h7�t��$0��SӮ��t�<�0��Vç�����!�Q�����wS�l�%�`���8��M���Q,1 J�L�F��6�^��-[�p3=S嶓U=����6%�17�~��&���A�y��T{����V��RfA�����A/̔�������"���qN5G#d,�%�[g#H��8����� `a���A}�� �%��K.�^"D���!����#�� ^�-�h��|Eϰ~�d����>�Hz�WZ�^S5�����+%���y���'��eQ���{>�("�W�tQ�"3:�����vyj���D\ǐV�[��uiq%ԜoR��	W$���H��[�nBU/BXpP�ș5U��<RAM�k�wd�BM�Ye�wnhO�����bk�U�ETR(V������I1?e���rp�a�\��$�|��H疽�c|��}�+9� ]���ʾ�ħ1���X�[��w�/�5Yu-ܿ������?tp=�
�6V֊�^u�<}�0"� r�|v�n��� ���As�m�ܣ(y^��&9h�M;��	�}�
���IY'@k����퇫��(:���]��Y@p�&ԖK5>%(k�Y�f�)�n4���`Rڈ�}EX��hP�'V|���Qs� ��\ëYJl.���_��S��9�e��/��1�{>ŷ	c�&�N��M����0fo��|�8���3M�@H�0��{�qݥe-_�y�B[Ro��P2��M��ۈ"|����r	4b��S�$撇�u��H�0���f�٩Y�E91��YK`���nΠ?�M�";D�N	^Lj�-�ɦ�?%S�y�����n{I#?dtƓA�IT���g���N�F %�~:u��R��cQR`r��`�Ɵ*$�����B: �i'.�r� ,H�eŮ+����2̪�0�4�e,�Il-�}'�
���3��_�7�O��q��H�Oa
fg �ӌ ���`T��Ǚ���B�G�ңuCR��R�/�N���/&�	�p�XB�+����X�ccT�����\�:]�Rўп\�et���ޖ�o��b�iPF�22���%����R��"��l����%i7?Y�Y���J���H���>�'�Ξ�[dam6�Ġ�X���r��%�D�ꪧp��x9T�: �-G�N�s��@�P��tØX�!���bB����}�b}�*I�EboA�d��N�U���O�L
q�uGl	za��vA�)����-6m��Sx�g���.p�QPW.Zɇ�� �i����	�&��M�)�%_K�w�*��v��g��y��.�TR����gs��lb~Sʆ��p�]�%��f�Ws��J��\)Sɴ���$�?�e�]�1hRTg�zWZzx��kL�5�O��?�����.}�x�Si�&`rF�1P� �bɁ��H�8�cmS<	�����W^�Zjs^�a��G:0Q�:�F-l��"j:�99�g�@!pv8�̿��@R��Q׭��A��AM���f�x�=�.�T��<�ԧ�2�F���fQI�KbZ����B�@��@���sc1,W�[��W�7�ȡ@�3m�����3@Y��iv.P*��Y^�1�p�Nރ�=͑�Z����%���?��I)��aV�'J���Ⰳx�r����x9x���O���s>%"�%��Vt�?~�J���hm0�qH���V�dX��7�H�^_:6��4g���<������/�h�r��uE�\5j�E�ŀ��QE�D��D�$������SS)4�4�R퀣G�����||�����VB,ޚ�l��$'��K��vz�j�5���Y�����1G�I�V�����������m������X��+��� �ਖ਼�O?�M����������O��+��6���V�����V@˲Ѷ��\��0�-���(z�[:��|�:��ն�4�c�	ߡK�x�Y�q.qU]kj��!UH�-��k)�;��B8\]H�D���]��(�L�cɢ��5>5r&�l`Ҿ9/�3��{L�Ÿ q�6'��:���!��7bYu�ŧ�*
��vۢ���7%x#KS:��6r�e���*�p=��f���/&���n��F�::l/ˍ�*�kЯ��˴��`�}l�
Tw*O+�ۿ]�z|���o�X8����F�U�H�u �f����T<H��RF�4�B��íl�����J�(��z*98,]u�o���駷\�~�~KJ9i��W~ʡ�f�a��ψ!�f>�f�+z����ҷ�<��k1ؒ\L�$0�<h���ΉF�%9F)����|:P���<�j�=kG�F��"(�n�F/��{<�Z����/Qq�2������� ht�v��k���cBpx��7d_����jrC��*�w�Ȇģ��մSܵ�;<H��w����C��{�K���
�~3/���x|�g0�Yg$a�s�{�|b,�N��xi�#�y�ǔ�0.�q�b��\e�T���!t��@����55��AJ6 "Y|I����Y��f��:-C-���mͽ��C'������.���yYR��g7�B�֥��+pu�bbd��ѝ%2�]�X��>����w]/�����X:n\+xM��jU���g�2�h�bs���DW��5D����R��q)&������]��?��������U8�_!��a�~w%h�.�'��s��zF9*]=~�S���9�N��޶x[-7{��%0l������&atJ�[Lہy��ƞ�H�7k�ؠ��l���{��`U)���n��8Z���s�Wݤx�$�,�HҥO6��1 �p�x�/ѣ$�»1Ǿ�6�f˽�)%� |�)6n`�{g���T� �!�ӲQ쵡he�iu4�h��3w�\�+�N� H��,��6�`�.�Y�	"q���x��9�!S�21�s��>N�t��/���p��'��9�|)O���r;�蠩�\b��������&)+�(�P��u�=t��8���B���332�"~��K9%e�G�[2Zcfjq+yYm �Ϛ����Nv�j)r��j�\���� �5Zc!���ջ	�)�m���<3ăGl��=�lhv����d�]n�(c���D����
��J�bi�a�;?|���Q��T��b0Ej��F�$/URz�RGȆ������G�V.<]+�䯎
�X?��at���|R����3�6�qF�Y��}ꗾ�����!��k��KȒ�u8o��4&��>���CI�%��w��¯�skʃeez�����P�L=G�r�!҉�e���x�n����ΕV�Ғv)& �����N|�P:Y��}sjE1iZ"���1�I��,J����	���:6O.�V�q!E�K��p(����P�՜�7��#|�:a�.���\��4ta�߮��(=��Yr���V��Z���a�T8}�����D+�-����������ί?7����8P�����^��0U��=ƥ&��D�Ѫ]ö��s����R5���֞q�TM턗��>vJ�{�f����w4��U���oK��m��s���F«���>��(+3F`���X�ں
�H~�x�]Z�z�����I7��"�C`
�<�R�Z��Y�����n򡌶�)R��9�I����#ɯ����
d^�I��3:BYpP��:	G�tM�bL��[��b,�mk���̱�/�`A��, ����N�t촺�p ��=-_9���9��KI�׸q2;�.�>�N�gt8���[��0e��@����SbE
1�a:.�*sϛº�d;r��碄��0S�B�f�>���cQ���ؕ�%^Eyq_?��s��rl��r"���,)Oq�z2;EW�%ѯ�XhOszB��qY2�&�z��	*Y���� ��.X͊X��]|\W�3(����ҟ
��V��F0��q��'�QF.�ǚRO�ފ���&2���2�ɛM��[���N�ĺu}V�T����oD|����5�g5��:UX�F��i��on?��Rzi�J�/ZVH�z��J��u�>�]��A��+͋?��>�t%��[N>0S,�k�B�3�0G�-�kơ��@w�@���򘀬c4��ο\��sq:Ks�e���z-\t�r��6�{Ď B��E�,N��e��Nc#A���?ZM�P6(a��(�����Q�r��R��Y�a6fO�-�Յ��b���P^.r6�w�M(��7� 0�O����m)��7r�����s��(M��r�,gv�p�_j�%e놑1c `��=�2��{�-{>� 	�x2ep�����,٨NC%C�B�!Ar�����	�L��hT��{� ���Ԭ�|��e`e���eE�L�MV�±N8�y�;����<?���9���DE��3�YL����|2���yE�I�I�d���ћr���,#b%�ҁ�����@���И�V5E��\�n��7�jT��]z��V��5����0�ո�Dz�/�胭?eE@�m~�\	t��zqN���?����C�%� �������bYO�H_i4��!i�t,��r����������J%rnсAeR��"ё�V��к�#��(�?VT>����v=$��+و�>��������xiBٙJZ�����/Y�ŗS �7`"����,#3K�lh2�V(Hw�'�8�s5\��?�9�Ϣ/����Q��;I��it��tg�j�.,�Kc���CV�P�&7�\#�3
�C"e�զ��B�G�;)�fЇ���[�����'�Z�^6s�@��=~(�J����~����Y1�/{>���߇�a�#�}z���!2���k�7-���+��-��Fug�'\@c�ʄ����2�x񼼻��zW�V|�>kS�e��ݣ�~�-�i���$�-����=`0Ip�A��x! �
a��E�4����������f
H���{G[�=��*#Q�|/�� ���]c�F��_:E��H]^��CsOVN�q��ݘ�Q�@#�/��cG� (M�^�4�S�^5/�d��t���x�@�����]��v"�e��v��Y��'n
J���Jyz�F���#��j(�.�F��Л�&f�����4E�����Ֆ[&��B!!�?FC�Wk��!��fMuĽnf��/y��=P2YY9���h��ym���%~������׺�:��ѿ_6���sR
�'���%7N:��B�!�����<>���m�h�>u��"����BL�ÁC���١�\�5p�
+����ø��:Ѥ�L!2ks�U]� ?@��f�N�Yǋ �<�e���AV�U@�n�-x�A��>���h���D��\���"���q$�e�n��,��r������Vk�jm���6�P5�(�;=�xm;��0����=�pl9������0ﱲ`^RCf���]c'I/I�{���:bT�aA��U�"�T�����.��?�>�A�����d�.۴`:��d7����.2��
Āg�d�!�[F�{�
�xڀ�f ��v���a�i���+<�i�l<9�%�Щ���X�t��Dv����a
!��C���4�$�]}%��RLk�*X�A�$TN���
�	5�Wn���6[nv�hK���҈�Ѽ��lچ��;}9F��[�E���հ�/9_��eʨ8��t�_ʆ��԰E�]ThЌPͽXg1&�m���/�&��,RBy���Pk�NA#2- as.�RP^������bJ�c=�N6��7�1�T ʣV�ʝ��ʅ�݋��AA~d��`P��ޜi���w�������Uՙ��UI5�e�J�2�����}�R�o� ��ܼ�iM�ު%=��H�:@QDH�����5�]����3m�>-i��n	E0�N�8�8�/�\�A�z��Z+�
��8M�6Y�>�}�ӟ�v�������S�F�潍#�NP+�NO�o˲�z�X(�KqM�.�ϓ�GWa-HP�z��`�Gɫ_8�����s�:S;7H۶�O4O�Ay�����[0Rc�l�b'5����C+���νZի��6V�W8��.� -޸������*`_�5�[�.ˆ����z~���\����U�D+>xZ8P�7�T���`���z�Jrw<;,�J-�-�{�P�^�⪋PeU��� ?��FK�����$~�1�B3�<�\ص����*���8a�n�q�h�2��d�, "�&�׭�x�}-��&��3�6��$
�UO�l���s���pH_���[Z ��jdTƟ_F�'�O�,(��!���gv��\�ѵ@q��P�gC;�~k=�+��
�����ɢkw8D�o�;�b����G�C�<ʥ�`�-��a�vj�_;P�7t"D����`<�i�����,������D<��^�3$�j�.傩��	�T�nlmh�R%n�� W��+q��a���>R#!��e1������� _0Ó�P��>�7��c� i���� ���;Lm�y�)D��US(��a��o��c�_G�R�s:R�{�����ҟ�^�x�xǔ->
>��C��*Б����H��.1w�)�B�Q����LT�����Z�A.��i���e�ʸ!r"��������A���Ɣ��P]�a�)���x�������L��^;�����re͏�Q���8�V���R��f��/'�ˠ�KȦIi�;2[_+�A��9�Y�w��56ѷi�6$����f������T����טR��Խ(�	=�*<������Ĭ���(���\Kʇ$��7F�UDf���	�i�E�is�%n{lKo�!�>���h����s$��cmNJ�����8�}��.�7��L��ưv�sv i"��<�U/n�l ����	�M%�ʳ��b�������!',�G��D���й�*�%��2��v>��Q�a��0�7rxy�3�Y�[�����"���I�w��*<��Z�����*{���]-hM�����7Go$����h��Ό�z���*?��@:�P����f2h./	��iL����}�w��z��v��q�*GDJ��N���� B��☊KA�/2'��U���i#�C��N ���I���|�Hlv
���������k�l�BO"��
��ۃ�D���q�l4��k�V��,R�B.meZ��Kێ/�s�.����$�C}$�$Ms
�&�nR+k��c\j�ܶT��x.P��38|���������ޥ#�rG2�*�|b�!���}.�]��C�ؚ��ͺ�5�9P<�%�@'E��.+ί>7��q�P
Sv��PG쀔��bҲ��{�%]P/�]I�?�j��[u[�Nbq���~�f55���3����{��k2ӛ����q�c�I q������ �}��o��*ex�����TM3�9���0�&�I���b�2L`g��ɻ��B8"蛲-�Q=П�!=��7
�.��4�K�*V%*3�@�$��H~hFZ�%x�'�"b_&��!��G���m!�o�O�%R�[�h.>C#�ZG-���v� 3����*��=��cW^uF���֦�wAW"~�GS��^�e<�Q��u�����R>�cbk�E)�$��ꋐ�z��Z��U��p:ׂ��k�	&�*]l!�
0F�P���QiOD��B�u8� ��k�#;31R�K�i��1v�e0���Cv|�G��{��*�>�Or��E.��_D�����l����OH����Yc�V���`�0��������ʦ#w#��p�vs15"w�|�� �?�����2�Z�vQ\wjG����є1��1aj�#[�iS��b"���Q�tY��d�)�̎|�Xɖ��qa[�n�!C�(Je����0�F�3O�8���0C���M���Ķ���a� �B%��g�h1���%Y�®�8铷1P�y�q<N���}�痧�ە?��7)�Ϣ��z놤~s7��ǹ�� �f7,�K+�s��7�!I��l'B��rJ���L\Ap�(�|�*�}@���*�ٮ�b<�W#w*�/����оK�Û��%Z�s����k�B����� d�LR��7P\�ss]X��s����(�fH�a�Ψ�W�_�^&3 �9����[���o�k��	��x�w�6���������-K$g�a�F�$Y,��GT.W�j�h�Њ���(�k�����z��`�SD-2C������#��/(>j����X��&[څ�n��2sP/^1�-�nm�M\�1+��MɔW�"�q�ē9
�]�>�ʁ��������~!���<+\;Td�m�qe3-����Vx��C"r����v��E��ǹfny����;4��V��m}Qg`�X<UH���B��N_�"u<�=1�Sj}���6W)t�������(�j�k}la[7li�z��VIvlԷt_��dy�/;\[)@�	W@ڿ��|����"�Z��ߪ��J����	�IXR���bװe��OM�	T[�f'֝�b%�%^d�o�����h��x��9b��;}~N�����<
gr�7�:-L�./�
n������L��0�z"`�M�0��dV���	�4��Ȇ8戃dv���M/��+3��l�@G���mH@Y*�����Z��5�cz�����vUoAq`���:�� B�'���Hs��ϱ�6��VA���(~��?4��=\:yꫝ��|'�;����Ìnԁgk2y�cBa��&�\���-͏(�:=f��cQ�nԒ�t�9���?O="�"�cC�O⏁��K�1{����m��@^�)��%[HI�G� �����F]+�^�}آ��9 |����.3B��~�}Z�|�<J���uz(��Fm�{���~O��/oL���;2����~�7D�X��l�n��"䢝�C:�y�y�T���i<���Ci��e�8���<"�<�r ��wͫ^I9a�%�ϩ���Φ�H�?EkW�"4؍��6K�H{�Z����R=�-���v�z5�����Q�zX�_��o҉>֋b�����x�Fb4��Sv3Cz���Y#9)
4�k]fu��qd���"#G���Q��GWؙ;��(�]����p�}�I��`�=���msG��W��Ka�:���ֻݚ(����Q��n���0��
H�p�Y��}�]l������.-��K\@�6Eh��f�hE=y�k9��L��`@����]�dH���உ_ɒ��r܂�&*�� �)�-|AXr'[q�QU�CN�aF�lQ�m�W� 
�KH��Μ3u)}J^�Oj������C!K4���uP���63�L�  �ӕ�����qV@�x�X�?4Z���y�{V�W"1�\���wa=��$��f5R�FmÏl�� vp��R�|7�لyQY�-�g�=}&Y�ֆ%+/MB�����V���o�
��^��@"'�n<�9�9�����"�J��mm��� �"�R���|����.�̕��b`f��H�����jB�)c %<�oM���N\�HO�V����)����	VY�p௲	��
J�_XD�-[��E7_��ͽ��M2��.{꾪�r-����Y��2�/�(�`ܣ��&�8�A�ksmyHxqQ�9���Х��ÿա�=��s`T��@*�=F�#���1��LZR�����,N3�c-��9�EmM��c�!F��@Ϟ/�=�0�� �җ� ����>=سI�9�}_�f�9��#"E�_�3npe��.@�����ey��x��B�D�
�#�ǋ��8��/�?� �;7�<U|b�{���.�}�������VcԺ�c��{|�@���t^��q��l�
��l"1�![ yZ�(Cn��@��T^���8�~;C���#���x���$�kp�+CYqBAŕ^F8������Cذ2d�$��+�`�֓�~��k�!���������ˉ���Hk��}v��s�V^��IE�s���kʶ�5j=����[;R�n�K����C��Ѫx�$�<��KA�L��G���a�O�����Y��)Q��sB3W�nN���U�!CU��=g��>�L����ڢ�z��+;��\�盡
�pP�|M�!�Am���J"o�
����c�F���H��<&zӱ��s�.e.p��:-tғ'���]۟���qSd=��e�Ԑc/:#R)�2�l��O�S$r\X������O�u���̷ܩ�Jn�
�Z	{4Q3R��m��@��5%��e�$Md
gZ��be���s_�	�}�;09�KЖU�����/��w�D��Wk�͘�D^�F�'�Lai#�E=G��*�q�R2��f��
�=�vm�����ҩ�d�c>�9tW�yb.l 
�-�7�iax��l�RRx�t'hZ�A��\�%��Y�����p����ң��9q(��e6AsR8L�%Zk���UT�A[�&��EPo����|����jC��k��8)4�55!4T��{����#U�u�1��k���>m\r����y��lՁ"�|��3��d����0��I��Xӆ$��P6��k��xï46�����%J':��S��kx�I���8k�5�Υl��/��DQ��l;�i kn���Z�݈�f`dl�a^��M��7�C"~wנq�aE5��G�?X��I�_X>�``0mK��O�/�_~|��r��/��S�ʂ*ÙjJ�O�S؇Ę�������G�0��s��jL7ȁ�*�: Uw�Ȭbk�������j�[�'����g�Ďz㥊���8#)��vt �����z�6��K.��s�2�"�o�����U�0L`	���L_�I�' ���W�ր���[�ʨ�Fo�`� �3�fr�输4�pR���1���Qmܲ�@�?j�7�T�W�����iXH������0�i��(��wPS�Be�k�ыVC�R�����Q��M�z�v��Hv�1,6ywl��`�n����Y��!�e#üX�bV�1a��LqS2����o?T���z~���Ku�S:y,�I!r�l�� ��F.�������Nŕ
��o���p}���@K��ت+��,�^��K�0���]SJ�g���. �����s�EaZ��r�%�v���Z	h��
���5���O(�������?du'�=�(�����0&X@F��𳱖$Q���oA�>��j�%E�D}q���WeN'Q
�Դ^�����p���gO �'IR��Ӆ����Ϧۍ=��L��j��HFVr?!z�5�"D�~�4�l�C)�������ʉ9�غ�9q�),���L3Ւ�4u)Fh#h����ަ�L��?#ӳ�j8I�~�C��3,s�$�	�Q.�z�;�0s3Z%1�V�}��tyV��~lka��� �xX{�;�u�u���c5����൲���Y����#��V��w��axy��9��F�F���X����l�@+9E"�#��G�"V�<�ƘE	����_!h������p5}l���<���2M�6��c
�\(�C�s�Ev�6<�<m�N{���Ch0�Y�Wv���j����x�����RO���K�5t�3��n�h�آ{07+)����ׁ�ق���u�9�Ȏ�4�xH��@�- _�esY/{&T��}V\�0iI�Y�y�1Gĝl'FTcw�$2�m�y��wC�f�s芌	Ο��U���Z{����j�0�;�w����p5d���J�Bb�'�P�����㣌�5��Hn���#OR$b$r:v[Ŷ�I�����e��j?�D��#�5_TZ�eS�wȂ/g�$�H��Km�&��!����kM�������7�¡p��]�BX�0V��E�v��:�B77G2��wN*�6W��_St�$�[Ӧ�J��X��m�5���1h���WqR8V&Mlk��8t�L蔄�vp��������s�%�%�"z�W�F$蹑���.2�׷�)ʕ��V��ݱ�B��B.wrIaN&ړw¿ ����?��?��1N>\��-�=k�1��ߞ]���zL��tO�i?-���Z_l':�nu�uH.�i����&{\�6��� ��i����������U�������3Փ��Y̶���Ǉ�|�,ֿ��i�W݀v��r����WS\0w>F	9b
V����ᰇ��^l��Z�a��?;�@�i��1������-f�}g��(���Ds<"�ܚ���1��=�>���#*��5l��ݵI��+?�prk���w8"�\؝�0�)�3L~"��b���Hl��dE���۸�x��}�m��ߞ*x���F6�Ɂ̇a�[��1�|���K24�N*h�K�M��ZiI�t��x6�&a��ԙ͜����]TH�85��ʪ�ÔkY�w�]���q2����ހ�n�mыF���,�i���`z�<m.���֩������3�
���是y��U�+	�t�7�)�2��cЂ,umg?�T���/��?���|��j�к`
���_��*���?0�4|������K��W�����O�ќX�NH�6��B�e� �9µ�ķ��m��,1�ߊ�b�P�����6c���;�è���
�l�D/&;��vewub���φ�.��|5c?c�t��R��N����y/V�}n�^W������}'to��:ǝqJ��A3�GU�}�ld0���
�.@��L�J3y-�R��Q���N�7y��@������*+'b|�n��w]�(��p��%jp>P��ITR�7�A�S��t�ͷ��&,�����;	�AC�eZ{�_*�s��˴����p&T�"�t��4|�2���[���Oo�(\��]q�ь��iQ���W.��8����;��!($]�hg�&H!�3�{7�{˪����lHA�'~�dR.}�Ye�vp�H��Y�<�MR��gˑ�E������?X����U+gC��D������Z�x��վ�C�}�������I�x�������[
�j#s����pL�g<˶g���L�W���~y�r�,⾩�HHa�>M�u�h�$�=U�vE�<�B!+���{���S���/M�{T�� m�3S#x�j�|q`<9�"&eRŅ�k��.K�����TWb"��P}H�i]"��k?�I�O
��,#x[i�5�3eeT�� �\d���N��x��#�va��ڿ����E8Px:�	q-5�Va���*�:�����+ͦ�x.)�f"}nO�\�����]I"�I(�̼��� �`�(5l��EI��LS?U٩v��u��|�lU{��s�K���@��.��,s�*���FY�!|�u���ܔ����K6�?9�^��q-��.0�X���f�\MR���~����������c�̒�׻~X��ݱW5k���
�ʤ�}���r��N�n�K<Z�l��Ka݀6uh߈���@<�}���g��.���]�T<$�i�S�Ϗp��$ژj�K�e�4^g����x���N������h�����>�S�w�/:�WTpOC�~��=|�#[G����XI�8;�?�ҕ͞�h����r�������P���ĝ���SfL�|��af �v�~L�g���9m�i\���N���~Ĝ��z�1�p�˯�@̶�k���$-J`7GC�S"�u�]���Y����<]�vZ�����<�M��" �j����[���X0	�`�Z��FH�ndY����ї'{�-�p�{ cf�?#�=������c1�L8Ugv�����v
F86,
|���#!�>+bwe����T�����.o�d'0�c�F�����f�_�9!"p��
�orT���F�����Eܙz{_$%�@�K�ھs�����Ͳ��V�>�f>�Hkӿ��R_�����2�.�&ǲ�,�3
C��*��<���%���`���&���Z��a��w�5%T�I���P�����fA��@,nZ�6M@�O��1����!��3)��?�b��Us�s'��е�ԑC��4v+�����ّ	��W�a�Z-?�b�_�Y*��9��A�LHB0 /��Tc}��j,/1��Ț�|j�!�"��mj;}����~$���;Lc���[�n����4O��+���Žr��}�W�&��+@���!l��k4풹'��T�3�+�K��eS�� ���u,��!��z�&�$���z#����t�l�XG�)��a�����%�K]%a�SLJH; ���/`<�t��zel� �= W_���S�Nb����H�Y8܏7�,�E�.�zK�����8B��z��	?�"VD)l4
�Iw�+n I���������đ�i�CC�j�t��N��*�^,��q�-�lZ�R���Go��>�& =z���z�C	�j�7����Tn�.�_c�x�s��OR�:)�NKo	o���dٯ[Me�G`�-�����������Лt�׎H�[�Q��m���1��!��֑��j�,l���-G���"d-��

A9��>�38��=1.D����5"2��֕�2��o`�Ru�;f�~E)�wJ�Fs+p9>��f���?�S�<�MV��1��c$��h��T`]����n;��|��c�6c$#Q�k{���UFn�!pc���:� ���*�oNq�obb���ɸY�[��P�:�à�D�T��r��s�-��>%R?~kk���f�_]첟�_�_�e�h�&iX)�x^Su�{� �=I�jO�(�6�O^`�fh>�m��Ϡ�@A��O�vB�>5��N�|N?����p@�G��d���F�݌(�F����c�p/Y4��;����&⫓��<]l�)=~�=����jS�Nؙ6ӝDb��Z�0���餒N��_&�LC��`�R�#�S4�DF�M�~>�=f�ó[z�me�> ���Nr>�ڥA�&��0���$.�( �y��g�7vH���h�}�R�ئ�����G~�7������10��<�߅�o� ��?�#SE�>�e�����5��*i����@9~�Z� ,���R-���{ �ξal`�����l�NV���*e:���I ��#�¿A��yNî�*�`��?�Y��2(�#�s��^+����$�����8|�xPH��I�>]�k�*i�&�e������*�|����)�N�tu�Io�ߍ�7X8��>(������/SH�rj����:��a{n
>�'��;�êBDC޲O�Y�F�i����S����j�7pv%{qpTUh�ư}F�h,����2XV��	R{�Rs����r�Y\= �V|��4��{E����� X���~��o6�F)�D���v�g��Ԟӟ�R�gs+�m�iEЋ��q�Oϩ��>xY�
Cl�1?�?��E�ȹ��흮�"iqZ��������TԜQD�ӮMyj˷��ZD�U_l?z�ؒ0~gw�'֥�[�%h�֛���:�lM���c�0���L����jE��l$r�J���b�G1ãwo�˲ݢ��"/6)e���Q��>��+!���Ơ~Wvm�|~���N۹�uHҁ��r���!��åq��fE�269.��r�ĳ�T�:i�`~��z��Iƥ��g(3d<E^Y�̌�<�����qot$_oc�����u'7$ƒ�+�QoDB��U��WI�nR֌B�[K��f4OV����z���mw�
 �2:������4B�>"W��8��>řh,Հ�S���{��EM9*W��f�12.d�rtk��e�9͡F0c?�\����n][pn��." O�I#�E,�m��x����0����Ø�$Q���w-�z�ɣUDYo����J+g�Ϩ�����Q�ߺZ��T�$����|��;.tvVw�/�e/��/k��7�e��iV7���P��4�n�q��Wd+'s	��2nΚ���_�����FIt�B����J�Oc�ӡ̅�˖/ze�<-��9�`�zQ^���'��xC��+�zWcY�P�Y;�J�@ȢC
3�r�-_��D�ܫT6�`F�ZBޱ9?C�Fch���K8E�
E�;c�i�e�iMLo���O4��I�C��[v��J���"���K0�9�'&	�������c!���I*r.q:4;Nw=�^Q�.�/ ��l����{mj�==���GSS�ܤ��C�#*�CNp��#�-�cdKR�;+EKP|�xi�N��F%�n}��_��!�(R��iU���O�繟�c`��t�v(K��}m[7ICQ�6�5c� ���-�a�êZ�q0����7�{Ȣ�wX������^�
6��W�>-r�~���K��_^Y�O\�>����=�.v6��O��8�M"��6�m�Ф�&��z
�����Y]2�8�6�T�{�]�(��Dz�an�H�ҩ3����?k�GZ�fCZ��?��Rm��$H��[b����eu��SS=Q������>�?W�\qMM�V��t��"�ADؽ��d����Sb���O[$A��?�m��J.x��R�u�c�Еqt��o0L�0$|��'��M��P�~c	j?lo�"����T���=�VM��e���q�(n��q࡮A����M�U�Y6���a!c\�]>�2�J̱9u�V1���ѡ�F~>1G=����c�e����[��l���M/�5�q��:���|kQS��������0���A�1��O���e��N���yd�]20"�0G	�Rq�ڣ��[cub-h
�Tlƣ_�hªd��'{;��-����"Ű��ɒv�ca<�v�j�Y�HíHL�@�i,�!�MU���f�yjOM&�X�Wq�/� ���N�F���)&��F�[#���"�嗜Ү�h���QJ������0�3��V�+�]�e�=�ҔkX�#�Ǭ��:��ok%��N�#M�D}�bAܟ,[4�G�<�ў�����82zi䟒���9a�s*�T^�����Θ-��v jK���+���s[�>jc|tn�k��Ǌ�tlj;��~�{���*��Iף������q��*�`��Y�Y
86Y�����0[��/�Ӻ3�n��wm���oP��Ѫ��^:���qn�_�^S�rԐ���M��V|�k(|� 8bh���BPhQ�Tv�R�
�&��+�y\��8T@;����0�c�l�[״,��/�6����7j9"j���`�Z�ux����)�biA7�l�2R���5�9���Y9�/3��H�m~/�Wy�r���ZkFO"O'Q5	:\MO�H24��Ҹ2���f�b�O���UA��S��:� 6���<�����F�b�ć� Q�Tֆs3��|�#�a<L��}A�7'K�1JT�$RJ��U,����֟�Ωt�x�pO.�N�t߄��{oJ��n k�J��� ��"�zI�^=��V�s�⩃a�H�`��M>TځW[#r,q%��<'���;��k�6%>��]�����	���	�K�D؞�[BI8?��;���1�ɵ6Um�%���i����bD�ui�ЀE
)���	��n'�슎���t�SGaY��O"�3^gz��J'�@$�����Ķ+?���.Y��<�������#,B9�V��Ġ��e��uopA���A���w���@n���(JI_�����,̾&I�oo��t���}�?�,BsD���� S��-e��a�$� %��e��B�V߸�LR�.��a�D�[��e����z��4Vp�.��GC���>8HM��k�_p��,P�!Ъ�>�ڳy��g��W�SϜ2��Ȕ��uuФV�PL�ѭ���FP�w�����|�?8q��;
�I74f�٤����W��/�����oG��4ś1W��� ���kϻ����1%5��4��
�y�׋/h0����E^=�O�m�e����ۣ��
-&�3�I�n�X1_���P|R#A����h�P�N��*$�F���;8 �V����Cr5_y�������qQ�CVi\�ہN���ց`��8���D,ٷrl)$���l0�l�@	\2����q,^��)�$����˴\+����WJ��٘���[��*�/��y�C����Y1�,����������]00^Ϧ؏�Ӆ���[�=_qx|3�I���2��M���-��!)�ݛ���\~y��tv������)���h��<�1��:|B㯞�A��j���ZTE�Z��#E�:�3���|����Šm2z���A�2�5r�es�h[ff���q�^`�H�y@*~)�ݔ6
��8��q��o�mm���>	ּP��=�(��ԋ��� b��De։�6�?:.T�i;W�.�d�t����`v�N�`�'ę�����|)Ej��2{F�=:1�y*��.a��tX�E>��>\� ��	�F�����˥C,��J����9��՚�����ssP�(�q1�%,3�L$h[C��4L��-���2,]Ҝ[���/�L����P��$W�G���ģ4FC�jA\�xM���]ظu�ŨS:a���?�v`f�����h� ǷX�Ihw�Y��~��T�M �G�R4������r+�N��~�Y��^�\��3[Ǐγ����q$��^(�P����NW�@��/+�zɥD�O��`���~��ȣXؽ���?* � YZu�dfp�*�"�V8oK��tO�j�0�''����ZB�0��7}�<��~��s9]̂q��IZ`���P�l�AZ�>G}�~��9�)����Rbz�|��@�g��8:4{��h�rY����	.��h��/ia*G���0�z#Jʏ�P���<�G}�*�E��eY���8���+�� �tÖ������K2q������qbX�r�u92��A�T�#�R�}�#���&��؍����A���iF�n�  v��wr.�r�if[���2�G԰�J����P�_T]�9�Zy��#n(����Ѝ�t"�9��'�I�A̍��`�`3싂�>�d�z��Go�K��1׃*Jtp5��B�<6�J�[��W�+9�r����n�)أ��]�����5)�I&,p�;i�1��Y�,�� �8�lpH���4��m/�ā�G�!�K�:R��:�J"�,�s�;$���s�g�w֚T�$�]��L�Ռ"m+! t0?'KXj�-��ѥ^ЏU�vR�>�����1(����c�t2(��ב�o���]@�
^��m����ቷ�����z�.`"�ɚ0��Нf�VV݃��EU�UO�Y��׷.�lF|�,Ч��-�&���l3r�D�!�$ڄ��Ɲ墓��?�@-n��vA��B��c� M�:
B}e��_;.*y�Y4�}b�Et3w����ڪF��ɫj�>��2�:u�����=���++����6m�UL9��Q�P��n���<Q�!��`�l�Jf�a8t�"��`��}	��%����1'�w�kȽИ1r�Js�j[�;;�mg[ɘ�Ŷ�������E@��!�o���ߤ陶���{i�Q���):f�Ӣ��	#M̮��`�|AT
����2-�1��CgU%��vJ��.Z�2��)�s��;��0����3Cnl���-�#"q�s�ab:��FX�k�>3N9x@�?wP��i-����#uV �@"���\�=�����/�{/We4�;tҷh�O�VJ���j�C7n��<�Q�]mM����M�}��rZ#���o�:�����ywh�ɳ�wi��O�ǲ舭)��1ҩ|n"��=�s$�9PU��o���i�1���0_�NZ.����i���'U:&��6+�-�+!���B�ɤG֪�-�?��UoӼ�7݃�F�-e{��ĉ��U��r����k \o�rH���Fܥ:�ϸ��kE01E�� �(��:�	i_�K���C0Hq�lgcwC��q���QZ�0����GVq�,���t��f̭NJV�����r����ȧ�u��M�Ŭ���L�%�Y���E~�״d��>�B2����c�w���ŀ�m�F���E��X̨��u:2s���"t��^?��rt_��4��z���d�ؑ�9��C�wG���>����(�4\.
V̊���iэ�=�A�}�S̲OΜ���*������@��y5vV����h��@��?]=�H�Ӊ������91�.��ņ���;%��T�+{��o���������0�)4�rݤO��}���*_�w4�)I��8%�ӻ�ӻ�Z������e���|�Ga�X�l 0<7+��e�<bIc��6�Yv"o��lY����%��B[�n����/��)r4��E��â���b���#���e��k���X x�1�\��� ���9s~�E�z-�:#���S��u��-�Y!��� �|�xr4~a�]���64*�L-�b�~k_�Y�t�e��k����O؆�:�`��!��n|�1�PR���`�N^ �
C�S�m�I�8��^�2�2�?�l�����	ͅd�ZD��p��'S��Q���3��ü�G"�U�����9"��)3K(�8Oh�&4d���l�px|4����Ցe����E���>b���,�ِ��"w!'U�vҪ�WMvf�G
O�#��X����� �$E%�L�X�s���q�9���o�U�4�a5�S�Fb� B�TΊ����-"@���֬T�a:i�㛃���=P! �Bru�L���e駭��a�}M\\�QZ��ƹ�!�������/z���
Mq+�:`����َki�R�n��dӹ��5�Z�R���ø�Q���@�*f�}�͔E�g�X��������3�]����ɠ�c����w�L�{�^��W�q�gos��r��ܑ��[�riX��:aò͐��v/�����`���JM�)��OAqM�M<B�D�վ�HA#o��߁A�s=�OYhe����5���3��pZ���q��H�~�T����<0t�1+.|*�K7��j���]�s�f�Ȱ�-���B�Fȃ��q���.���6]�,X��[u����)d�3��>/��	���������$�3�)���N�똦�FN���C�S���G�p��k�O����|���LT���h�+|ը^gݠ�E��x�/в�r6m��2�;�E�.���,^�)���ю�Z��;�{ûc�x%/���:�u'���`��9KV�/�ZB�°̄sq�J	�U�ҭZS��uɂ����,C �8��� s����Ǧ�e+�gF�gh~�&]�s�������Lali��Y�u�y�X�t�b,�k�jIp�X�|� !"��l�����Äs|�7˗]�\��~HRM���6�}�ri^�%ZXw�״F($$d�_&BG&=�m?�yKot\[���2�Z����V�����7�=���.�LS�] f���#�z16y5�\{qÑ�|�Ik�%4L�,ǫϠ�A������i}{G�U!JN��QAg4O�i��*HK]/ƿ�h<����)� �W�Q�`���7E�}U�	� �2�B2P1F@�J.��-L�ER.>�Z�[�<�L�k&8i�R��V�2fTZ��#H�$���
C�շ&�M��8� �'�<$���˄	W�)A�r�?�FGܵ�A�d�@J�[�'�Е\�Q��������N�q7��Ȉ��#^��Xi���P&��ӆv��U�45槛49�������ޑ���j~m�L��/�|À�\qc�w-@��	�
 6���i^9�5�����I�8.c/Q3�
2�8@�0����0/�$��iBk����WM g��~v���J Y��(���(?y*;-8-��Z��>Ô�6�w�R����K@Bå�2�n�%�#�������QS����V�"q�=D��[���Q��Vr!W�Š%��PC�zS��-/����m�$���5#8i��{�����	,A�+m�mF���m!U�q�wiا��Ϳ&@���n�u7�fwp�R˄��؄|��K�FmM�����K�R��z�i��N�~�>��G���s���gG�5��=��#��/T�Sv��Tٕ��S)*���x�0mQ��s��O�Nm�G��j-Dܠ��,o��QL0�?X����ɘH��_���ԡ��eh�W5%$���_����f0
�p�n])?�͸���a�����Q#s���&�6�60�^��p��_���RZ_�S���:3�N�&2����%p]�#a��vI�"WD� ��@<��u�����gꡢ �T�N%x�VW��敊D�P*�`K�}~�5�7�Pf�et�c ]��e���I�p�v��p#ws�b�������� ��M����x�:�ѻ�"(�I���9����p�=N����`�gg?|�:�mVߣB2��b�=�����G�k��� ����|��Z�uw��p���fՊi���ۆ��`)sO)�-vȵ���-s��{1*-R��Rc	Oz�6�zŮG����ܦ�ՇGY��	G���*G.Y��A8��[�����O	}w��V�����.�����,^a�,	ׁ;6$B�Ä&Xd<mȩ�0o��vj�yL��2�}~�{�_{DI��B����߾��'%ٍZ�]̹��(Y���iT�eOJ0�Q��̑�Y�:}��G��HVj��,G ���)������LUQ��ӹ�I"��B@����-�^!B:�$��D�"nlū����k�֡f�nr2�6�6�/��&L�:�܈s�6/9l�a�/a��+���q=IiI��ܑ�d�xQ�Z��W��1uz4$����e�h��K��- �K�J~�W�v�ή�h-��>q����O�n9��kp$�h�2���1�R�@�Y߾UR�Yk���{������������$5�
P���JXF���?*`�D�x{�f�c���	�B|�3�l��(�_uI��ۯ���.���=^��@i��G�砼mW��8E%�s�`Y��7a]6T�5��cZ�r�����ڋ�$���TW�!cDm�%��yV�"�ۇ�|P.r[��TKj��HCti��+���]RH�E�|�*+���=���NjY�������Rqaa�8|�J^�H�L��Lu�m����]��>��񡻾�� ������s��Y�@������t!������� ��Ly�m�Z��dJz�K��Lu>�׹j{K�G�B�h�+P]L���Z�SF_�P�?{k�Q����ܻa��s�30'˂@O�K�ǿ�%ᆙ>�|B�L��ݢdQ���O9�ˀo4�/�
Ȃ\�l��O�[��o��s���[�G������,�`�oA�s�����%Xt�@�n�t稌0�ň�
U"5����~*>K��>��T�X�?�6;� �$��/��jǃ�.�*�(�$�����|z�pA���w~{p�h#4ċ/\o�s�WN�_O�z��SZ��l���w���������M����͑�;�����9��cv��$l �3S񶅁,�c�Y���y3*��wƦ8���0a7� ٌ�����~��M"s7g7�C��^^ʧ�.ܔ7P>y��.8�o��0�I�mѝ���I;�����3������,vO�N�V��� z�d��!������;��F����:��T�ҡY�c0��֙�3D�����t_�"EVh� �"D�"���i`3G�q���������)��y��y��h��9�O#���qN�Э��� ��<Im��F���!�!u�y�;\J5�y������J����tr����B��E�2�Imm���Eu#�6����<UnR&�d!]��2p�D	�Z\�̩.��N����#��YP`����ߒ4���LT�8qv9PX���#��iP�jes1�뢯�y��J���O���U�D<���g�rg}�.�e,[�m��E"�Kڔ��S�'�}ӣ�z����Ғcm��Mx=aE-��wU��?�D�a�|Qh$�]��ro�̶�:���B"9���VV���@�"��C�5R��Q+�s;��k��|���o��]_ 孓D&�g���	�&��Q��WңH�N�Q���9�H�|��f��P[y�%�]�l�+�x�Q}�Z��0Z&+kA�V�W�P)����)y�fƣ�!�#��}^�\��+��05E��68ҋb�|{��2�E+B�4���0T��@6W�dW�2hj�0A�6��$Sd<fq^���GJ���X3!<�a v��
~4{�(Փ��i1���i�U��9��lZ�/���^���3���l����B}��=?ˈU��"���lr��1��Ey�q��Sb�S:�b�9DU��[hH�ž��Eu��'���J��\�o+�t>p�׺�����i��_a�������������� Sqr0KSۍoe�d��	-��S��^��og"=Z� K�Say��)7�Ky��DA��Lt��kS�����_.�#iC�����@k�'>
�F�����@ ��?#�Rf�2?'}<'�d&��٥J;"�F��Vo�(_�t�>l����HU�a �M�.�;u��}��sq�⑰��A���!g	�������hUq�o�N�l�o��.b��$ v�df�&�Z�>�LZZ�Z��<\�1|f ���)��K0k<iu�t1�y*�4i	~�"S�Ɋt!��(���5R��8x%웽��LSU�8���	So?\&2��v�66�t-<N�d�S��de�P�G ����/�|�����ʓ�t���!�+D,E����}�9�}��G2�j�,�O�ˬ�HCyl�j�C�䤩���t�@ns3nv�Ul^s����R��	�^�b�2؞>�nЅL�#�ls�*0(��us�t3�t��Pu�O�{vZ�b\���
��=�/F�A�ysqG��R�U/d��7�q˸h�Fs� *s?���_[<O���R���M�^�\���"D�c�˼�F�<�v˧��2Rw(���������is�7�%�,P��,�<�XG���]�_����-	d�$Q�S�X���ǳ�����U��q#����Zm�Ȃ�N���{�v��N������ҮWꇮ尵��Ix�?f;h�?t 6�m�����nyU5�m����%��~d]`b�R���
���*� 9d��|(P�q�$y�X���}@6_R#v����1)��l>�����{_U�
ݫ�nA��C^W��K�XP��P_;D��	��0����y���
�R{)�G�&�!� ��7|	�/�����j��M��Ԩ/��Z���44�ʌ.��+ȵ�L�SWK�����zgN>�I�iv��7o�!��*_Nz�Q���L��$G1�D���I�g�#JEG�m�"�_�z;f��*M��c�+�������	�+4joNV>�γ� �[�d��x��k?��*�F��ؒ@��q��#V�&|e
�/��:���h�2���V�[�@�۾�Аaﴳ7�9a�8��x:zx��Um�!sV��D��Vs�,�k�@�Y����6�K�����HP���C��!��l�C��)��]�~�4�����VK�B�ǖk�����N��:	�'�\��>���Os �^p3�șxo^�L�&�"�sW~��W6�L�,�_L"m5���Q���˱a
ve&�,�(����t��A���R�����W�<�'�D_m�:Ң@W�����{�r��a���g��i&D1Gs��f�l���(t�h��*;��z���t!ӱ����F!���;N4#����@fp�p0}{��z�W	j99vobbw�DJ���t+��|Qc������>�ʟzt��B�3I���,v}Ȇ����ʇlX���E�1�`�V���򽔄tqF��(_�W�"��j3�M]\�����ǌ�	M)\��V�����l��EZ������VƂ��/U1���)ň�'��)Y�sn:V���7���r�?3�������/Ӈ��h���Ȍs��?�҆�՞��;7f}D�Ke"j�m����E�4�����W�5U�ު^�n��<7�w��Ԫ��	#$|���Mx cv�D�4�q�t�A��Ն܇K�'Q��hf��Ox�XŅ��?Y���Pp�zJb�<eKN�P����Y?���XL���XV��K�|4ǩ{�˃���p	b��XP���.��h�4A٭�XW@z��4�y_I�R��c��N�&��n��]��<o+W�J���]g��1u�ɰ**�X���� �����|W �hg�
�N]�����E�l�7�!�]@f7�{`�RfU#�TQ��9aj,;�Lh&D�xr����Z���g$
y��P�Fk�������Ց0(?�V&����幖*�z �F˜�%���j�5�5�ozH�?��&Ч�SbJb��<e�b�kf�xIm4ّ�v<g��&�8�`�	/�oP��
�v8n��S�́��a��CKaa,�`2޵�¥T[��T�}�ޙ��t�I��o�h���m�4?��}���ixZ!U.i��,��N0�y+���?%vJ�(*F�<�[������!�Mx%{�ay�����Ѩ����qgU��/�l�^��@���것�ʴ蔬x��}�Gj/.�ÿ��(��FQ����6q	�Tv��y�������.~j�w�)=��<��B�}X�o4W��q�4��sr�u�&�.B&@�h��@-^L��e��h �R��1G]�B�I"�)�VIX�V�zw����!tz����b�-�*�D'�vԟD����\�����=��͝fT/�y��K�I򦲘���_Ks\���9˞K�2?=��5�����\h���🷑_���^�zt �+�H\�J�BE8��a�_q����!*ǼvK���t�$�ջ�3�<ψm��E���]��"ڛx�	5;ö�sÇ�_kė_�x�`����� ��y��d�!���xf���u�q8������4kN��ɤ���Q��$]0�j���|@��D�5�7q���Ъ�>��k���U��:1������V.'�n�X�n�H0_�LD����'x��}��\_��!�����!{�; ���k����λ4��\�1�qzv�WC�ac�
C��[(�_����U�c�4��3��p�_��]g�	zg��5Fë1�m��%�$Y�.rG������ꛘ��C������a�tk�;�r1��&��[��x=�ds~]іZ_op�P�(�����1�@��8~g%��aB�@�C�-w��_׽}5��{ȼ�#����\,�����vY���g��L�i
�K�F�|����|?ԧ�6wWt#n�Jǲ��\��	�S��������Kr�K