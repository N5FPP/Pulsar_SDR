��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5dδ���KdXyݕ�2�j����B�}��AlU=w��m�C�}�S�[U ���c��6��u�������K���ֵZ$�<���?�ޒO 	��ȿk�Ƽ�o���n� �����4D�������;����l�{6d�0
�Z�^�^�2�;�D�
�UjR!�1�2>��Lb�`�D�l�W�?��9�J�ס�Y�u�kK$�ɓ�#�NA��Y�o�~8g�!'Q�Qd���1��+j�i��|Dσ:���x4����j���g��6��� n�벙s���c� v�f�GMcˎ�����0���6�R��$́r���E�^vq8g�O�jl\	��ч9ݢ���/�p-Zo;i�c�at��zb��M�պ@
�G{���CM��0Gm��w3���Q��ɛr�v�^7�<��cq��Z{ۙ��]l���gw��Eh��v|ۻ��&�xN�I��X�eъ�_�PB ��'%xRWh���e}��w��X�ə*J�Q7�j+#�1Q"���E/n3L�r�~��(>�,^�"O <r�b�?��cN2}�8��[�sA����+k2��\�8�YҐ	��~��@�D@�|��u	T�IU���|L��Ms���<��ˊ��U��F�5КkvП=5Ǩ���-�a���ow���I�@нr���\��.C��JxNV��IO�,�{�F�\��kR�[$t�c[��ܘ:^�� ߐ5��nV��m�H�p�m�:��y!o�k*y��P����P��U
���܂��BQ���,�O�/a������2B��1�f��oĜe7�拙���{� &���"�G1����E0Ja�>��񻺼�\�z�aA�=a��2Oq��VG��6�H���c�1��`^��uKr��Q�p�Fj>�ZJ.�~�:�4F�eV7�^�q��M�j�����V���]����W�[S Zc�S��9ײ�?���o��1�����Q� Z��]9��ܪo;3!;�qE�a��P����X��}�޺]P�MF�UR9蔕4�)��NG���SI��fP G�a��BĕxP<5��o��lH���7�!6�)S�]����AY����+���qF��4+^H��?����B� ��8�\��&➆B+���-ks$)߄�_�=�ګ����L��Y���diΟ�\��-�k����F�]��l��kz��
��زɏZx��+�������F~q��9��Qa�h�]-=�o���9�}�K��
�ԵgV�N1f��W��A�\ӇLO��E`w��$���HC�]eS���Q^E��Z�Q��)Y;��ĂQ�8�O8�W�X[ЮT�?�m�����L��/Q��/B��JQL�@��r��Y����������f�A�B�6T�B�����L(�!�Om,=��`�	;W(p_������Ϗ�̽�����	�Y�l�|���c��X�>�[�5y0p�i�Q������p��\ك�l봌�����hm0�ذ0�9�j;6X��a�o�;joXke�iX��+���W�Γ"b�/KؚtTn�"�����$7�a��R/�@� �0���#��q�� DF��I��G�һ���fq�b�$l4f�\���fMc"��[M<���nĜy���uKh��@�^8�X˕
��W��T�~��O�F#��T��Am>� ޕ^�����D�,�`~:�Yf�׾WR;�ɸ�p���lp�~ C�B�d\�I�Z�ۛ����$ u�@�����`~=,	�	ǜ M�6\d�E4�5w�!��߮+ �|�*���C�η�8�H�j���Q�͇�P�`�Kܜv�N{y���N�M�R\Ѷ"��p�e*uk�oL&d��?}������l��������c�CeX� �g�����IN�5'AͰ��A:�(%u8��Rog7�F`疺j;�ġ����} ���d���W4�Wl�rNn�fUPҭ��G*��L"�� b�Fgic���d*O,��X����)��ca������,�-�;T��a7�ȆF��9ȡ����N� g��14b����x�6�����U������M��)J̣����i�9�2ë���kޛ�/��U �� t�fS���*i{��6F��C��Ha�4w�~�EZ�{�����{�xy���ٕ��%9g:^j�<�hڧ���.)G\��f<j9�JK�O��� �§��)z���Ue<��1�]����]���d���u��!�c�}펓�:S7��~��NdUݪ�F�������5b�����`�N��K��{?x� {O�F�#(���I����|�vv���ɬ�u���Z���8�P�t��(q����b�T����%�_���Ԝ�����O ���(�T���=�l���/h�EL�A/��2���UOd��]#��1lz(h�����@��*����~'���;&|��vE1��b-}���p�Y#[E�w�����i��.�+�1������'�o�ur�SL�M��������D��\E��|��(�T�-^�g�C�s����k�8R�"����m`Si�D�MM1���TS�W\(T��R����n��{Ǘ���%D���g� �n�� v��ٝ�UdB��U!���rD	�,ݫ6���q:�!��]Ľ�x�G.F����j^�RI/к��_p$ɾ响 ��s�<4+��ܣ���z��w�Ŭ��OVO��FuT�kO�ԝۍ=[���nk��Aj~�h쉪�!��\���1'������PS�o�d1�o�W�����6�����X�EW�<a�#J��C��MM�H�n;����j%�{$�01�2���3��g�Ի�����jwI�\1׻kd���.r?co�d��_J�^ў�����0��q���C��3+�{Az`�	�/(C4�9��,�b$SBK%�4-�<�� z�����9���&r��'�A]-��f�hpง��ś�Fo�s�)���R�`�{i!}r�(q���~q����ܛ�iN