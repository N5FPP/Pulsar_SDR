��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��e�ik3�������w$����g|��J^]ؽ�2h ^A ñ9���s�x�PJwBE��FI4FoF�H�TS8��;7}����v	nv��Ԟl���=��1B��8���Z�m�y�WL�߭���O'�_�).O�Սۖ��C ��D`E����97K����C�FWHٚT/j�TҐ�mӇb,�q	�>-���L?dխ�Z��U���L�$��]Kt\A_��
1�2�z�G�~ ��Ru`1՘�^#�>c��p�I���	�c�(L�c���J![*�����Õ�{B�}�hu�ⴓ�긮��ak��C� �|38a%Q�O��چ�X���˲���C�6�-��̢����v���R���AG(��km�DMbէ�^ao�0��b�R�#��J�X��Q��+L!��/�4��!?(V2�mM}�N��"��5M�ء�<�����d��}ݼ��c/T0!м��pv�y}b�R$��pAM�WI��!H̭�t� P`�n�zӮC�t@eI����s�+��\��������Ż+�� 9�z�����vm�b��.�c���m��- {��Q�Iyq;����a,7�L�"fx�e7��r^���]��GV���21V���w`�Y�m#KI�a�ݹ��ׯC�NN��n}`�y��WV�扼���46�<��'��}0���+7�Yȩ�OYi�O�!��댙���9�nG"�r���$�p��1��+G�&C��������7'�F����}ƅQ�E��fN2x�-�x*�t��fo�Q��B��e�:q4�mK�
�V���(��OL��ǔ�+Y�c ��Ϲ���Jq�z7FT
�<�=  1��w���b,	E�s��5�?��oxN�v��~k���� S�R��'������[�u����|x-mt��	��]����ӆ>'_�3��%|h�]ɧ����a�ݤ�
G�[�V��N��+��0]�xP�M�v�"W��v��̧�+���s�x���Mm�*]Y*�Ҡ#�n�A�S.A�	�A��l|�h����z]�$o`�xÎm��I����#Ce*�=ʼjos�^�"��T��%O�>O��25=w�����P2���z��J���T۝5B�kD`'a����}�������\ߧ���4Qo�$���:��C~����tV�H�d���L��3X����X���.�g�\1
@��;?~��ރM���B�|ސ��$��-w�i���*ٱ���ap�CC���o�K5�$��� ;&2��� L�aI�����	�O��_#��KF�qn�� ˛��EU�Ų������ֆC���]? c�GR��I-Pbh��$9�k�#���g��P�+Ӭ(��N�o��~��Qt����
�s� 6�Y&6�J ��v 
���AY��7Q����B�|I���������%ʶajm+p��]�_ھ?��8����Z����˻��iN���Տ�+�]Pf��d�Po^)���r4�`%�{`vQg�נw@���1$�ir�Znyr��գY� ��]�҈�Re=;�;�02�TZ �z�m�ft���c�!s�D���_n��܃aJl��`�u��Y	�{���.���)�h��z�gK�'�v��c�`*�\��'��1����)z��BCk�#/���((B�=������R�7ce��VS|ۓ��Պ�.�ʬ�E�X�X���>�` ��;-�(�c�w������.Q*��P2����9�n�TC�U��/���FJfF<VMYo���5d{y23o��c5	!��L3��w����rq>�*Bd��X��?�4@fԖ̓��8H1�}�ȥK'���@i�KMU������?���*�\�ͩ�G���}��&7�@��6���#ߐ��͜T{�:X>�y"9� �����|�^�K�*��T��JU�UP	b"e8|�����L�}צ��;	�}� �A#��{��)T���B.���m�V�p�ד�������031JΠ�5�W�����FB��+;��q�b�uV�yr��$`�u1��=����/��GϷ*X5 [
��!�ҁ�
q�yh,��GF ��S48;9�t�K3�(�E�&�(ʟ��6�5Gt� 8�xD���YN	?�a/\������3b�֛^�o#:Y�8����0
�F�1|_V��\�%���d��4�݁(�H�jb�Ra� �s+�cPE �%A�?�x�= y���̅G!Z�jQ��ia�w�3�PI��`&�[�AtҾ��m��R,5׹�yGO5`�v�2U��|�@+��T��Fk��]:�L3T刾%�'�y����X��:��,pN:N�2���;�ߣ{���a�s�֜�����]Ε������lU��Vm��9���Fӛ�wҪp0@,��pH�C�0���:�ﷹ�;�L�H�����kS�EU)��u�q��,��s'���zx�{����Rdh�-C"��[v�\�k�g���
�\�N6^"�d·��DR�Nz˰���p^�\�XzꏺP�|/A��V���Y7m����*��sG�11��r���kk��u	+��B�$��X�S���*
� �l9������_�T%�X<���~\��:�e�]���A\�-�xyZ��k���U���\yz�0��߸�����c;�����v���%F��:f$�1ZV�	��$Î�\�&A�v۷�R��u�\��8��b?^�}� ��@��Y-��$E�5��?=��u7��2W&Ŕ#�f��c0�����	��=/ M�7�tp���b<
�(��=#�&	�Jf�n������)�0�i�r7�dL�Ӊ��v���7ɚ�:�7�<��c���u`���:�G�%�\fR��ĳ2�e��[��47���d��G.�3�76f$�(N�Ef/�f���	�+T��oZ���"��8�H���d�>j<&"͠A(��������Gt�.qH~����љ�k��C�u�p�RTe���|����]|��hJ���WG���c�n�{����<�O�_�FY���Tg���),#� ô#g�� =�;�<_As�}�MKa<0��rH��@80���!?�rPi辇{��?�~n�i��U#���{h&��k�!ٚ6l�D=;b��&6�V���s!�������Lq͗pД?Х�l%��E��H~�kV<�Hu�+���ó�1�X{�-N��2m���Mg�#�/8~d:��ӀY�3+a�\mC�37MϜMtU[�m�8&Q�oAl��t��Q?_�&�+�'�K8(Ok�z�S�N���r�����*ۂ���bT9=�g�YL2r�4>Lk�FN���G����v�,/m����)V0Һ��9�y� ��ʵ>�6�X��`�&�E��q��>%���[?��>"]n�` -����(ȱy�����{��\�\��9Hڅp�M�5�H��W��.�qQ�v�G�R�0S����E�x�VxQ�2��N�XwÈ�5��D��Y#���K��{���
�������6�I$�k���0"E�L�Ȥ��7!Gݾ5��N���u<�g��t���ת�U$���,�\.��o�s��۞X�W��U���-:j6������>�e���nA�ޛ��i�s\>��2`�,�ڠ�" �!?V������w�S��7=K����쌜Qc�ދ+07p4�+��o��;�
�|0���� +0ѓ�5�:�V���ˣ���]��"-�Z���>O�&��H7�&�����Axf�����x�&2��{�ӴU����ǆ2�� �#�AB:��� �a�(�G92F�gJ f�����Vtv+=!ly�@�%�j��$	����2�bi�k�(�Iy���7J�JѠPI��Mi�. Z8&OH��N�>k�|�B�'ġ$��&�]gW~*�t�m)����1��{�[��"߼��O:� �gq{r1����Ds��=J� 5H��E�p�W	JC�g�`�Y�ɹ�8�Ia?w��Z.����3̃�|JX�B�[�4���H,R�^t���M�Z��������ϙ\���Ưx4���j��I�URhu�R�$�W���oTN��|6��؈F��.n���#���_�y�ot��nRߝ����T��&�嗤�[X�2L1����N�Ј7�*�Ȅ�X_�Ȝ�x4P���@v������k��`��-U��6��.ڔ���au��ZFv�E�gAGM�4T�-�����筙��*�F�k;�/&I��uI����=���ى�MN;4)FO�cvVz8��\Xj�j�Do�f��p���y�߽��g���ج߀*х(�����h��Ut�Z�
UH�6�����4���e�9��:"W��!�b,
��1֡Q7�"�b�;"�y�ɴ�1ߙU);H��G����Ě���Z��&�r�_�8*&��^M�u{]Wr6�۪�;��Ԩ���Yס筡��ga�D�e��ߏ]7?�n<6Q%/+(:=O5�E�f��hP����YF��5f2������Θ8�K�:��/��������~�@\	�zc��S�g�����kDΓ3E�E�e6�6Яd��N?�!�F=䜬N��i�n�:hD0N���]���(�.{��A7�|�lɠ�l�8����3+���7&+�u*���K�cRN�e��n�.�����6��N�<;��Է�ܓ)�����r-��dvF>d`4"g�f�K� �I�t�;�w�c�:YT�ն�}',ħ�����}�/� �a����?�*��XI�kAg�8�-�:�5��aH@�G)Kf�jG���ݏ�G�/C���C�9��_$�I[�՚I�(x��ŵܽEh�	W�hc��mq���|�N��P���xY���u�5k�E3E����q-崰�����픛_Q"�~���D�p$�8�\`+8��,.�W~�����`���$������O�z'.N�0W�Q]ao�ަ�8�L1@7^���N���N�W?B��Q�E5��:��Ip����G̈́�Z�����bl��I�	��C�k�R~���t!��0���P�X�\��Gkw�wq&�yL���.�ؾ	`pa����;F�2�l�	�BC�������(Ĩ�z�}zAvq1�,�PZG��z�FP�Ŗ!��ѝK%-�|P���i��ժTvq��8������ P�יO�k<����d���[ ��0�
/ˣ��Q�&�̷����n3}ܻ�r	X��ѹ9C�O���X�o 2��M���9�u���nu����jG<����g�6�б	�3�$��#'�S��WL-������0�S�~Eე)��=m��M�M�����3D6)jv���h����=�k��ۡ��l& F��E7m�I�R�܎���y��c�A��$l��F�0�^q���'�I�hʸ�\5�Bjŋ"�{B�zzG�9��
��a�X���[��|U{�ug���.��Pgݸ<��:�Íǽǉ���Fh�&� ���� ��0x��P�+ǲę��)�, E����n9���wV6�܌�N��F�3+{��8�}�?j����A��2�j��V�_Sih�^*D�5#�k�R�l�z�[��f⋶:Ð,̈��K3�ed�k���v	��-+�:���BH<ݝ����� !�|4�ڝ�M��F���
�B�z2NNh���^�{��_͌�z��B�������A�y�K�P�d�R~,g���k 9ҩ�_HMt�+���Cl�6�M`X*���ܱ��K*�Eӓ�'����ٸ<��T�W|k�$�?��6�$[bExn���Q��`� ��Ʈ'y/fC`�4_=�o�HGF�� �I����6�|��/G�kCV�@Em�5���s_��D�$�r���(��Q��_�-�\�{��i�e�ȍ�yt���M�O��n~�r�ZIF�(ʑ����>^�$���>$����-�®@3m\Y�K/9��ԃ}��W�n��y��2�r]�m������?���V�T@�>�f���#=mFg@+y9���VtM�ImݼX�e*ޫW7ܯy�/2��vyV��9 �n鸞�����~YL?�څN��X>"i�W�@��<i���5k�xv�f�]�ʭ��3B��Hp�շ'I�Yz�K�D��c eui�q�
EJ��]Y"�D\���[��Qh�{��͓���1�\ ���՛�.(p((�9�̽�H��qE��]��.�G�$4�i4#�'� z����˷SLtW.��9^�Ȁ5BҪ
H�I��PN�����uB���/���*�I���>[��}_QV�����:��7�坾�� �(�����gpG�G�����r�K_�׋I�\�du���&�u�,T���T��)�o�����o
7��Jn�����ǉ�l� r�3h?}ڂ�	k�	?Kj@TH1�g�.�9ݿ/-�s����1����8���ࣞ/vLMf������8y�U57<����^���6�|�#H�s�I4YV������ <2��J�tû�=Pr(��d�Ә:V�wD�/�v:�i8[��c�ZS�Dh� ;QK�*������h/>K5^��F��~�r@2��'6=SC����c$D |��+A�F�T�G��^uC:�����{Fpe�ʠ~҂2_��k�e���rh9�b \l|��[�X��V3#	�
R.��d�9�>�=@�QqN
k�7�P�;V��9�k���)���/�0�V�9
�E����Y���'FY��ނ��p΍1����KK�dJ�E�ڈe��;�5�*�~�����%�iq"���#M�$w�����,ǳBYm�
��7���c�^�����y�{�#@�l+/��� �՟skϚAY���.Y��0�+إVJ»�Pʷ2��G��[ɨ.oi4�č�{��J�b�MOzP��iɉ,�<���W�x��2���T�K���^�"K�; �.}��؞.���8
���eCpk!�7�#T��Ru��S�q C����4 ��ś��ӓK����h��]$��)^ �*��f�e�5�W�	Cu��� �V Jŝ�U&˙��lM{}��%N�����{�������Hc���;���}�v�{Ө�~ U<*���
k&A�Vy���1)?q
�J�=AlZ>��,v�O%<	ė:��(��؍E�z�L<��!���=�������#�T`)����T��뭉���5�;H���=�	E@:;�""�� 6ulԐB�5�0@�L�gM���W1:�Œ�r�S��B!���=0���O�`���ʖQ�Q`���Psz����R���;œ�Ѡ�8R����� )3��貘[�/�*lb�" ����~y����T�߅�}�e�K������Lk���RƮ�w,q� %^�������w���	o�υ�������eZ�v�Z/iJ�͈P�C�<�'�%��>P�����I�� ^�|f�7(���I��TE���-��g2qIח/���L��H�?d�>��>��/����"�?�#��$Tl��ԍ$������՘,r��Ne�j������Ķ'k�`�yK�.}}�����6��|�2|ge+��+���W�r�;�0�t���AҤ�/G��7\����F}:�d~ʰ.����]�N.x���J���us��f�����2n9O@`��`(�ʱlGGż˰�c|U�(,Ҋf����NpJ�N��fS;��m�#ѾSI=�D��l�"����Ž�9��1i�$\����!L���d#�#�����<����sO�=�߭�r�Z4#p��~Wi���.���idkb�~p�t�ָ��M*l^�.��Q�f��N��
�\�$Q��zV�tU��J`���� ����?�v�a��0)P5��i�^�<t:�I��=���3�Ue��5ԉ�U�Pv�q@Y�l�^��6����Xa�.#��w)g\@�fW�ٓ��l�:�F�:n��tC�����n Y`��2�%n�`o6���&W;�)aJ��+�4�񾹜|{�}H�C���ji��䤠$4錄֡�}��b���s���'�eG��)̗�yM4&����������F�\�[�:�=J�y& �Y�E&�H��P�����Y�숯�[�����o�ע�X�	Q"��\p�s^�3׵3d�3`��{�X�؃���~�ʓO���?O	�%���7����Y���8W�Ĺؗ�Wi����b̱q�U"v�g��Prʩ��4�,,�~Ä^Rn��s���Q/�Y���&6S�-�C*_��P+ b��ߙ�]'��:/�U>+�����@��8i��ۓj�	D��O�Ս◐�����e����p���cIH�qi�a����n�ɘY���?�ՍX�>X�>��U7SQ�%C;n'0�kq"�;m��X�t9z�ɨ�n�i�吠�$n�P��UQ��1=�.)4,���JNN?��o�b�������iT��f�j|���=�T����c]�������q}��I��6ۍ�x������<uC���Tt��o�T�rx������k(�ho�"��j���K��`1	��c(1j> O(`!G��}i�����Og�r2����~m�BE�(58Ӥ!�e��X�ܭPH8Q����)�mI�ߒ"����i[v=�f�|	��ߢ��%��j��R6c�5t8��Mߒ\�Y�����)?�-F]��y���0�G���s�J��v�F�x *�t<��
�~�d��V�g�$�k@�9�'ZV��cb��0P����뵙V��;1=H�2���:�9��U�����ݨ��KN�)�����>޾�3��<W��:��ʡ@���Ɏ8������YzTV���LS�#'0��~n ��[U���W��+��O��hf#�h��*:Kd�O���~�!�ׯ��UR�]+��#"� &įU[ ��1⪉i?=���&��@} ��иww�nj��:��l h}�j����)��߾�5׽+,��9��1=�m3͜�{�xq8�L���U��1X��O�B7Ke��%)����`�i�ͩ,�qH���>��maQ)�T���]�#.�W�y���s��i�:����q�|���o6�M� ׂ:��J��8�}���Kz6�v��
$0���L����ƮTϓ3
�&��y��Ҟ:gufN��T<���M`�#�"Nϡ��t~��[�x���x&���J��8�J�-��tɒ���?����m����B$|�t!r�t���p��N�.jk�袙B��D�(Wu�7t����+�aph�5h���L����xnEζ;�q���.��iu;�_ %m���8o �}2[����t�����o#��p�s��X7CMca)�燊���mr[�Gb1�+G��&��l����S�W�V�� .G�L�1衊b���t^w��dYg,�.wW'�Sr����,/9u��5��F?.�~S`m("�a����Qr�
���}�׭W�3L�!v�0
�U�s2�D��� 5��ͷ�^ {�K�u&�j��&W0o�u+�r� :�sی.(�H�'�W����=�5<���fن���|�&����scGs��cZ(�|�������0��[]��S��]o�򏦮-�4��(��m�#������uUyCٹlPe�3:���1� '�#�`�)(=Ñ)�M0�0.;�P#V{ ʸ��s�3��n�&�O@�bݓΨ1�EF�����;����A���o;�w_����W����!�o��5�mU�fN�.����*�U����3��E�[*ՠ7�	�eVY���.�`q\�}@�i'�>�2hi��4��Sş�� -��︋�$���i��j4)f^9�:0�q h����&K�%��9�%�Z�4���'_�����:��ԛY���V�!�����k��a܇���@��Х��J��0	�`���H���u6zI$�a�6]v��ɘ k�4'�d���]�/.�5�����%�l"��A��	?f&*	�ˡ��i!��
�`�c��R���$�R,)������~ss��(�W��Q��(�Sw�U���[�|��{��۞-q T�<�ASr"]�C���Nrg68�<�4� �+��3�R��s��{������$�|g�i��Q��ȷW��4����x2�,'j�/�_i?��/��V	�L����C�
8�ނ�C;$����Wl���N�VϺB�-�����(͑�	�]Əy:�,�v�E���\����դ-z�qXZ�I��XC.$����w*I ���6��Nv�Ҟ�C���'5��nݳ�uv�s�&V��O,��@w��D��k�vRs'98�PJ���Y�q���⅚�g��clwQE>4R!s�8�� j���Nm|R�ڨ&w�9?m/�N�!��Y�k<ʽ�/�֙<��`G���QW�կlL�$�r�����9Ӵ�'^�[
�|V�
a�ߡ D� ����PE��#�� ��ˌ���x��`rL�CWOѳ�i:�a�;����2;5~��ޝ�s�AC���^l���U��c�{$��}�I�ệd7o�|z������>���,����<��2=�m��y��B�D�o��,����,���ٌv�����q��(�~�?3�^"�s����L�����3�G��$W��lO 8�K��d�w��tQ��%m)�/����E`�h�k���l��R�I�Q/X��xRMJ/?�Y�I��j�������R�"�BFh-��gY/�7X$o���������s��n@���xb��l��Sh:����tᆘċ/����g�
�,�J�z�Y�5'sQ��h��8�����i4Ar$?Ȓ��2�;���%�Qx�� �bA˦Jҭ�Xi�q�&,���st�V2p����q���l�ZE ��Cz�BI��]m�7�qpc^�����k��v4��Y�_L�<y��]�(o��݋`��cz��W_)�����Q�����?t��x���D�@3i��w���v$>TS�f)��M�О}tCb�fi����l�	�����M&q$)-����M)k���h�<ڸ���jZ$������B�IF}Ζg2UtQsN���|���Rd �1���A،dvSB��]sE��|MpӮ���,�a�ձe���0	��ƅ�S�� �k�����cj�����69����5c�.Ҋ�ᇴ��BV�����U��V;k�Ҹ���<���Cp�����Y'����UL��+��Uǡٌ�+im�g���ؓ��/�a�R"#�JW��G`���5J~���*��:��>�#zٸ$�_tG�<I>��)t�)P�G�QY�r�y�6{I��l2t�6.D�gDrq�k\s�Il{�M;B:s�w.\���WT�@���k�C��^Pt�%	cG�����@	;��xq�hGfc|�Vb'X�x��1Ą�������L��E~��k�1� @5\A$x�Q���a�g	�P�zȐ�.sp�s�cf">�4q�H�[��b䑐/߁`��4�`�ꖶNl�K���f�@X8DH��{����L�2���_����>�2��0[������ι{&��7��{�e�mg�&6Q�����7�	����F�uP�����k�srk3u�n�_�H�[Y����m�u���8��!sp+\j
fN��쌚2iA�^���Z�t�D�>J��I,Q)vדw��]�"(��Jg��d.�����z�d�v4���ፅJ��(����Y��`��p%S<�����:��R�K�K�"_�y�������J�!Ȕ"���8[���B����� *��#D��j�yo\F��p�M�*�_�A�^�;����Z��{�g*
��%�!����d�&�˃��ƍq�mrS@ۨub�t���3�J��w���q�f"v�:���_�`��^^]i�g��<�^Lw�I��QiN�V^�ly������$�eMF�*�^���������B���Г���9�#D�S��s��אK%���֓�S ��W��Fg㾏s�-ݟ;k��d�� l�� ��MSr��lȑU��>�������#;�ѥ]�\�'ӑdv�N���] ����-�_�]%�h��Ӫ�#�FWY�e�Ug>m�M	��J&�ęRa��Ѯ����
>cO�;̛:�*[j�(�^A&�=]�!�i���ņ�Njr���VUOJ��L�JgM����: �^E��t��B)��΄�WI�r|Hi���3�����6�##x��$H��	� א��$�-��c�.���6c\���JY�_Vh!~|��*�3K�nO��M�yc	�;�4h$;yK����!#K,�be�#���-ߎ	1��q�z�B�Wt�z���g���N���RLf���O*�:?!�G�r��k��
.��P*�xkߓ�}�X.���Y��i��[�3�]�=e՞MǷ��FO�֤��ƭs�ЄO�M܎b�����}��x�^��0	�� ;���M��̝I��SLf�Py���%?Յ�+su�Mg^����lS�����!&�8'IEX���cJ���0T�fm��ú�Q Rlv�j��3��;M!�WP�?R3�+�M3i�#*ʍ�@�p�|{Z#�[m��H:P�飫7�^�]NAq��+�5fp��[C*��vI �UӖ�rc��֒���Ck��.w�&<���X��+L��~ ���~("�wo���T� �W��r�����u�E�J�P�����m�E�`�w` ��3��i28��ߤ[Jc("��f|G<��;��d�օ����z�a���#ND�ܩN�f���`24ν�Rt��o��`/)�Jg�./7}<��3k̣TE�*�ޯ�:?䱁J��yg�����nX����D@yY��О�P�o�8� �]�,���H>��v�q?s	p����FQ�k���1Y���Z��50�\x4NS{�WYaN�Dr2��~�b����eq���Yɴy�F��c��
{�#7��&��F��+��64k·�wTk��F�������(�ܩم�\b�'����Ֆgk�O�<�:�a}��� �$,�*s�7�g�y�NbH�#J���Ȏ��^FE�d�SO�з�DE���<��*p{-�Qi{|�2i�����ȸ���+2�xh^]~=��k�1�F��:��=P��/f�v+�X�x����L�Y�m��b>X%"������Y�f�>g�vpnĿ��T���"w�ަ�$��� g#����"f�5��5g[���y�P{�ͩl�h"��m��'J>\ ��@Dk�Zp�\K`��6��E�t��od�g�ع���#l��\@D�in D�;�p���uW�iP�a���¢JYj�U��%�rMaݎv]*��hHdi)����t�}>Y�,�ѕ��'�L�����R�C�Ƙ}Z�X�a��c_\;qwmE�8�UV:5��G^eDT������3D�mǅ��G� Kp̲����hG-�,�3~D�2&Fm�m�(&���I�If����}ߑ�4З��'���@EG/>�d󪳨�����AԔ���+U���]���{���[�3�IP�H 
�R3�fI� �;�Yb������*#L�����c�Bp��Gu����U^z�7���#i�X�{���:j�?���O^`�]jt��H��o�(@�*E���+���oH=R�u�,(A����!��U@=p��r�<��K�W��1/�N.�t!�;� 0캟�	������B6�uȑ ��iY�5 	w��ƭE�5[�/�+��
N��N@=toϴ������m��3V7*9h�����q+�{��r�譿8��Y�(q�_� N��K ���|��;�x�_2.�k�`rv��v99�Љ���-������8���������y��d&��L/TZ�O�E2������3��!���,�Y�$^������z����V�ǻ��<�N�[�lv�a����@zS��5o�܉:9F˸��T�4:�uݹആ��ǜ����؋�����귙�Խ�Y�pŚ'A;��l`A���U��<_:���>^�1�*^r.��K����S��Oc�O�5 �(?�W�BD8��*ln�\�"Qp�$ᅇ'���o�����m^?-����ņ6>�;��>�PGf�5����%ɬ���{���E�i�aO�ҁNU��O9�M*����s[>iѸ]�o�4O!^/{����\�U�|������C{5"�4�C.=t����d�F;��-F�/�XM#1�������¶{gG)X�g�{>�_�Ӫ!�H�Rru��=9ӈ�������݇$�%' i��p�uУ�"s� MK�bU�g�2��a�T��O���qg���mک{�ZD��c�[~����(�G�j��n������\}�x�	��&���������@��2.����
�0����%��,�����ص���8�����V�(qcg;y����P��;;�儎1������C�n���cu��	�WZ˙Vb<��������H?(t?���Ď�nn���ɕ	N$��w/-#�㓾7���X:&\	�R�(�0�n�=M��s2�K��?�e��m�,�DY�!8T��<��_��~��2���
�V@��l��vԺш)��`�v��4�� �G����:c�p�1M�}�oFx��蘉Y\��sl!�`�f��J���m�a.�W�m�8���5x�ES��P6E�Bǀ�����ο��E���\�0S��,O���X�2�i�Vgfaf�.@��4�'�E~qx�����F���� C��g��,?����B�m�Κr>�����D��q[�6��0F����6f^�R���KO�<I������
��7�1�em�ԀJ�M_�Z�ȋ�ɇYl�p�ϫA�5*��$�6��L��m�K=%>1/h��h�Z~<�9�_h�\M�s4�@m=7�B���޸�9��'��^Y�~�����̞���,فu?�5���B��SB,h��Ju�G���TҢ��tq�G>X.4b�:����c�|��H�S�ǐ�6�׍B�&�Uy@���y�����[P��;��Z�چH<d�;�`1���Z��sff	��x�M���A*�g.z<����q6��7������v�+��H������D~+1���~>,!'���F�̱H� �^cXhg4r7ۃ��FG�
���49�)�|	���C�}���!]Џ���*�k�����T�J" ������U4�h!$b�fG����Y�c��l1����uWհ�^��m�b�d����km\�!s}��0�YY���ڲ@���]��A���􆱩�wch�J��I�!��Q*Uk߽�A1����E5I�ZjlG�Y1��Q��)Y6�]�'�ZR���]�~�a��X�ڝr��ɻ|Ed�V��X��V��9�S
-�Q���,mؗE�	�]�w�P��ʜXJ��]�s~�Ͷ����S+bgb�g�� ��r�v��rl��L	d�J.�P�d�u�=�&���KOO���m"#�YnlA��������f3�%�Q�M�k�b�C���%��C�>](�=���*�e2�Pb?&s�D�^���*��/�-MEZ�~�����d����q���!�nz�"���إ�q����qf�H	>�CIϠ�P���VP�l{����֫��L6T�Mi$6�ʞ{5�� [�N�J�
��xQ��c�ඇ�ԉX#���ZF�D�����!�TW�86~�B��n�J%�QCm@N������Er}�6�m��~?������ФaۈI�E��N'�Y��t ��������ҡ�F�ָ��3��W��\+�q�=w���}ip��☦D�ٴ򞀚����|���������3�l�d_'��F털��m_��Z�R��H	��?����ܥ��6�<���AL<�Uw�t3��X��? �¹�o���k� ]����V����f�u�;��v�8E�@
?ɀ9�n��A�\M ظ&�%�8I����}�g��Et�P����cy�sc�X�ub�=�V:_T%�!��!���Pi�(�RtY�ʡ[g>���5Ѭ�NG�%yp��+`����i���߾K[��o�S��\w�̴����r�3<��Y�+�c�*�v��x�Z��:q��5=�N��6�\��'S�k
:��
��~T���Z�S���26�2��`&�}����@c����D��q�+ؓ�ڒ�N���Ǐ>��Ծ��B��<���+�2�Ox��_=���8#*��V��@J���/_���n�To�fi̧Iv�4V��1�銠��G��@�\�,Ȓ��+���K���:̠���c�]W��<��=�d�)^3J����
��;��^T�;7W�c�:+kǜ�'�v
wbM.GL��6��0�A&*ͳ����
�~��y�}���-���Lv���)�[Y�%����Q�.�x>C�Tݻu_�ˍ�;�.2��m�'���pL,�d4��dH5�vdX�>#���d�p�٤�pЫw���,�_+r��^i�D7D�x,AUR@G`�ch�,)iR�CÓ���@_*�՚3�����0�6��I��QSX"!q�v8+������B_ �-� 蟂ӻ�
�儞���I��,�L���Ӷ�%|���eB�P��
J���ثe�'U#�4�����l ����M�P�@~x��*x�o�,w���`�!zH�|��0�AlX��ˎ�@[�ò/�\��d����5'�tiS�?�n*2��C�������ɱ��:��6�zҽdB$XH�c������v�g^T@nQ����F���F���W���ND^��ڎ�'y��Ŏ�{2��-��]��t�}��BE>L�
�uujvZ��R�	�^��3�CR���lm�=�焒��o��_6��)�F��Y��ʹiΥUtcr�G���F�1�h���M=F94��)�{<CB�	I���`�N��3�%/x���uu���ef�4���O2��ƹ
8|ؾ�#RRa�T���o�0�z�Z�+�(nv��јUI��٥a��wT�Ӌ�@��:�9v�4�����	�{�p����ո���-�'��4�m��H�6�4����QrZ+�Ճ<i��x�Sp�_q�,˗M�Toc�����~��Xi���`�2J����)q�ECyd	c�&JA���\���o?�`!�a� �X�[�f����d�7����y�|��d}�����]�֕gD�]��ݬ}"���28�(�ҷ��j�u$�T|�6�p��_�G�U#H�N��D�j�&&�e���,��b�[qb�e>�:DG^ 6����`0�9��i�:�`���i�^�y8�v�+(b���������F!���d����ocU엓h�\���;��N"������}�)5�/$��8O,ej�O��X���[#�D��J��q�XZ�3�B�������N� Dr�Lm���E�Q�	"&��0mh~j'Irm�>�o�3}�9�4�ϝ����_�����ǈ���Fx�bo��lT�0_��r�T�(ôjL���G8��H,�t_�N��D�s�������ͷdUr®.>���&������z���hiB��e�e�D>	����*�"�����U�٬�1�O/��z�"�f�\q��} �<�p�6������ꂋәV���7���Z&'jx������JAh D���u*���"[�Q������~U�pL��.�Z��	�,��>*�!���^���ƻ�����N�C-Z����,��GUM��3���=�JXj�|�a���|,p��O��Xy:�����*Tb	��7Y)sv.q�t�� ��&��vz��[t?&%�(��ŰF����>w=�;��;���k�����|�0ϓ3��#ۃ�H��8��p�(:�}x��G�'x}�N9�7����j�/f3��[!��ZD-):�*�S�������'7�H�����x���6%�'��?Jhͭ���D������J�e�w8�_{�~$��@�q5�>QȦw%�Vo��)�&�iP�����K���RW��[2q��}W��2.�~�ͺ�%��IxᴹBEZg���w|C	Ƞ�<Ps����k�lF~�9-��WC��������2�*���Z�����x��2��N͸���Ƿ�0uQ^��u���S]��Z[T]�~D�ʮ誠�}��8/��~�ͧ6���}���n�ۖ����hV�5U:~΋f$^0�8~&*�H�,��E��4��1_��0�l�r=Ċ�H�#$�"��q�EU�Z�(�S�W���	s��S5�ą��,yxo�;-eL�3�=�=����b�<�X��{�b���f]X���>�=�IS�<���H�r�a;*r^l�ȃ��k3�$ f�J�r���A3�6a� �bǪ(Nw��Xqg֨��M4� ���9�y���t�N��v�O����}��Z9�XW��Mc���P�a���F0'G�sT,w��lȦ�w{�@������J�;g+��(��DH�J��Z��r�dyk��+t�p��TWhY�R����bdV����@_m��R����YM�\�2?!�X��_�䞎��E1� ��{�e�*`t�  q��v�=�DxS���G8���r���D�'�&�u�]�e�P��ɒ�z�,|�W/�P�j>Hm�[�<O���ur�z"��&�M׉}v��-��l^(���QjV4�� ���	���X�u���%���C���a������ȫ���ĺ��x{��r ]�����2����s_S�$|O��R�،��Y�T���%nG��fܠq�u��z��=�k��Ntm��4^q�F�3@\
Dt|��v/������~�/ע��Yi�nZ�TLv�	����HB�G����p��-a� i��K-�,�>��(_�o5��%��#纙[t�����+�q���B~��,p�k�-��0��.}
NG�<�S�8��f|$㕚{OE���xD�N􀡜������H��WnZc*en��(Rb��9,�=��Bg����:ZG�V%��l���W�Ұ�������������/���}rЉ��A������u?�8di/�lx��
�i�[ 39���U8�~78���DuQO+�_X:��0e0�Ӂ7"
��C�8�^Գ��[��l ���w���/7�#B��h���u5