��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4d��oc���_LG����*k����۾�T>x�/>:��e�=�C5!)f���86�$����ԤE���oZ�&�x���� ]1����V'���Hci������I���-�;����{�gr�HR�l�q����~�n�2�����̴S�c�6�'o����f�?L�2���r�����uq/�Z��a['R�)9"+",��:�l/
����#���U\3�$π��`3��J�,�;K��=.�ʄ1���c��ą�&Y+[&��z{��/j��?|��~:�%��?�!M1�3?ߤ�	d���j"VlVg8��j&84)�|K�\�Y��m���TU-�^V <h�Τ�4XU�/6�����X�_A����W!��i��o��>��B��.��9C��iżׇ�2�%>+o��q�(t�
�%�\����·�*,U��y�oxmX S�`���;�F�S7�
�(���!�e�5�I��Ey·���e�`
&NTv��n�������Րae�m�d�9�<]����kw/��׼3`����ǧ=��ό����d%;�4�����"?E����R�m%���<�:F�Z�䕼jp�j7���P�U����AX�����:;��}1I>�[Z�洽��J�(T��(A���ik�sO����al�	�y�7�Ady�3� Ck�ѐ�9���#O�XM��@ŏ��X@���6�-i�� �*D�ӆZ-sa)K�7�
�3�`8�"\��u������Axw|*�>�y�Z��eDJ��rs�?���P�ι��Q \�f�Q)hQ�&��c�'��n.l�.'I�X	�D)!���s_��@U[%�Q�A���"��L��֢��۾����KJϽ�U ��T�/�f�MYA�����������=��D����e��|E��T��_%�����̸;�[�T�J������i���~��9׾$T�r�j?źR�o��*��C.�������uׇ<V�6�ĳ��Č�z<\�^?�����h�%X7�mp�Y^}Oa�V���_�L��������|fMX���M�T�B>�W�~l�z�S��v\���	w���՘�SF�n�:� vX������?�xS��3�!�}� Ŧx-R��&����5�s�+r�i��4(�01���mw0� #:�B�Yx_�=`S��f�$����O���J�~�:O�au���tܟ]�%;3
K20��i8��Q���kV�j��d�ԭ�����J���w���}@ɦҙ��v���`-����׌"}��J���6̀ڽ�>�'�z��Ǝ�xF�R*e��?�/�dt����n=n���/�7
�RB6�,-N('��_Z�~V�e��fd�yB4,���	#��-�ز,FF��f��C�$H�����]���.���Q���a�n�v/sB�|r9t��=)�>]�F��Q.��ɵ����������K���Z�]6^���d�����������iB=%�=�t���s�j��L�\��i�0^*�x4I�̵x�@����?�P�*����0v�����4�yO�xX%g�li���E`Yt��{�S��+�@K���%�8�|v�w���IT?P�&��ķ��L(G���T�2�����v���d��P��2wN��$3x�
ں�%�dU�#�߰�e>a��y�LW�>�W�������A��4�\v��L
�Q��n�vj�>A6�N�0F0��@v8%����R�����מ�G�&�˵�h��p�U:FD��-�<��D�ʉ���?=�6��� 6�51�	y�f-�����1`���Wh��i+H��S�8V�b�Q0�N��0�أY��?�x���cP@Z��a��Κ�A8�#�Е�;هf�Κ�>n�|�&+Rٞ���-!�}�fP�Z-����2p3�0����ٸeVQ�ԗ���<셬��%Zȇ�op=#]�%Tf=�J ��`��9��!<�맥����P�-�YXͨj��O+3�D��A��,�1(�K=_q_?�1:|��a�E�Q��vQzS`b�l�%��B�i�[-�@�X���d��x�d�a���[����;Y��]����h�B��O��R���|<�� ��� ��Dm��s��F82����������Y+*MGN(O,���y��a�)>v���:[3i�����*�c7�,������-mwf6�)+Z�i0��V���R����褐�����Z�u>Z����-��qH�eY�����]N���#���'��z(���0~���o�(�罄�
B1��!	4(g��v�%���|�Rc9�wt~����N��ndg5����6��������\`��:�� ҹD��4���ы7�W�����_6F�U9�,�oLORP��0u3��˟����&���4H�>?F�Wa��N���W̍U9�zS�vZ��P��!�t�>�w�ױ������ll�gI�À�eW`s(�
�﮴��c?&�aA����~�Kaxwd��{�^U���:a�}>tLK"s�;'k���|<�#%�51���b�o���7n�Z	������{(��Qn/�S_�Q\���U(~��썌wz�A��z	:��B���1�	��糲h[��3�h	������K�YQ�.��C_�M��/���ũQ���nJ&}���P^� "��l\���v�k������:�bQP�Q�����@���(Z�w+�Gs"&L�_p��i��󱪶j�������;G 4��2��]�k��;ތ���!u`+�kSt�,�_ܰ�^�ĩl�h���ei��>��BH�ג��1PE1�nx�	�Nm �G�z����5� v-��ᾪﻋ�[�L�W/_�	�������A!*��cyX_��pnbR`�n��
,���DH�����>���_��?-;���cg��@���`w~T5W���xn�h1X��
��γv�W�֮��_]g*�	X-�l����p���P�~�� (4Q�-���4ā�PU� Ã�v\4�O��~�@�wn�~���{*	����'mc%��:�����ac���jkgpނg��8������K�^LqX��8���+$Ԓ�$��b�[�Fd�s �@=#߼�f]�������TF�֞�+���O���gtH����qa���4�s䳩""�E 5�r�o���YǙ�T��~�:(0�p���Ӝ�žA�K<�}�>Og�����`4��q\ Y�l�;,t4#F<JjF~�=�,���~�	<^r��^���bt"y��R��w~�4C�üͬ�x^""-C����6-Z,D�SK���)��}T@N!����w��u����ld���iۑ��K�Rd�6\�:�mn_�B����5{�q�a�q���'����j���vD!��,{k%�����}'�J���̟�E��F��gD�_ե7�fP�;����rk��ɸ�Ba��+A�#Y2��4�ąW���Ba~��_?��1��d��f��/"�S�K	�����%"��蚠v��Uc�&�_]�C�/��0DuR&��~�`������ׄL#
�>Q��YL�N1Rri~V�{E�L�E%Ǿ���9�*K��~�&�pQ��K"k#:�Ir��,���Eq�3�(����jZ��I}�Q���}Ps�4�	���9��aZ���fhd��۠�������m^FK��u ����8�r��(�9�N�,��Kk�J6Y��xvW�Qn}\���y�ͻBLC����A`�@�ϧ�o?l��~��pa$R���b�#�!�χk�ԳJv��~߾7aپ5�if[�΅�Y�rjQ�Bc�G�63+�-���+�NU�b7���,��~�ֈ1�@Tz��-x�pn�8��KC���'�������	���8YB�8�Sʹ9���-Jj���
X
~�Ԭ��/Eq��?#m��?�ļ�z	�|=�L-�H�<�e�\��/@��ۓˤ��M�>��a��=~���o�	TC�ޥ#�z�j�"�u������ڴ���3??4a;�qX�Z�P=����y�0$�������"�*�h�@�놮��ן�f��B+�.�n6��m]�yƿ��;d�Vl���Ovzχ������cȷ� W]����'��+OJ&�
4l��/�<�Ы�(U��ƜI�n~�#`%�ʹ[h�wVMr,I��ˬ)I#�m�n��mc�� �cg)c|SG3O͙5C>���Y�@�s�������xf��B��N�w�6~*^��q�8m��-u0=�mp���D���)�ʰ��Q���:��y-s��l�D&�g",�ڽ��e�J ��%��m0߸�8J��z�E�u���Ĉsz��+�L�eh2�5,w�@A\YOn�[Eh�+R�F��e��-v��x�#B����\��� �Z�o24����r�L2D�m��'����Մ������_������p�r�b�$��� �3FʽC���PdvIOҥ�������lwiL��P���@y���T�o��S��F�sg�	�;�Ӹ�h$F/�'����W7>����௱�>�Rt?���_��Y6e9ǥ#��eI 9�R7�ԭʲ���ũ��82�V,����i��Q�;�d��h@5n(=�/x�j߮��e�x�ƹ��~���"-��qh��v���E^��{@���K�7*��36W��U/�+�%�'B�c��l���J��i`� !�B�-'�ok1�f�	�^��W7�TA�����4�1!��BO<�dC��[�{���Dķ���/Fp\��R9�O�2@���)Nf��0�I-kk�.�V�:}e��^�ov#-���ӐF۵dM�������X�°j�K6|��k۹Փ�#�T����3�N�2#X��ɼ�ɐ'��d�w =�z=�5-�=LL��lf`{a�ԃ��B��0o������E�f\H����]
wr����|��{�N��Q�j��?�݆�Ik�}���Z�Aۗ�ʔ���qmӖ1����Wjtf"�$O��n(�p���30�U�*t��}� �3�+���m��Y?Z�J�?�@�J�]�Zy���7��EoFY�}�A*������i�ݏ����n ��[�I�O�r_���)U۴��g��-wkkf�>y&�Z��#��E�xd�-w٪>q�L�|ɕqo+�>}4`r��K�,Tz^$o;%R�8�wk:$�`�cd����ԫ��0����n���[��N�P"��HtXaa��lR�OS��'.�K3hC\��{�N��M�#k��5�uίj����cL��������24��
?x�And�M���+dw�,o3�2rC�"�����Ą�d]�j[e�u5���uY�u T�`0H�J�n�M������~"���7�Ԯ��i��j����k=h[�w��M{�`ʱ
Cn��
ԘX#6"�.�?�Τ[�P���/����^��m���d��.���C;���YS�}�`x�/7A�a�M�ݪ�&���W��%d�Y ��u8��x� �F�&��0��٪VG�	`^�)�����ѡ�׍�jG�@�}<,=�F?m ��k߷'p�[w�U>�x�{�y������+F/��WK�Ԟ>�$���ǍnnRN*�F�������rY�9�ȍ��9�C ��K�88�p��:�����6�z;#\�G���Um�+�GE�Q���1+N����ӂ�Vp~�צ�p�9��2�CG���[�<���o׶s�0k�WN� t�&�`N����WQ�ē�Q�%
'�w x]9��y-�+I�����(8-Y����A�`�,>2Pk��ͼ�������~����o�˳��2�a�$Z[f#�-�D
c�=~�Ȕ�~fv�0��