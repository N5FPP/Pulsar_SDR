��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*���D#����=�6�c�p�GCE�N��+�xh�Eaa�Ƭ�z�5>��>s(�oƤx]C��F�i�TϚo�2���E���W�۠N	Rw��#fa�E����ǁ'�iM�$r����?�W���aݒ�3��L��'�ފ�q��p��FU����vJ�k�~���l���wFpe [�29��Zq���)Rq�� �CPu�)�;��/�V�2��'cu�*�Q��펊(�Ľ�|�3ڟk}wX��r\�� ,��E��:����B�bqr����Ǚ�A�Ǆ)���Z� _̴������v!�Uy�=�y��6��5���f��>�Pyj�]��z���
�y?���H,lV���B4�b(��\f���� �~�v,��
�� wz�B��C�n�f?��RN�IY�O������G�v3����Ё�Ԣ���8E�$��ZH$[��d�H�2��*��U)���j����s��߫�fѶu�E<�F�� ]J��b���)��$-#�L�Ѳ�Y|���ׇ�������e���Ω�`�@ysҥ!x=3Pb���#@$�j(��0`+
���"9ȣN)��HX�`���Qk�S���+;3u#���f#|���	�7	���&���ǥS���;�|���+� ��3�%���N���@�?@n,�y��&'5 �(�c�+�Yhd��������ǼB��.<Y�~a"��m	/s+�	�c�e���H��)�yp�`���g�/��u_���,MD ��eD̈́�u��C�	%VI�S�B�����#�Nƌ*�nnǕ]lB�y�_�Q��9a{;z�փ1�H8W�J�ﾕ�s=!���0�p!����ܱc�g�>G�e���o��$�|eԏM>"��e�[�C>�k�D:1oo��6Ȉ����n7��E��v��F]^�!%V��j�c��fAK�<��/�l�W�F�*A_�b�/\���k�0���Х�Q��Iν5b�i�}1�m�Ɨ�:��;�T���0O��؉V��9�[��z�y��-`W�j�s[�K�& h �c����G�hP�ُ����;��4���>|�����G9��fe!�C'�Fk�-��S=Ȧ�X��z��#�~"��x�Y��sN�
��Q�[�(�i�(W�|��M�	hZC�ج�u(gf����e"4�q��tGL�4�e�xD�,3��jI�0�U���O������U�R��)�\+��%>��r�������c��x:?���<�R�Vp�QP�R����! R�t�Jԓ{`�j�=x�~ϗ�m3|���n�o�8���g4�L�*���#0�3v�ӥ"�'(�ǙGf��Z�j���� �,2Up�ބ�C�����#��tj�!d9�h���s��Y)��\jm�A�|�^.O��|.�+Q��d���VIW!ʛ��r6#�Wz��� (^P)gb	'�lU�]krO������c�v6�^�hj��%y؏z�����?�m�8�5E�b�H�v"�ܧ�sX�Ӹ)b>9���m/��q�'b�JF��"�9��H�H�%�����家���2�i�,(��w�$n�k�og�ؙcS�x�h)���.T$`����O�9�K�*�"s����c�������yY3$�4��C�
yjݺN���}0; XI\Clqm��a��6eW0��#���x���}RI�#�S$��'��&���B���Y���& x��Z��>�L�J���~:���XE|{"���bm����y�GDA���#+!�
�z��Ʉ$N��Wh# Zb� A����Y5�O=}����(�G"��P�j2����R!�����o�\G�t
�lo��dH�PC�Mv�����&6 &Â �W�'��ݾ<M�����4r���~�jB��jդ��;��j��RQw|Ow�%-co{G�O�'qb��H���uU+6�*4�;>֫�u=��KU)���fu�f���� 3�a�2��v����O�"��"WU��tJ���;w��\�0|�Xq^G��oDs�a�D�:g�"��|�0	]���i��0�~q�T�p��by*
�ױ�z���'�Tvq4x�Ch}�$�I�ƕv��{���:���H �|{�5���98���h�˭rsvC�|9���^��r���fV�&�(�U%j�Pɿ�v S�lX{Ց
��o�BB���!>έܐ:_�_@��ڪ���H>fS�A����b�pob�W�3��6x��H@8O�ߟ�-��|1�\%�E�Mܸ�j2�]2�Tgo���i5w/R c���w(<h�T�P��n�y	p�N���O�@�2�sN�;c�,�U��L����.�S,��Û�� ?h�^��������"7jJ���>�$��[��8R3ۅ�7xF�y�����腁D)�mqK��5���U�����c�[�D�D��07-qG�����b���\�[��89,�\�ldG��u����Z&�8����!���v,-�_�yQ�^ȶ^��	��ŏ;O�����������^�b�*Ұ���ʄ��ͭ���&iGQ�$�"��>�+����u�6�$���XF3g������H�qh�Y}�-s�M����\��-�[�*BH��&49�($�>y@T��VKc6��1�G�|�* ����0�쓇�ZJW���R�W$�O.�����_�ݡh�&�zI���;�$EW�3���&���-��z�Z~�QFl0���y��6/Ȕ���B��)����������T�X�{.t(L�������u�Fp�5��D�H<�Qe��=BS��.��f����K�FF�%�h0s�q:����E�C�*`m�6t}��p	P�;28$|��cڢhK����N�;�/z����fv7��i}y����E�@Y.�� z}�[/�O7�� ^�S K�I[�T=M���Q��rZ7��s�%�jHS�h1sI�ŋByI��_�0x5����S��C�6��߂�R��i(�g,�=���"c�G�l�e�߅�3�U���ٽ4�a������ڡ�Įل���X��y����Nֹ���aZ��+�ĲX�dL�0��v�i|��_�>r�"�!LCHe��D�#�5+6k�Kc�g�V8�'��]�2�ޢ��l���L0J���<%��H�;�0��9u7QA�_�V��i����k���v�a�3����N9�:*qr���=���-�t"Qz��uL��|V(�05�W�����a/`8L�;�%
o3�{=�������4� Ɩ^�J۪�Y��f��"��1��",:�·e��i���xa^��g,�����x��lR����L%���L����L���,�|�=r���<o^Ea��CxD^�qÅ�)�g9�zG������O��x9�q�l�BG�<��Sʬ}Z��1�N���2����#T[.� P@���Y=@vR���L�M�jW=�o�*�C�P�����E�(d�hJ��Α�@���ӊ�`+�5���yr��G2[�G�������X����I�H�sE
Ñs�B�(�Ao�h���bV	��`z�U.+�%X���1!����M]O6��~E�^��4�����E��At1���H���t#ᣟ	|�<���:s�e�,��h�}:�ʹ���J��,j>b��^Vee��j��U�6����1�W�W.N�(D��������sq�޸�JW!�ĩ�"S���̏ױ���1�.�;��e,�;��9�a!7�{���X�}��na'5��VO �W����{���rPPχa�f޸0�fTo�1�_�Cpo���@�����!��&���SYk�xՙňO[�;{��J�<�5QH�9:���5m�Z���]�/ʍB���jh��c�
�z��w�.����!d4H%��\i�&��X�����F�b��@�Y�|XD�J���0�c�7c�4�����v(gP���fP�]	e���W`��W�iV���t���C��y��$$�oDc#Z- FC���Il�ҝ6���Z��ܶB�����SM*�{ё�D`�tFh�/��ӂ�T�͞������|O3�5q ��h@����`:�����:l[�|76��I����y���r�\"�m� �3�(���A�BO�6��m9R�e
���h�H��j��1��m��g�̽hE�
�zYh�ҽ�s0�J4�lޱ�r{~�{i����&���+�a���J#�����I�X�9�'���h{����'­G�|$�������b���=<[Ü�L�ܔ��t����P
t��z_�Q�m�����p��ٍ���;�&��)����}V������D5���?�C4+[�Ski$�������L���~�I���i�7�A��ZZ����|~�u��ˉ��3����q�݇��#�~�fhD���]�'�i��G�&��w��7)0� /�,����,R~���H�:���[{^�γ������I����n.Rn�+;2�'`_rSq�V��W-p'&S���̯գ/}�-��5_�hb>>�K�V}��o*������-�}u���w�є/��j���׋�d˫A��7	�ݤ���ٲ���6��+�s����Vl�Yt��%��Xƞ���[}�Lr�Hi�Gb�&�75�rNlcNH�c
_P���U��5~�
+e��c*�0q�8�:�NYн����� ����A-j�9iN�"�놁CL�Ck�(x�2vr�z)Zd��\��c��R�I�h��-�4���Q� 4(A��r�E"��5D�=[3)���u|ԁ,��L�S�]�� �>fI�kq w�����/�Cњ0u����L;.�����+N�=^~kw��T�hc�D���I�e��07z�����|aU�aHr���+��J�ߍ���p��m3_�k�
�rn�Z�A���65_I컐)Y��� ���d^#����jc�Ю�\�d+7��X� �TZY�:�"
P��G�Vx��5tYΜ��<E)���������P��T�ե"����3<���CD��k7�P5L���ʆ�d�j9)�BM~��!�������0=M�=�����k���ݭe^��H�"��ہ=�z�8e�rk��qUe�w��?��ͧ�"����;gn���	[0|���~A�p�v�t�otI�wtW�V�i��}�<�[c��E����1h�`��YS��.9��R4���y���ē��g���v���]/`�n	x-K2�5�:��kaB�ʽ��M�;-
A5�ܵgz̬& ���� �v�|Rp]�}G�L���H���>�5'e���ؔ����bE������Zg��px��?#���2,~=ZϪ"K�G��}!�ȯ�w�%�D�P{��zB�wK /��pIu~���c�����h��\�J?m�e��XG��hg;Yf�=BK9zm��>ٺ�_�!Q�f���KpWQg}��p��ܵW�vL���u����� A`��G�r��v/�&��%/�R�4��m�T%���y�A}I�E(����t�26��:T:��g�KϬm���ǷӖW�+CS��%�ؓ��,̜Z�)_���|�䃉�&�+�݃X|�f�1�Q�_�����o0'�����M�xR����F��Dl>F�39u^��g͚(���U ҄��J��4��M�z��0~Jߓ��ʳqw���V7�gM�7���{��X��hk�b.S��
�;<�@� 5�C݈CPK�gb@�:�� ���ú�<[�җ�����~;�E�j(-����+ed�lt�3�;�42I��\����x�"n-2 �K�.�:�(�=
H��y��.[vN{�&��`�	y���I��W����O� �N�3�-#Y-ow3:|�:���
^J4 n���"B�ϥ5��b������<a�P���p�{���;_h%;8~�I�����~f.�ZZ<bWDE��Av�0�!�8l5�����m� aͱ��N>5�K(|^:	������=�Ǎ��s˴jV����WfA�Ljf�75�[�F��k�h�tm��3�!�L ��AZ��.Q�/�o��m�L�)mT��'U1��r[!�K}��6Ս��;���s/c��� 	Y���'�*����o+W��U�Ma���{�^˷����
�; jN��A�6D�*�5�e!܁���mH"���>��"c�B5����ck���X���� ����T�B]�k^
bF
�7�:�������k�c�B-������,���(ܶ�Z;._+�7�co{Y�y�@��(N��4�M��/�,�7<O^���aH}7��2W)7Ρ�˂զ��Uh����Dd� ���:��ue�#IE��>���w�s�\��x��s �zB�'��E%�eeȺߚ]c�
@V�ک�{b3P�os�|1��]N�c�[����2ͯߣ�!�PfƔD|�b���Tx�W�L���Tׇ8��!u��@z�}~^$��_��T�
�CG��2O2�)�1
|~H�<Gp����:]U_T�1�J�0�������	˸v�+�����z�/^)��=MA�/T\�<�b��P����G��o�	������SQ����V�L�QZ9��d��WY[�6z*��;�s�T� �[�{��Sm��1t�ԷD��Ѳ��ʈ����� ���/uy��3�R��&�X��A:�Bj���Q�z~�=s��¡w�"^��D�"��<Sp����$d?똴��w��Vo�ķ�z�#y��b̸9P����;{�`J�l��=Ϲ�r���������7y��b�ۓ�:(�����^� 4�����r�b%_��R��@`½`(��Qܳn�~ۿQX?�bd4��`f͌�B��\YL
��`F4����VB@���i��z!?�e4 ���h�]v�_�|���yz�XEFJ�01�s,�M:�ۘ"#&[���"���5=�lna�����U��o�(uN�hz��S��#O��O��n����f=�st�P��o��*� �O}6�;a�f&<n�ֿ��<٬�FS������){��-����m��l���p闑Y�Y̓;b#�|غ��l��S�@;���C�3�j�I�fƢ����<�A�ku>�)g�A:�}}�þ�Ft�eE_j�����
��u�I��uL���g�p�e-�?3b��q��xQ�b�̓�e{D�r&�J���b+6�ή�X�jUl@��c~T�?wjN��v�8���r���&|#�-��@bT����H�!��\�pDt������.	�[����ݓ��@����X%YΚ�	djq�'M��0ۙ��'<�E	�P�i��A�2lsRm�vD{������:���n\�9�e�,�2�8)����_�֞s�{�N�.BZ�6��z�6d��N�"�)�+�Q��d7�/��#�djʄ�fם�[�Ξ-�L��:L�k㹳�'/e��%�؆)��&�%��i��8�#l!�=i	��6�-�,�Gv��/�ߕ�>���'�x��݂� 	�lkv-� �Wz2�����`h8����޳ ��ݿE�ôݨ��ȋla�w���>��ǐ��G:bA*ը<�TWQ�0]�w����c� ��j�Ie�{����#V
UP��=�+�3�0���ĸ�Z������XN���^G?i�^;��"�N���W ��c܋i���}���򦬿��,7|3�0sF�.���j�D�ԁ�_4�a��%wX,��W����/3�6�Ԓ8ă*hB}�(���P/b�b%_�>�

�������t��<��N�`e3�D�qH�6��Ƽ�i(���V��� .|�=Cߗ;S����ϒƣ��":�1�n?�]$��H����+ :�Wh����ޫ���4�E�l�����}ʓ8�pN�g�i�Q��5u�Zz��X����p�F�%�M��DK��2[��c$�r�nu��Z�7�QS�%�@"&�D�����W��Z9�Vx�`�σ~=v�*=�_��z���\��������ٺn�UЎ<�qr�1�b��S�N�t԰$.'�G���Ci����Q�!#:��{k�d)����FY���,NL3��̡����5t�f�BR*����XI��@Q���S;(u�k���el_��ݺ�$������f�~7��t�beb�Ri�m	���!�I�j�%[(�Ϛ/󼚻~iq%�t����j0��"Bk5c�	�<5M�-�8���օԨ�W�^0|��U޲��Mq�^�\�c�&�`����L���@��Z�R&C�P
&�d�0O�tܼ��E����o=�)�	��ik��En�!E�%��r�� �vl���3�Nws�"?<gm&���9���O���Z����?�K��mo��0~C��+�dJʐϡ�V�����Y��[9��h��]϶/z1ㆲ�P��|���fO-�b�U��r�6����?
d\#�hr�����3���+�w:���Gtg��@���Sx�\_�p����e4T�m�r��������7Z��3�qȻ��b��Đ���ne"1	�_�T� O��o���7Z��2�:[� l��3iw�:&2�t3���r�:P�>��f�wMg�3;��a%�B��}���&����M���C-�Įf�\�I�� �r���pyI.���۵��4���M����C�B:���T`'V�pM�-�Hd��5*�����E $$�����>��rt�E����m�y-�h������W�}�ݖ�!�T�������'����Dʙ���Ȋy���4�I�q Y�Q���d����m�4ZvU��=�ɇ#4�b]��O����|���=���� �o��v�L}Q�>n��g�w.����4�����}��������F�"�d�������7�+)VshkP��6�����Y�@N�02`JC�}NJn�=��T�cg�H�*mꧢ�!{��L�7��Ɏ����L�l[ƐG��20LU��]b���Y�ԁ���r9mLf%��@и�	��s�}U� ݘ����Buf��G��t�c�!�d2�<��?[5|�2/v��g�/��;*;-;�
�W�9��"�Fd-��h�n�Kd�u,w��i��B�cɇ��ihM�������xo���{�}���ohSe�D�3�vl�c��*�D�H�3DD�"�M�f�\XM���w��mG�+�B��p�}�ֈbe���G���_�L�麸��od&���U_���3[�nP��? �v�/� ��e�2��V�зm����&.E&m?[%�>ָ�ѷ�K������_?������ �< �.u�QS�r��&�9�}��$F�cf͡~�qƕ�u���v�7�uY���X���Ϗ��}I���+c���8�m�vv����#��[��u�s�����a)h��̗�W&֢�A��}��!����Ҷ�T�7������=�G��T�T�}��\t��(�#U�T�*�棫؉y���ߨn�%��Լf��)��eL����!����V���mq텅4�-��D�=����Yo*�Q ��M䂪p�+�[c��Ӊ�@��H7=Hp��8����>u��Ma|ipr�����FзtI� ��ۭ�J���$��;�y�%G<�8B�m����낀]����~��H�h1�c�q��$/�e�CT:+����B�O��hfY�)��-��~���\:ZuU5ׯ�Q��E�W����2L�$������7c��Ч���q�L���S6�J�$O9J��25ʇJДbC�<RJ2�j��J�Y�p�	��������*��QPnpMϒ��M~����~k��(_��#��CT%���ZS�#�M�{N]�<�3�"=/��lv�l��q%I��i]q	A�J�-3���>P�����Ce��kSD���g�����ux���%C)���BHTz���6a��qs�r�t�b�r
�}�,��:�� ���?��g���\�D�5g�D,��;�;�<��t��`�n.�fҖ̡n�r��Y���d��DU�fiI�"juv�����&Y����=m�o�#;��w�d�ќ	��u[�i��@�(�b��Csa��	����%]���bk�\
�K@�ѫ��|�?�2fk��Jy��\����Oi�N J��`�7�����!�q8J�uSG�u�0�Nߺ<��ro����i�`L���wC+��/w�;�=:j��G4d0�gWb�ȇ��	�u{�F.;��`� �н��8Z�PNcx0�7,����ZX:L��c��h_n�1��hH	��9�q���9�sə�kH�
��|��K�Uf�,-N
�So�6M ����Z����5�W�r_O5�"H��"(�kDTNF&j���<�@Z�.����*���q���x�9�T�"������h��/�d^�[��:{�f�� �:5�ňK�)l�����2�f�R4mt+�Ȳ
�B#N~������F�X�7͡7����!:��ز�.�~DKFޯ�zD��IU��#K�*7����O�U��/�W�U�--�O���W�e�
]�Ԯ������qͱ; ^X�}�� �Iu��n��S�J^Q�ǳ��N���\����#��ܻ��d�9!�6�N�-���M��N�~��"̡oA���"w#b_X��ZTQ�3�찝X��/�Y�4^Yq�S������b���O_�a���U.ʳ�P�=�ڬ�OW�������Z��f��}�e����*K�1�����H�����^VeR[N�jQ
΢�0�Yz��j���b����j#<�MF��xb��p�����lp�����C���e�V8��{~#�U�{(784*�Z��cb2�A�.{*�����9��M9z�׉7^`��b�~��A���ߕ-ǒ��3z���c��@�}��N��Yx��)�ԃ������BsxlEqίh@f#9,1�������>�`.u/���Q����l�UM�4���~��3����ĂQ�m����IS�z]l�aa�"�w�?���ҭzy���蜫�<�|0����:�裶ώ��������!����~��9]X}K��I�_�S7�n���KV���"ސv@�[P��w��Q`�{�Fc0V�C���Ȩ*3��v�ۡ��׆\S�v׏��nB���[a�_���.l����%ݬ��U�e��ْmR|�P���| �4�x��G�$�}Ԓ_6�-6G�Ts��++���lh����F�&��R �YV�L�Az�e�q��O��	�Ut�=³�yU��Od>��\��:�T9�W�4#��B�1i�� &�u��F�#��'�G?����w���}���Z��翽�*9S��c��Z��R��B�=�
Gr�n~��gCD�������U��mc�17��C�-����&�� R�R�\V	�6j����l�f��������~c��yo�����R�(xp,�r���;�f�^i��N�EM�|���\�u{���7�ŋ��-ơ.OT-/6(�h�hɊne4���g�H�� �к_-hcdDP
ın����<����%T
��.�9��?H��؟J3���W��������K�e���C��0�޺�ff+�	_g���e�\��uK��2��)'�ھ�(A�W�RAb�i���- ᪩���!<t��3֑oCX�"W,K�������G��R��o�N��RK��M��-���wO���F]P�1������>�ン�۩��&�w�bN-��L�/$d�݃��H�Mai~T����YƗ�R����T�:����c�C����\�Z��1�(3��ăE�}�,N��O��W;#��&�e�>[i��o5�6Ε������JϘԋ.�1i�% \~x����8ҊE;r�4�������o�VX�'�zj�ȃ�+����vr�ds���h�����{�ߔK��|p`[���w�K�M����ҢbH�j�D��d�|���6#��a�����F#|�r��Q"�0<f���s��+f�&��o9#�<a4Uq�u�LQ/�|�=��N�7���W��l،�Ov9p��I����D	�����tb#���yF���[w:T=fe}9�ܳ�x�+I��ϒ'��Z�^~�����9goM�6���B��h~)ǆ���3(\�S�TNq;d%S<�O�#�ek�"$0.�ؗ�h�4��}z�W��,����Y�����y���i��;[Pjj.��l%9����! 1�>�����J�R5\7�N�K	Nb�ӉSwx1��"ގm��%���\���U�K���'�Q bC��^#��N~�K�b����&sΠݷU��"pSd�l}t�˅��P��r�9	�*�E�a>$�ږ��O"�Y^��T_�!̋��E>�ϧ�hF����iK��!g��@�g����W������|j�V�4�q$-v%��	Y9.)88�*�Z��s<��7�Y��D�	Ж���ڱ��K���
��!�_�v�K^��Yz΋٨� �6A�:�0wu��հ�t{>�g:swK2=�TA薅ʒ�v佀o���ҙM�ǚ}��d.�@\q��0�Gٹ���p<&��K�RU����VR�5*�<G}���׌��'�	��Vİ�ۓu]O\�]��(<��k�=���� �� �A_���lb� h����k���N˃Ȝ�A��|�/Q݁^��0����.�Ø������ZbL?M�K.��8I��
%��^��U��I��Ѥ2�0�h�;�ˢq˝��P�[;�ěeۣ�;tWlK{)N?�9��`���B�:&}R;�ihZwF}��d����-zX��X��˹[���/��Yвh�QЎ5�Nm�z,�p0,����
6!?k*��<�#��=?�Q�������>� ���gɀI�+̾ ݜ��-!�*.�q�q���ޛ_�(_![�����N�/�Z�S95h�Vg�G(��ݑf#�L����v�G���`�>�_���6��bmGq<0�C��-���}��tL���s�֖�q������E�{�����T���\�i�L0�`<�&��?�	���w��uQ���]�~q�}��: Z�R�$���6W1�;:���%s����;�0�?��ғ��=���X�l��d)�ڇ������>ƛt8{<�hb)�HsB�H��c�]c�9Ud�Ը�\�L�T��b!��MiF���nyͨš�8"'��jr67����J�e�$G�X}7Jb� H�;��Z���͚�EN�,�F�0;Tl7�H6�C0���+șV=6Wv^"'�<H?�f�3�i@�7�r{yQ�������;B�_�V-l`:Gl�0��v#+�}�:S�*������]�U�{pJ�o7ߐp�С��]�����ʜt�j@�k���ļhN�O�5��i	<̭���[$�1�g[ȫ[�ࣀ�A��c���P\�M�[�:Xd����M���v�%������o���B�xGE8����4Hѐ.@v�����Ώ�]
m��u�1vFߘ�!$�&W�/*$'q�Q�R�|,3�|鲷xK��g�ޙ�nz���M�d��s��D6�.˸*.��DΛk?���*('D&�c�75��Ȯ�M�Y;* Z�E=�@���Z���&���{�e�[�����v���B�:KmxȐ/�H��%,_˗*t�7���W7�k��t瞮 �@�����4�ӻ� :���-p��Cn�
���q��_�<�?�}����K�$7�� �c�Y�ւ�R���_��������)1C�	�GjQ�H]5g���dyfh� ���{	X|?d9D��wK�J��YxK,
йT �)����9PƛQ��+j$���>��
���G���cf��V����P�*w�2�u�D�!�A̎�uYi&#"W�VsԐƧ�PE��a�����D�jCH��QE���}���It:���y�s��o2�RAF.T|���Ǜ��Z9q']+Xx���rad�zߐ4/�#kQ�O�]0�OT���\F�5��k{u��C������X'6�h��qr|x@���r�v�b�� ��<
}�C�/��Y�i��?Ðu�"��	I{ʾ���<�9����Y˓��R��y�`kiP�� +�W�ih(4�^e�6�h���$,s��ԫL@0�%i�	(���8�J����^7�L��r��ΞN�g$.�O{��2��U��k��Qy��2���]�:NL�g�L�#1=KwZωw�u�=�À�ّ�!� e�R�����k�ϯRI�#�����yg+���\���v���[����m�cƗ�^��s��t��a96$�Z�N�o����#1]�OT�_�%�׶�	�w�_�D3�n���f��!i(C����[ ���ԇ��ZV1"�5�
|n�k���H���6�V< ��p�|�����P�c6��R����x�����¿��J�x���~i#�b�*;[x��e�og�����x�'��f���q�W��C�q�������l��e�Zc�m>���*(Sh��'�L*B�]r+W�M�����E�A`��rg��.�w�ri��8V1j$H���cN�dJ3�C��i�}�'��Ïq����~<���m�*J���1�J�@�e�j���[	F�ג5�SR�7�����;4��\�d޶���]2�Kuo�NC���!���=�B!��9տ�k����(5��2�'��_�����xNߒ`L7�b�)]F�*�_��]}�����{��	VVr�������3.��='�����R��bN� ��a> ۍ�mu�J\w��k�']0J�Yھ�f��IB�cq~������?��������n���`��X�������l�sgX�9���t�I�0� ��?�ވ���(�*_�S��a}~8K0W
�-�o
F�6�N�v������? �ч���f�_�t�Q��^�;W��{ӏ�?�-�6�`eI����;�PmBA�0��k��j���<TaʹH5��ͤ�c�,L��t����ޜ���Sm����/�?�Д���S0�����i��6��Gt�Ջ���c3	Vni����
Y�{e�,���@�f)X�v:�k�%�}fvvb�8�����=_���b[aPM
��\�1���6��& ��n��8 �M��,Wg�9��ctj�ͪ�D�&�BJ%��y���>E��^�#w2(޾j����l u�l8[:�UhɊh��Ōb�R��T�^5��*��?�RR���ǃf�H���|��t��Tɦ���"j��3�L)���D9�v�)ݟ�摣4��â֡��@P<8� ��1�7Ȏ�b���}������~�~���T��_x.|��y&uދ��G�5�A��0e;+W�7���}n�Ԋ$hjL������.kp�ܼ
7�<@V�Zٍ�����̗�V�#I��z	�&�r�qY17<{�G��	�A����*E��"ou�˪.�D5�����5!��O�C��b����Rv����	������-�e�\ј�E���n�sO����i�r�A�p��kVcN���X5�;��|�MX��:�$�)$�<�uJ��"^�Ǐ��v�zx���BɈ���5��8N�[C0�1q���ȇ-IU��7��<�����89�UW��0�c��[����}����K]Y"ty�0Q�	���P�Q3t���n��{V�!H	*�SwG�xoH�.wkp1B��Z�y"{��$fSSr�Q�s�_�Q�B�(Ο=�����l֏����Ruw+3�M)�x�S�z�3�I����#��Be�Zb���(χ��Y�9�ū���n����"�{�&�o��B;��mX�N�>��l�nvj�5ߞ���x����C���sX���'u��+V�� ���N��&�J�hW�]��Ŭ`R��[♙&�C�`�n�[2Ȧ�D	��#oo<B8��>�'uíw�՛I�S��mA��a��{��F�tqf �e�����$�ruYD��$�3w;�@z�/(��ֿ����d�8�]��X�WL7�i^�����ͯ�ۤ��ɘ0G!���.�p~�\[<���Z}�%������	�����k�n}=3�5N��K���)lI�I��7��gx���Z��4�;�J�z&�pZ�̸�ع��Ml�S.Q�]#���P�P��0!wQ�{�bg��kq��"���7���>��,��x�m��F0��l����+�9g�;��N�c����7��� �7��{�[��y�]c^�6�'z�94�_���^0��(مK��J���BF^����G_��	�)���v\�
�jd� ��n�ú@��9�^@E{�ӹ3�Xj�e1�#��� �I��L�!��d�K��ۻ����*4/��xiq�'�YT�N��1�BQ������t���d8d�[b�(LA(7L�.t����LF�ĉ�l�EN�a��Pv@�(�j�$P;Lo���:C	0,�6����T���0�'�d`���;y�w�zI�CV����D��#.���U������*��L�!��>�%��kX(\� �9M�XS��ŝv���A.�x�_�fw܆ǩshq���������q�L�b�;`��/U� RrY��s�NΏ�
��R���b�i��mp�l��[g�3P2�%1�FjQ_�!�k/���[Q����F"�7�G�;����rr|IO��޽yO�˸��,C�dN���\g����[#&��V �s���ГV�<K\y�ez�8��|���"ª�.}�D����������m]�ⶒy��~([ �=�U#����2�Aj�����h��`#0I���~��}7>��Z�D�k��:�����V;�/|�q����߁.�u��P��Ҷl�Š^�ׄ�&A�#���X5��C�c��j��F�zKʛ�"0w��B�a}�Ϝt�SF�ӊk��G����8EeT7��Mg�+/$6�i����vǹ�\ëñͥG_A�ʗ])z�w8T�x�h���Xm�G�:�m�ִGK��_y"�Ά4Ћޢ��J�	g�a�;�H���9��(�!�,GhA|̿to }Y��+F��u����;�S]N0�gKe��x���7�t����#��!�c\*��'n�.t��zo`��	Fϝ��`c�FXhp��{0�E}��!�$9���j�G|�~G��6u$�#ho����T�����C��Kw�n�Iz�}�j��j\���{u^u����'���{穛�e@�!���_���cnO�q0�hj������/�ų�q6�-�� 9M�T��>���)�6��S�.������3�˵�%�-Ќ�E+C�O�c03?�^`��W'Σ�<��`�����oG�>aҾ}T���K�����Fq��rFl�5�gk2�9������w�P���B��Iǖy��PD�y�f��������C���o;\Y)҃��1�/�J�HEo��>%���!�0@&c6s�bHC>&��߼>�k�� 9Ǜ�d�b7�.�q�m%̼���������������Ҽ�=%�����X���V�.Q�����e�@�k(�N��o9�tD�B��9��>�Jv������r}D �r��:����,�����B�C�*��]�q������u�m�e��GQ5�dgh/ ���'���5�������hL��$u{����+����0J���m'��il�� VAT�lh�U�PQ��*��U�{=�4WЏ�l���1�*7�E�b������m$�6��������K�;�ޏ�͵ʮ�����[O�4�O�Z�T�cǼ��m��M�5>jtE��<�#"Ċ�Tj������t�&�S%v����c�W?��
:Z8!��n��]�c���C��`��-	��}�am��l�ֺ��N:��p���-����94�Դ�I���h�z8�%���X9����T�<2wx}2��ɩ��w�[R���EK�[rS��$T?|O�Vf���|.�!�- .�+͌8P�B�z���Uz�:�����Ƭu��� �&�����W��<����}��m2�&��'����P�Ve\Tk�^`��^,~q�VE��5����T�cy8a><��[��z4�r�S�UUu:t��5�p8O
�D�m,=J���Fv�
A#5Ș�,�m�D�:�6#�Ղь��gLuH?.%�*�9贤�ߩ�i�S2���'J�ɞE�k�AA1y��9���c�-���/['W����Y4V�B�͞W�n��;�=�NÐ��E
ｍ�O!+ѻ��͔�Ms�Pʺ�F[��I"<�� �:<��d����G&�7�2��5G4v�	z�oA}�Y(ɯ��n��ϝQ�0���
��W0�h�wHè��J"J��O�wH��;��m��+����M�	c����'p�c��L�GYީB������L�!��R㻻��T~2n�{���4'm�IkQW�t5K�Jl΍�9�o辝]͂��#�����T��n�|�]��+khZ Z�i��p�s:OpP�a댨�����2K�k1E��rhj����'>�!`j��1��42m�RO=���$S����~��:�ʦU�uv'�h����p��X|� +$XkX�l����6�Dq>x9��|����,yI��"��%1�F.h������� �A��B�q
���F�M���Ej��91}�z�$��@���{A6;�^ߒ�;]rL�/�����/�N�։}��QN�:��b�`�/��+�p5��Q7��T5`f�9(����E?��sww�6�,���_�^	���I�O.�[t�ƪ�-֙�ޜ�%�G�+�y<�5�	ޚ^���\kW�#��;^3u�U���B��%OiQ�TxU<4`|aa�zQ�}�\���[���Jb�����[��b^���I#�PN�dP ^�u`�u\q!?����6�F�6;R��D;J��S�WC	�y0��V���~q��?���M�C�o�j�n� ��ז�s�Qjƺ�§��k��d(2��2�>��Yfx��N�5௩J��$)}]/4(��`dH��5�P��M��M�����d��09�ŏ͟f��6��#���33hPO��5dh�A)�5k�䝴���x�/��f��9F,����0A��\'(�{f���x���9�D䟍�����Х�E�i� Cz���·��q%�)�k�m��M'b�V�Ь�m�mWq<)��Խ���@"��N�!������׽Z#�3�3]��~)�{b4<C�}%��z�q��ue-�ݳ@�eN8]�]5��z�@��ݮ��˗	H��5����Ef{D����$c�I,Θ=v�Tx����;�wU�a'�G�4�� l��&��n�%��@^sh<��P0��r}�R�p�T�@�� �V�p<]v)k�`s֞��~� ȼ\];~Ѭ�:I�Y�-v��Qb:��,tݮ+1�J�XL����;����So����kc^��+w�������m�,4V=��	�W�����Ү¶�k+,���K�"e\2Ly�%d�	H��V{c��P�q��=�K��[�;����.P���Тi[E	����`�\Y�{�|G��&��s�j�֣U
����sX�j�o���+������P��X�I�Q��>'��g�L�����YՃ��z4况́���Gp���n`0~���?p�.X��i�/KZQ[�bN���a��5c�ܵ��d�Lu�U�E��;y��57fw�����?��������5j-ʉV�;hSU[ ��94������P�{�z��&��27[��$�@;7 �s,էrVZ�^6\���Ϲe�YZ���g�u��9q��M�mC?�q���X��N�`�_牌u�+���V'm5p�KPZJs�`����"����Z���D���T%Ϝ2[˿�Qy'�CzZ�&��70��a���:��p��>�r���7��#�V��8��%�j��D\m���v�ZXؐ���)4mpd�G36�U�C��y�Z�,n�?tT(�v-,��4�ck�w��/z�?��>�@��dA�d���CnO�x�1����ר1S�W�&�g� q�����i'���������5�7���;�V�?�����'dp�[Z��`bc���YDs��Y��r�l�ߧ(��8�7O�	xm�,�@yŤ����0�[�>������3�6<�I�S��_T��71�f�%��n���i3�K�Ѯz쒧�/���_���2��Wr^'��jt���N�?)�dZ���^Pr���GgS���_��&�tB\cX�զ�
(�R)Uڷ0�pq�0%h�'�A�4V�a�:��U%�'���.�:�,G��T!XBR��K��!��]�̻@�2na��+c��{��.ފ{�<�&�9B�m�__Q*F� d�S\]Sb�,���x#4c���C���>P���j�AR0Z����0��:���.�<�U�����ڡΈd2�w���U�������|�C���ڸ~�6М�Cm+��H�#F�'���w��L0��5�!@����Q�VZ��*z�]���e�i��,Ճ�4��g�"�q�V<'@����U.<��+��3.;.
� �����lA�!�xIbs�xʚWH.���&(#��brX}��(�g��:�}ғ&���k�$�6e�	ISg���ـWs��r��[Cm�iBǽ$���g����0@��D�/���cb� ��H�����D"n�S3���4ݲ\z6�󹋍�4ETt�9�'P��'���}g�\v�;���W�Z���W�շ �}�h��,�N����%i{�H����L��y�*�e$�0x�j
�I,�S��K�(-��:�o�l/�LD,�Z.��Fဿ#l�'�wouy�Q僈�?�D���v����˝�W��i�K^��iG�P�Ħr��d��75�`�R�@�x���3��*�9u�)��U��)\>��t�ܓ���+ך�������b�Z��`hI1*���c�nh�UXc���s�F�^LCS��� ��FX�а�yx�ai��<C3� -�7�P�r*��5�G�F:>bŠ#\�ɗܛ�y�/|g_���q�:iǽ��j��z����RI�O�ڊy���f8 ��8y���Sm3{Im_4/g�ΐ\$��y�l��|o∣��2�w��&�,W��1T�}�^�~�����& ��VŲ}\�q��l����((M�ѳ��'[�0D����r��ʩ�Ϧ�,�QK�����Σ�ܨ�?�����AIE�Q�D���ص�.�U�U�LP�ٚ��P/@�r��2/8��fE2x�h��{���S�q�(u2�⁕��n�UZ�u���4n⏠�1�`������,#G����}��>��\����`=�+�s�vfF�rS��X ��{�)�s5*7d�˛}�����-�G�fW$���]؏���*#
�P]!Q�;{哄�v����>�Vˤ��� � ,;�1�6qd��	S�)��3�C��!P�,S��(��mO�6�M
�pҡ'��N�th�?�w�Y
��-- ya.�����=��&�T��
�/�J���;Qw_xn���� 1o$g�,���}�H����Q 0�ڿ�Pz�s-\�>�H)�m�$��y�1C򶳭ţ_��z B� fh)�0�o\�?�E��{��T��.@��le�Zd>�:�{8�.�A���Y�*x:�J���5���ʵ����l�q��生+TgV��*&af.w�D��Uf�:����X!���d��^m6��A�p:�la��I�P�~�}�|a�J;�S��0 �U��H�u��,�跈��5�v�L,?5P���!�r��$���J	?'���!S��k����B��ݾAf��P7V9��̪�SH�m��6�U�
F�0��@��K]>�ak��f���X�q̚��G`�bf3i��MJ�/!y=�ܒ�>�d�I���=�����y�z�R>�'��^����uj`}��|j�c剬F]!b�zT���O�O�����!ŷ�����$1���3��-�2ҩ�(VXS���&��bo��\w7� ��Z5ڠ�s8�9�S��"����/��)�	(�)�;�J���z��%�3�t�%��j����-jńqSA�b�l�a��h�7^$��J�ｐ��5zE�v��|���\�ރ�2U����Q��p����MK�V�P������ ]lk"<�uձ����KO>�JA����[��N۔x�c��-/f9��xH
�ʹ��5�9��f����G_�fp_@N�8.[]��3 �����c�� ��/$s��˷^J��\C�,Z��v+�1�ǲ\��h�����5���Sh�iSF���%,�+���1� osk�Y]�Vjq&��aE|^��~���x����p�/�[]+! �K��q���L<lg-��Q2�n�z�ǂ�fڿh�4g*���!�[������j�^K�RXv�/j���ibTX����qᬾ�YF��g���F�h��J��#6��7��!�ؔ,B,"�[�� ��iǹ�j����2H-��_��D��[�j�lP��䲄6�OQ���"�X�`��u  �PS��}���=���U����wxaBN���d2����.��Q8��{)8�� �l�����{e�`�J�ϥ5��Ɇ�y��C�$�n�/W|=�؄Xmu��鑦O *^ݰ� eV����[=��2��|���'U�P��E�����>��{=��!5B7�*�E)`k����G4l�������ܺ�D�J�W?n���B�k����>|��u�yERwf�Kj����G�]�@ߋ�lR��əF����}>�9���np�`|-���=�(!Н����	M��5��q]�-2�5��Ɨ��A+����p�۸^�F>��[2�U/5A���o������s����໥ֆ:Pz���"�0�3S?�YJA�:A{�k#�� ��+�$� ����c��7�6���bB����s�)�n�x]J�~��Gn2"�q�����P��,��o�(��J8��'���� �$iLο}�@g>��k�����*�v�u��<�;��wp��S���<�����U� /�~������g���Xb�nL=�x5�L��#!,��z�|f�����ua7("Q.�&�� ��ϧ��:�%e"� }ڊM<5���d�ZJ�g�u��rr�lQ7p��j&	��DRԛ��
��I���F�Xj�h�Yu%�J�f1S�E��u=��=�mk����f�:�[��邚`n0��&u��.ߌd �>]Bmj�x>�8�)�W����Sr��Qd\����N>��a�'`Η�LU�G��|�$�>�r��h����'7ؿ��c���Y��v� ����P������rcu�3���'e3oC����K2|&oB�1�� }cz����b1.��|0�_����3�� g�U�,E��z8�ġ��"�,��B�M̏�S,�Y��h��ӣ��4���f� ������{dPB��eZ������_��0�;�Oc�<�uWW�./m��S�(�p��)kɶa���uØ�T�ܔ�?3g��i%)�
*���y�2'�����!b�9X���p��blk�_
;�B�i[�c#�)hk`��˞�7!��G	�?Q%$OR}��=d S�_h��S�Ul>� �]�pˈp:r�uR,9�;}h�TPFSn�:�o�~�/ �hv�"$�-7,>+bG:�9%�n�t2���eV��>�q��ʴ�R�D�i������������u鷐hҴ�������=��pp��V�?6 ��c�4T�mL�!(b����cGgu��#&U�-��`r�b̓c\Q.z�_&HlW�&r��� 鴪'�|���G	�����t��n��Wa\n�6�]�s&�o0(;�g\U#�2h�!_*��c����d�Jgl�"7gFF���lCc�z��2�@F�Dog�l~����r����i^2�Z��Ԯ=���k!O�PQW�a
�3�S� ��V�*iX�c��!���R.}���P�~׬�u���E�S��*4��=׶���%l��~��i��w|]��`�aP����Rd	W2즷O�/���xE�R��]�Ԯ�Z���VF�`�hĘ$�"��W��ڜ��\��S�xQ����Pu�c�K	�Yʧ[@fp_M[%J�!E�ULn/��SZ2�����&h��y���p����U��ŝ��A�j�3�bP�dvm@Ee/��嘩�t�Y�Ym����%@��ƠsFG�뤥�`��9��e�&y)]��9�2�O�����~�BT(��^jhY��g��쌓`����9�+D~�'��'nOR��Y׶�1^\��ZU-SlB���	�ۯM=��Y{.�}1� ,�����=1e���*����Q���i�&\�U�>@9�|@����m|��9I�-����&k��
�m�D�����6�o��'�|,|=!��2�2p��կ�c߽)x��c�\��7��i��AO �:=�Ӈ�y8Ei�%;Ϙ�O��Vi��d��+� �=���Tǰ��4ϫ�2|�_M�Y8���m�x�������-ö�0wI����=B��fF�9��z�z'T$�! �g�lb�h��v�5�C�|�$�w-�A��#�*�����=Z�;n@Ⱥ
%��#��U��P��T�d>�{F���|":�Wـp�����uR%WW�ܷ�*]��N1����Hv�`й�ɩ3S�3/�A,؝��|�2�����7��/�ݎ�G�&���_D��HGI.�e���:�%v��R�
�K��C�'\l�CC�����	�ӑ��`�a	��º!]�����M�T�J��P(Y>������I��%1N���J��n.g�Kj)2OF�$���}:R�xV��b�ʤ>O�����%�Q�<��8����j�r�?V��$�c�t��lM��OdS��{~7�E�Rσ��*�x��n_i��i�Iٶ�O6�j�`2"x��ǥ1�"�I��b�]�� �
(�	h�z�h쑵��ꦞ���ƜR�or}]38�7u��/eמK0!�d�sE�>�(^GaL��h3�.mj�JM��߈���]�ٌz0G�~�~��ucrǒ�O2���x���7O`�H�sC��0���7=r�s��bI������L�6h0���Xc��=x��U@���J�g2�g5/1��R�].��\���5/��j�[�u_��0|t�^8}��ά��4�� ��`�Z�,R}_��9��?�o%\W�`vmh'w����6y��K��r�AD�SS���H'4�p����x��6G�u�:���'z�q�C�M������u�IH�Ś%΋�s��eQu����p^B��1������T{�e��=�<ܐ��|9�7���)%�@��6�!�ri�B�!GRw��N����d���o����px�^�||3)�R���+E��(Hè����Ż�zlV�-xj�� �	% ��3�[�T
u[�SC���Q�oy�/1�H-<��*oq8��n���Ą \x�+1]5b��6��50���2�;d��v�&�E��ܕ��������|Vvd���Y��F���4.0E��.L#�`.r��RL�0���Q����W�g�^�y4��	�M�3�ܻ�H/��|��{��ӈ��j�\ugE�#�"�7��!�X��1�-�p�m�%��s���=;^a �t���Nь�n�>�B7�_Iu&@R�Jm��u욮2k�jG���F���|{-jkd��lz�s�NS\i�s�3��6t"���v����m���Vآ�l`�#���g�<�)�b�^�;��Đ����n����z�׉�q2�=��Iv��,S3>`�F�T��oL��`b�䣫�J��B��ǀO'��|�Y�M���dȀ��b_����+1U�^��Pء�*�lXu�}��u�y~��D�����X��[�EYstcDP���w�ߜ���!��_
�АI��84��:���TVup�jX�{ p�UM����6�E���������j����/z=F�\����Z���+%�.C�2�s�-9{Y��a�ȿ^9d��r�j�3���i�,�,<��,1�2��^����L�{���?�5A��5��6���m��Y؛@�~{��j3��Ak���1%�B�Ө�Z��u�fO��#�/��?�O/g��mI��̩���x���QJ���#������*�5�I�q�rz-ⅸr��Xcg#$,�R��G�L�oX�W�ᓣ^=���	�Qf[��]�ywf�_��!S�2u���MkI�^�d5��l^�Ռ��#�0��#�_�ML�[���H��9K���ڏ���DWI��D������SEH�2��*T�}��}0K�k�96 }��~��+�N��" ���r���H�=��4��J	�;4)"�hP�A���t��z�|�.R�C��zS�y��UWL��c:�Ɖ��Ě(r�R;Y�� ���ұ�����
��i�w�Ma������>B��"zG�@��}6��V�����{�o3@�c3�5#���~N�8�%o�!C�D�Q� D��l�Ws�Bʵ���!��5@�g	�� ��Y�vTa*H�iŘ^���Ͳ���x��l���M,��J�e�5�7/��I:A�mջ�jL	9�A�'��4��%� �h��S��{��sJ�������9N(j�D�5Sd��xC��6���9.��s�_p��R�EOx'E�v�1Yylb�������pC�͜حP_=�,����Sz�%�����CFx�jP��\�`���|k7���y��M{\���|tD˄_`�+�iǗ�y�W�Џ�O��3yk�tUgc&x	ԣy���;J����'.�Z6Y�����s���S����J�k{�+J�\�}	?�Z�����N|֤ɗ�;�V�KԘ����8�P��
y��h�f�;�ĕ���,A�M�VW3<e���rUDŚU���`Rg+��Yu�AGK�J�>7�!kqԁ�� �cHi� ���6�{ň3
l�l��m��X�t����b�˂1����ݖw%������nfPא�Q�
��֐��Ø��
�Cn
3�Ѽ�u��o�iN�.(���C}�o���׎:���� p��a2^���/��`?2�����uÜ���܁�&(ٰb�Ժ�Ӗxk6`�O���9?�x�8�c� ߿�`L�q�ɍ��_�1r���A�?�1���j������b��d���24�����7�Ih��&�A�'��	n���ݬ"ӽ�r���=��m���n
�ڨ����ZL�K��+,�"�3lYm ���$�j�s	M��lH�rf��%|�8�'F�4��(�Y.wJ{M�J�rՖ���/���J��=�O^�C-	�9��$ů�KgR���ij�a���Ȳͧ��!�D镽�������ci���ɯ���<�Eq�/S6F.�j�&;��) �n�s�xF֘�%�ok2ǩ֭�jG'|�cLE����l�����}O|m�7Á����^�L宮�s��p\F��Y.?N���� ך8Vi�wУk���@�2��n��#��g�7��m]��]�Jp��¨�~�w���B5�fz5�6�}� e� �#*h�j�G� �r����f�0����T3�)T��)\3wM�0}�|Q#p?.]0�Dj����x��"�ɔỪ�CS>���dҲ�ԣ/D@�b����$�O���3,�0r����	�$�����@sx OrG5^��A�c���F^�/B���W'���x�E��<�Tk��هe�%�-�.p1"��l󣽣�Յ�0��/}!ku��"����?^H!�}�fG-�&'�*'��T>D�x2�<6���-Dd*�<�CV��)�?<OzR �:g����U��"m�Gs�.R{-���;lP]�+�^)�w��y��ގ� *o`і�5��a��wXzwt���N�o�Fb�lŤ�I����^�(
�aKs�)�t<�N/��ATB$=����G��@B<D�m�����l�j캪���f~�M�*��7�0�/MY�n-Sd<�G L5?0c�/;ld`��̼��#�'���������b��C2�ߒ""?b��9����mY�G��0+d���:�1�3��~[<׶�1��ÂqUP�$Pq	�w
x���mE�#��l�e"���OOa��N�q�{��+���3	���[i�7@���6��\|,�
��}���"��d�S����G�T���Z�����r�H�l�0ȢA�Y���-;#1O�����c���(kI�;c����
��|�`���%��A%Qk���z�ʯ���}Bu��/"$=�a�@8���n��C��T�j'D�������w�N�3	�Nn��
'�4�U�7U������x�IO����D$]�]R(N�	�m� �INQj����kJ�V>h��̄ &���P�{.�3#���4����o^�d����r7L]�[�F�ز�0+cq��w�V,��@�Q�ͽ��2��Ջ�y�k@��;Z���c��,E��@��6o;ٓ��4c�����s��?L��Ҟ�b����]��zm$��"ou�ȑ�xj	1��1;8@����)+^�;�/�S����g�8:|`[����p��E��P{�����=ND(^pł8䳒�P����e%�&��.�4I������O:��88�B��Q�:�����4��AF���Ě�!T��_�sb�8N�^��Y)��A�nj�B� ��K�š�%ߠ�5���g��<�i�)��;^<�����p����>��1���"�U4CqU��h���ī��`P��Ђm�� �g�b[ԭ�a6��s�6Kt�r�T�D��x�[V���dB*���=������9 G�w"E1<���(��N6ߓ��]x��d�Hd���LͤR&��f�^N�x�=�@��ŝ~��SDj��X�V��ʍBrt���k����U��f�d�����ˢӁ�>T�!E�����פ��u��	�G!���W�Mh�;.)�~qd_ �z�����j������f\�e���?�~;��#	��kZ0o�5�ϡ�?E�Hin�O�8�=h���T�F#��ץ��N��췽�E��6���}�~�ز���3]@~2���IM��Vȇ]��_Ayaؚ��	�q)H��Bemt��������W������b����5<�}���4�@��jvե��Đ�{B�Y��=\i�`va�7�K��I�%1nZ���Ւ��.D����b�:�ƨ��8��*)2)�$�Kis#�W(f���X���}�\�U~jJDf�,�r^W��8[�÷W
����H H�F�\�e�i���*�N4����~�ML:���@�_���ĵ8\]�L��:h���Vo�ų&�iMN�V�`����5�䤂���5�yH\:[����1��h���)�pm����	gdR�Pf������{��7R�W D�tM��0�j�.�d��Nd^5a�QAb����kIK_;-~c5�y��M�#���J�"�3�ł�`L��K�'H�`Z���X)L|Zqo����u�v�����hl���hI]��Q��xK^�Ò�`��\�`ȡ��L^���^��1]�n\�W��<���� �h'��fMz��'��X��"�s�xP� l�`�|�/zN���N`C�b%+�&�J8�S$KUʈ@�y.�s�$+�aCK������Æ���ٝ,�I��
��k�"s4PL	���C���BDt�7{5��hP�Ǯ�}3���"�61�m!�A�[�g�e�t���$К���*8�~�P�AЙ�'G�R�4{�E�C��[ز�=�.���3�,u^,�C��>�+�R{���E��(�},��I��6,����E��z�K�S�樾�S�"@^�2;J9�3	��訜�L�$���9���Oc��*�,KP%r�����|�:B�{P�e��h���ה�� Lo��p��~{�Y��׬�"�hk��0���*�{W-��e��D�'��	�.VR�9�cBO!%2�u�J�`=Uz�s�vl�3"@�b�<;ɴkְ)���0���t�!ba�%~Kh����CE��q���yQ���W�n��������7��x�jd��^
ts�CP��Ok�6�]�Xfo��7LJ��������
�B��u7�u߶�Py<"LJ�6 S�NM@E��o��B���=��w�B���L�em���V��r��wf��;(>��^ W��v өfm.\�� ��3:�ׅ�����a�F�hs��������Y�&[k�#?xsyB�ԚJ��8FfX��1]FD�=���!h����!�Z�=�"�\��=�]H^�VX�HZiG����.c��(�MhH90O�bX@#�k�&;Ipl_?�哧� h�[�Qkнx����x��+�7n*���07����y�]��y��DxXvg�/:Uz�*΀2�.
mF�4�h�����A��깚yҀTW�-�*� ���C�Y�U�>���7nX���$+
����g��cpN��Z�;=�)��`hJ�84�Ӭ(L1���G��-=�9��^��r1Qw7 q�'XǾi�G��WL�t��n׿ ƠA N����{"����n�~���X��!眦qu�>"�KI�C�3$5�:f{?m�@;�J���
J��z�"w	�.rv4(�| �t����u�*u�0�=��5�TBѣ?�%�D�p� ���j�}���M��C�G����R8q�$�_a�яr��	�)�?6Z�����s��t��l��sѭRKg�U�=3)4`9��֫7~�S+%`]���z*�<��͡�p� ������0�T��ðJ�5<�o�������$@ch�	�+K"۫��
��Z�OPs~/c�<B� K�/��QJL�'��z�l'�wZ;06]�
j�M)�Z�"7�Q�rO�}m3�ܷo!�Ǥ]�"����/�e�`K��v��{� �1T�����#G��z��#��,A�9İg���K��5�A�H��3�Ȥ��0&� ���Uf<�2�KF���$1f�������(�����΄�O�Ӱ�f1��_�~�e�[!�K0���t&�/:;!�i�D' �$:��ڀC�ޣ��\?�J�|%�X�*U@���P�,�rN�E;\��2�dEl'M� ��n�H�}{g9m�X��&e��͓��
�QS�[q�9-1�� �I'=��FY� 6�	����+'�2�K3����x(��g}�L�'}�T����* �y�������25�o.��;�&�fk�7f}ϩ?�"��.�=5���l���A��l;g���σ1B�=�"+Ѭ�-��P_Q�nC�8��{�����b�k�\`dyk�{ԡ�Tzb��������Ou�� 4�z�o��I��W^���.��٪/x���M�~�b�Z.rY��i�/���t�(Q��z����+a���z��1�ݷȎ�"ԭ��?$T�tk�*���rM��
���$��'�>��c|{�����̉]������2�������!f�CX��Jk�P�Ǡ勷@yF�F��a1��D�<
�^}��
R=U0I�4a�y�UM��ZD�M.�J�BqQH�'^�)�>�B�	7+#�Ļo�ۜ��>�S���v�U��9����7�,�$��N��}�
�6��^��bq&� aL�8S=};��` w^Z{b�S���9�To�|Ӝ��Z�+�}3�w���z�,t!@�	��~���[V��
������&�ru����0���c��N�զ0�BA��j7��C9��w�Q֯�YQ�Ò��.����H�בݳَ��nl����������Ha��5(b������Ʃ�Ŕ��6Q��gmf���A��w͌S�߯�#^'���������k���XZ����yT�V�B^��ܗ��p�E��ϕc:dl�0���G+cc�Ő��!���z:P<�F�pgX.��`a�˅S��|�ͽ�CdzVN|5P�(I�<���a�H_�b�c��v������^��Eqv��u[�*5I�m�6 ��dsӏ ��q0��O҅�X��9�l8b1�N��p��p���J�D��P����C\"b�2�K"K4�Sl�;x�-~ؗi����%n�����6W�̧T=��]��Oxꏍ�X��k";��a'9���� )�"�E�q��z��k'+���2��:4"����JRZ��������=i�_k����Ά ��������9�����t�@��������*�t�'�}}�Zz����w�3#�yP��S��_�J2��Y�5��56��X�o ��Y������/Ii�+�h�r�'�+�p�2>�������愈���n�������S/�j�]c
�Ќ~�X�K��C�~ݖ�>o&f�&��&�!$W4�O!(�iq
<g��|kD�XN]$8�͗���6Ƥz3���&���� �ȸuP	���82:���M<r��Is9_v���x�9FrB�h�נds3׋�U3%̊nG�m����4N�}�����9A��Ò��]�Sc��kј�U�����+��*��bn���MwS.4X��3�_�"�"\̎��}d�#4��rr��ͻ�V���5
B�&��h�R,3C)#L�gl�>��T'��c���|�ࡀ�\�${~ҜY΃�h[���
��آ�xkU�-+��I��C�bH���`��s;gr<��	=1��o"����[Edh��A�s�X�p�doPi�����*f�b���#�K4�ty�g�&Z�U��]�k��'iBtƎ$�ANݠ��pOM��<�"L:s^��ă��_k$�#�g4��
t���#u��0?�^0���~������,�)@�k|t��<������Q
��7�w:8 �s��8̸F�='�=s��r,�C��_^��?PO��j�C�v#J���i�	@-Q��k=v�q*�1�yS��w�B�@!	i���T�xվb�ͪ�H�<Ѹj�9�(�~}1.��&�z˖DQ��Fbz�غ�����i�%���T��%��C��mK�q�>7��X`�_��_r���&����m7��O��gn�Ի�Peq��+�XF�D�R�Q���mۜ
�@�ѳ�	�P��gg�bq�K&�us�;�؎#��a�V|�c�v�J����溆��w��9�b[`z8���1��@֏)���{�#OH�T{1gUtDء��t�N󇴫U�'���y戺81�����j��J=:��R�R�a��>]�:2*�w�:᪂0���!��IR�:-Ы�A����de��eX'w	w��w`�D�e$�r+�r�=���4"+�q�')EU��(���c��Y:X�}w����� �B���뫵5�=m ���~�Ziz��4?�-K`�K��|��_�F��F���������/�T#��m�b篲�&��秩|�����\ �id���+loh1(�����R<P����7��(�_��O��]+f�d`M�8E*5��=�".�?�@Y�[����?�1��x�\̺=Ϲ���?��r�ގl�9q��v�4��=Է�gR^gq�`"}|�x��-��3Jb@��[�s)j��*�F�"�C9��Z��������I����݊9F�E(� kv ��ɕ���XB0��l�F�O->�E��q���Ҥ]`�G��w�44>�y���W�:�0Z:w��K怜1�ڨ�MG6ғ+�Xpv��g:M�;(���UV���eb��<�hV��n�����ݗDظ�=sJF��L} �	0pxWT�@bn�쿸�^|k�m��L��#ŋO��X/��X�Հz�WfD[�JT�:f�n`P�������y�2�Ж0m2k�n���eP�{*��%Ϫ@�*�0I�X��s� �}�9}�+A�b��!�@L��Q@O����L�%�"4�����iZ^�p<n�>��	1�t�{�{ƈm��3�.F,B�E�Cwژ3,O��U"����+�L��Eի2�ka闉�z߶ZrG�ѯ2�<jw	NW��:��+v��܋�����zc��ޘ�lWy�$�3qk��l(>��c��.�Szz�ԧ+H̖��ڟC5�!ƥ��Xb����-�:�g����[i�ܘ6eɸ<�dP #`b��<ͮ=,禕^�IP�$�ҍӠ��ܩ"?�EC�D'�o�a[o$.�9�d,XE�gn��d5ˋc� �V0|���aƩ��E0N�\|��!�f'R�����2�D��@O��c�@ΝCW�q��d�I�$5%U<���d��Ŏ�pR��,�z��O����hc���kjՀY�#\Cڴ:�|Uu� ��c���J=_�v�RR��ZFi�3B�s[��tԞ�9S��q>���]j)[�(.T���F���v����1�$tZ�/��d��k�
$I�da�C�N��dg	+! �����{b��|I�"2���|mj�ȯu�!����Z�E�K���U���JC�B�D��m~h�w����S��Z䤤�h���>n%��K�a��]�Xv6 WB���g��P F~�S݋���k
M�V-F�����T5�8��]�kj�h����(}���4`����m-H��[�
Cp�W�ˈ?�h}�Pns������;�p㣂<��	3�}$q�NQ_s]e�GOR;�1:�6N`�B��K&y����v/A&��
H�T~�C5��,��!Π���8\Q+ڃ���}2W�Uj�Oυ�7���۱J�!�;�4�[�F��]�V�c�Z�֗Y��2�ez���#�{"��w<���b��h�������EP���e���>N�����-
\B.�Ԥ��9��ѴO����T������
%̧�͛'�����	��;��~�Ug�(;�w6���^;m�o ��^��,���i���958]W�P����o���7>�Hj��uʭ]7���j��p�r��>�1s�,�~��qD�W�����I{ȉ���覾m\�yRz��V;@ d�� Bzq�[YVګҔ6]�5��7���9���n
V|E���ܡ��꾜{�W�V5BK���d��a������6�Y��ei�au�����a�.���A��Ɛ�� `��w>Io/�i�Շ}L����G��:�6b��@����4��|���G��rFq�rfE�C6����+j�ֲ�/�6����<8�w����bc������n���?+d�`�����V�Վ{��)^���7���,T��;��z6ˇa��ܹ_m�x/�5�[w���3�39j�[ͯ��K^�T�"�%��u7��r�Zt�R.��X�a�l[n��΃>�����E�۝���W|4������]\n��_�\d��B�#mBƮf
��'Ɂ#���Ĥ@?�j��t҂��i�W���3D�e?{~=��m��]�G#N�p+3��B�Dw�=��"��)���6�ሙ��]=3D7�ӕ�s��0�'I��I����Ղ���k�nʓ��"ߓ�|��Q_|2W�ozC��x��bDEq=�籵lo0�3�#@�$X��w�F.��w����`	d"I� ә�X(�&��v�������c���� �[Of���ݽ� ��\�˧g �ghb���̯�Y%�'7��й��1����U鎀E�W�-��Tυ�}E�䡥���G�h�C`���$pQ��i��t2M�}z����ܿ�S OM�ɭu@�*�P�[7���F��c�]¹uF���Bm2���9!�!�ʌ'���:"��H��_�R\p/2�K>�����\�w�=��7�]�n 6���ƎW,dH�F���/
ϪLE�e��]�����9oi�9�?�����ۢ�Σ@�[��N\�o�9*�-�G���.�b� �{�.�����)�g�	%�h{����s���[��(Z�f
�OX����f��H�.F�UKi��|�&�i7��,V-	6 *�j�q��r���B����2C�0�.���j��7�K�*��RZ�Ub[G�,�`{Xx?Bl�	*��פ�� �����7��S����Gpͪ�#?k�/���H����#�4F������|(.�^�TN�|�닣W��flI��7�� �8<f5z������ʵ;�rw���t��,ڏ�5�_8�|��J��J'�Jd�R$�qHY^�=(`� ��H?�A/�Z��E���~�\�3��w'�^��^�!4JT�0c]$G`�!գI��A�����+�)e�]^Pf?�%��kތ��]�7�d��G��г��VǆO�7�t��U2�����!�gs�wEnԿ�1���������X��]QƜA�5�^8��e��b�I���=��h��`�!]�)�T�	$�4Z������x�Iw��O~��[L�eS��P� �0f�ۯ����3��dn,V��T�w�˄�i4�=�s�U��GzS[��kԃB@AZ_������ՉҙE|r"A�!@���K2�)>����>O���k"ԙ{�9��X\��Z�Q֊3?;��s���W���$oJ�\	SV.���:h�K�a��˜�VA-� �L��!&�7�_朙�:C��9���jI��vK�*��]赏�!�Dy��9�T��j�\x8�$~;~�7|k{��������F�����z�$���2�YY���` ��+5��ư�"BJ/��s
�\ș���_��pmot�&�S4�l�,�u���\���\��9�u�ow�A����)nb,4��'��t�Je�6|�c\�#[tS���#�O��t��42�HB�>=� �F���sW�m
��ύL ��I���5`6d�C��NQ�<h�~���������<w�x��ah�^��M��[�?��?n��Ә
\/��P�p���m�صX�l���Ja�I4��L�0ݥ=-�%3�+ZI�fjp��a�����������W9�y�@�lm+�W�4�u�}��!h��j$�4ڶR�����q�K��q�?����; �o%�jŞJ���~�-ן?Q_���M���W��jD#��"���9>�f՜ �l��`d���ue�W�G�������bs��4��ț&���	IgW�/�wH6N�!l����2��:n	k��u��<-� 3�
�ݩP3m�s�w-�%���.L�@����WLaJAg��x����@��9����)����'H/�h\�f��1J��;[),�z�ܜ����$�w��.h�ϐ�u�P�O7u��25M�^b�nu����l��I�����,��,APοPV#�@[���Y-��	���#��3c���V��$7D�+}���M�-e�q^i�n�_D鿰ό��-v>��xZ���6t�)|������hOٓM	�~2���k�t�ٮ�
��T�,���*h�Q�ǦR$��#XVȋ�x2�m<T&��US[bd$�Hs��T���y�Y������+A�i��?�F��e�Z�_���)�О��g�z�F��Tp��MR5��5��Ȋ�k������"�n�2�T2+		D�q�{��U։U���B����Q�f�����&�m�!�'�Eb7�n:{=���]),���[�*�|%���-�ȫ&yH����R��ۤ�R$�:��Z_[��=%�]�������ó��R�����*T�Lɍ+�^��I�`��yͯ:v]]��|��i�Ӛ�L��A,��>��gܵ�ܹ7v�%�t�D��,̧aaY��g�j�)l�	��"g��Z�|�&�Н�N�ÜgB@�[:Ɣ�܊���܍�gm6����ׯ>�S�w���kOɶ�	�d����3L�A�K=�	>�������ʘ���)_Ku��H�0?��&P�깊F�υ@\����WnNDV��#P��~� �,�>��� wZ��`�૯c��Ra��-��/�&�b�'����2��ūO�-�OCu�:����"f�������p6��T�H��뢅�%{봴-R������ ��ۋ���
;XCpsܖR̡����.�����ewp*p�� �j~m!����Vp5#��p1t$6��W���<���g�Y��f�8�U��ľ*7s[�P?̧U��W�������݆	�i����&5�\h�f��	)��☱���&��%6^`[m�=�!��^���ք��:����ZbV�'�w��+���z]�گ�DB�ܙ���[)'[���Xɓ�vY�H|rr��I�������­�� �7Y휹q����5Fe�Rـ�Tx�0��mG���W� �������#���� �E�Q,��PO3x��������ݜ�?��x�3�[����C�gK��lo���"U0H��YC�c�f_r!U�1�O�xw�p+�,wJ�XXڌ�(�ihBd���G�,�qE��� ^�՝�M����7iݏw$Nxc���
��˲D0���ӄ�׳.gHA���ݲn>M���|1;eWў���љ�8/5�}򧶞���
���iW�� ��$���.y3�|�o ©�|�YcYĥ��io\�ۄ:]���<��^�I�ٹ�A��5�7Qk�q�.
ϼK��4�b���݇�'������"f��(��u�.rq���/���b�4ݏ����c!yK,�M��Kԇ�С�Sk+�c�aV��&�C���&*�}v��_�Q�S�:e$�q���}a�Zjx�ޢ-ԝё�8#�$n_���p�o,�~=�i��T�S@��:���?�8��ե�[g�	��9����9G`��h]:/��B�Wqx�P�%%꟫4�<��R��ܪ�-�`�,_7S��j��~V��t�p�6F���_0GN@��L��ꉀ��2��_lk5�B��mJ�]O��.�]bh<H2:m\����T���}A�[�uΒ'=�W��L2�������!b�U����-:�|we�?J&��up���
�ɞ����	\��1x�[��+��-��D��v~#N���7���&������L7\]_N��"�����2�gw��5G�h �*��F~�d�:�	�{��ԐNyҼ	�`�<�Y�Sն:�qQ��V\�%��vg탙���$�(�ęY!��B|)���PZޕ�Z���	���CIR�!�`�eR=\��	�cYDM�MA<㺹�\+�G�<<���: �v�p%I��g�^;6
����"��K���~<)�P���d6��N�*��\Q�- ���G$b��M�YK��&<�4�.^ϴ$픩�[D<K�Wk��Wq=�� �̴6I��q b=�2��PA�EbZ�'�3c肇{-�c
OTZ�D��v�M<s�A�jIX�ý%=\'3�i/
!���R搷h��4 �.�>U���ls�ض��/�#���z�`�<1��=a������[Scc�[&�z�I>��B��j�^�y�N��D��,�|<B�T�7�ӦU|�Y,���bi�s�Gn݃���vֲK
AU�Ld�Ҷ�U�t^�0���n�ׇ>p����1�H~�r¯7��.�o	I�И� ���F�;������|�u�j�����Е���,�ހCBg�7ʥʵ�l�g=��0�m��ۄ��_y�"O9�W�C���{|(��	mq��
����~��q������(b�(��� ���?� �Y6�q6ǐi�x/_��Ik�u��|��<�����v��
G��7�3>�ҭ�ѻ�q�<�x�4{�-E��a�EZ�:j���Ҳڥ��Q�>G\���e$5�>k�I����=�֛S�i�i�t9~/h��
X8  K�Ϭ������8�iRR3_=��!�$/�P����b���"�b���lW��^?�l7n.�=�>���m�K�+�rn�RM_n�tӸ,c縵vq�
���P��o�;�QP7�:��X8�Q;�&�~_�"�L�F�͗�h3UT��,ч�L�3@UW%7g���U�1�m{ �&�1��s;�Z�/}/���k�e_�5^=38f��V��?���q͗�0 ~g��ú�:��`��H4�q��9�T
�Ґ/���P��%R���M�@�m�nm��lQp㏽���@����S��2�ͳ5.�@�Т���J���+� �>j<�uw�3ʕuX=6�G��=�t<�`��}qu�L����%"�;UvV^S��a�������4���2f���q�4�X��ps{�<�V,(ub��
ǆ��q�t>���`�`���+�|����*k?C������U�/(��d�I��[nMf`p�-B��N�U+��:�۶�T��il4�]m�Y!�<�l0oj�M�|Q2���mh߮%0�_����r��[ĳ�t^t"�v
�͝�����]�	���ln˼�	sE�ǿ��姴�u���qnT_�t���W�sL;����N��2rp�6��!{A���ܮB
�����^+EGJ�t��D#ٶ<�ٛ��=l���m(}Phzx
�$X�"���Fj�b��1��T	!���>��Ɯ��ݭ�L!�Uq�b�zr;v�(d�1E�^,gM�ZA�x��l��HՅ7>��7�p�L���%����|w@�A��	ځ"8�m�!.o��\V6%��m��|�7qi}>q�j�(��o5�+:u���D��fN�"��M�]��V3�#Q_���X1����������7럅�ӆ���20���;�0SP�h	e��1��
�_�?�/G��^(mr���Y�xh�Z�j�6ż�)!y������ބk��d*0��BS�)�VA�U?>	��L
�֋uM~��Ÿ���*�+0�	]�x��E�鶦�SoR�_�a	�FI�W}T*�~8��� �"�5��@�&6�XPj}���eD�������4Ӕ���h.3�!�ž��"v��2~�vc��-�Y����I
t�h2}����!�/�P���-gbߐn�ͳ�u�w��rD���}�s���9���x6^)M���!M���"���qA��XԺx��E�_Ґ�!ɏM�2ƕ�ڶ�?j��eҪ�A`'3 �r�\���.�wr'8vX�Y³ج��US�li����/V5�S�TD9��U[�Xh-�磤&��#�B=�ܢ6�W���$�|=��"�Q;�^�{�)����vO	�~�C(u(�B�28�����JD���׹b�N>�> .��Z���t@ ��z-��nл�pX���Mo���fK3�F�COO�������%��7�v��|���R�s^SڶX�4Rw&�@_��*�vq�B9<�#���t?E�W@jx��T�^�8E�c�!����:z/p�Ϧ!�L16_�UTE~�Yɩ-���:L�-K��<�쨡�o�t�]걾{q�T�?�>�������@��˥x$��u9�q�� }~ꋛ��+{�lB�����Z �_|Nb�]�aE�9�.:[f�\���1�8s���c���K@R���i�~�f)�-��@�LT�H�G�������@y��wߠm�Ca���;C���S�,��8�D������Lex����`���བྷ%Gl���P����A�������.�WS�A>s��lY���@���˩w �(��MK�l��D����2��U���<*@���+�����CVh�l0<*e��i�`��_��4�$�4 xc�� V�5K��*@�C�*�}�Z.�e��ɠ��L��i}�Z��U?հΉ��%����g#3Y���#�NK|�����绶6��ri%�@��R�0R+}��It�s��� ��c�U^U�?r���FZ��ީ�C3U{ri�.��37�I]$�ivR�M���J��|�M.�*+�3�M�S�7�ϯ08�+�璚.��O���v�pzn���3c�����L�����N���)�c���SC������M<9M�*U
}>�ԗ��ڦ�׹�K�̗�K��R�Ƨm��;���Y��H��m	E!u\t���ِ���?dy&$���� ����%ۼC���,jÒ�7O h������c{��9f�,�����j��78"g.�I
C�cs���z��8+]-}��MC��w���ބ��#�}��D8V�{�AfX�a/D^��$��i�#�8]Jh{=�=Ӳ��#�O$�UI6�\p���f������7�S|�P�P|�Z�~o���GcE�2iTo�(+`V�4��ǋ�o<�e�$��'_�?�GQ�a(�G�f��ǲ�`��F��[~�����x ���m���M+Y�����6��)2o
[�}L!���B�_-㥣����`x̺vC���4�Sl�z����{zf�5�哳�o	���"��-��P��Ӌ���7j�08j	f)�Ğ�����\��J��&�xK�wgt��FY��)�?��<����8�߲�S B��Ri�8<޶��4Y�j�9{�- ���Ln��nQWF� ��W�>`���G��|^Im�:�̵c,��9cїŅ�+H�.b�}a<� �w���/0�#���vY�pt5���w�O%R��/{�^F�����.�q�Zx����&�m��9ݳ�w��~v_�̳�f�j�j��z��'1�/�"�J��M�HkGƀ7����9MW�UH3���4�#.`
��e���v{Ɵx���3R��6^{����]�S�Z�$>!!,kY�s�h#��G])?�mj�/:�(�a�C����7��ٺ�����f��/��&�(̴Q��˅�Nıa�~��]X���^� �
�_(���T��I���I ���4�"<݅>�H���Ճ�Z��İ͋"3����Z���<L%F�d����I{��e�PS��mQ^�r��t�O."�yr��u��g�d=�Όu�HԸq����� p(�lzR+4\ڪο�#x.��̓Q3���1#�����K��������DO�Uht�D����oF9
��H��)�������߅U�c�E�C��V��H���w���*�d�9����CJ�>  ��"�"��xŤ�1�b���?ߞ��%�Ǌ~㕃�.��J��x؉_f Q�i����]<u%�y���尮+��nݮ�����[=�_�s�ՀJ��n_|&b�MS]�����]*J��ӏs�3x%�|(�<g����@�8W��G�^~re�0�G�K{�R;�k�s�����Ok�)��|�����zBqy'��~���Pu����"z<;z�m.r��Ј�K���$Y;��.��!�qgρx�##PȠ$���_k�AlC�����Ъ�P�.���o�/ϱ��^⳺�+��i(kP�G���UEḔ*�v����ۍ��g@φV�8"����@Ⱥ�|Ț���70���� ��';�k�:�b9�S8�T,@�S��|2����7ig `���e�K�rKa�2%���2������0�,�$��L�b��p��=~�j�bS�5�A��s���M��(��ET���z�"K��\����V��\���qdi�u 2�xyFK�ޗ��� 	rJ�5�|f�Xs3�:��?� 'U����6������3(�Q��Ė� �D�o�S���N�E}����x��'"����.�Ɛ��p�T:*;��������Ӆb�*Q����$_���븶�y�����o��)/ހ@D'o���5q�SQ����@��9Svu��!���&���՜F�m�
��"�[�Fq�t'����t_��5�d�E�^�B&��H�v��ن���h�#�C�':k(���Γ"[z?ti�U�Y�����D��2rʇ�'��`�QÊS�9�'l�sl��xB���+ݚ�V?#3m�K5����|1�'�M��6��w�g�A'́n|�����	��V�	k ��h����W�S�졿!���$	p��p�yX?�-k?@��ȺB�u�uX�j�E�En�\��q���6��5���Scs�����E����$�m����xz�w�g��6m
��E0��{��4�����$��CW���ؗ+
�\�������5������"��2��q��՘��<�'���B�3M�g=�~��(n�ݓH1;�&�>�	ԡ*��&�~b�Upi�Y�|���[�=nb��A�-f��ι��,���s�*�=��V�P��l�*�ܳ�
��(����!D�;��Ay�T&ԩ��|���;��z�V-������Nץ<[�.�� -'D����.��]�������nU�$�C�J�FͿkO��Jm��7>V��B;<��T���:�8�)� �;%@���(�0����N��50 *�2#4�)�F��Z��N/^DbaX�
�2��=p��[����:c�������-�)�*������h\D`U�ܘ�B�+���6�E�T�T��VZ��=���2R����W��6�H��
-�i�
U���8�8�7��ƚ-F��h9��6��b��ƸA���9��%F�`Kfw�# �I�ɣ���E�΀~�0a����V]2Jy���׋m�|p����5t�z�L��n�K��~�澵M\I�bΗyl��b��Y��u��uߴ#�ˣ�d��e�x��֏��b<�s.1N��	����TVğ�������l���$�6�v�Y�6u�A��Q3�L�W�4�Á	�$�kc�^#�SݳB꼦�W�Qqf�Q&���(�.P~�lȚ����A�R���YX�I<�Cw��=>�g�'��}V���z��fO|Dm�q���I�׈�mz5:��T9v��߽����]��Ľ���c]>N�5�?&��FȶZI��,��n-vB�\ �����`���d��CY�)?Gw@�7U�ܐi�R��U�������5m���n2Ŵ��o)ݍp�6੤���;'iQ��k~�B�}x4�շ�U���$S��KA����]lD�����W��M@�k��%�|]q�-�T��>�م���~�5P�O�g-�J�~F�m�����i�h��} jd�>[f�9g3�� �g�\�
޲���T��)a��?�fcL�Vw���Nf?�i�C�^���W\'ޛ��E=���T�4��U�r7>jA��:y#��Юp$Ԁ��`�L|xۘ���|��yf�b�śqUZ��ʻ��u�ҷ���#l���M��[~������!���0w]�
zt-�m4���k滁����C*!� �h�����n�_�)�!ʟ�0�P��p{�k�if|��$�~�C�h�~�p�J= "j�-�� �(�RHϼ�I �6��/,�~��B�v���i�#޸�S.�}�/��&KTh��$��]څ���l֏g��I6�-u�V4 (�k���.GOX��o!J��0�t�)Qz�(�G���TM��t���w��ȼ�D�mPCz�u����S�^�ǵ(�l�	e ஥}�d߅>�
W��?Ƚ$<��C��:�R5���ƃy����u�h�Ca1��Y�`߰��r�(_�5��xQX�ۿ��/D��:���e 7˥���K�C4�����E�3�$ ��L�~�c�&���q�љ���u_y�DkI����x���5��a��9Ledz�GM.k��������P���#��v�Qe������rM�����4�c�l��Mr���^�Y0�fSfje�m`\(��І"� �A�[d	aЛ�����#���K�#>�_ڃ~���t�#��������I��j��%���8����;C O	
�u����'>걩J�t*���m)�1�H��5T6��WRt,12��q�Sy���� �_���5�9�
g�"Us��V=r��!Ԗ���.�p��7�W��#�2�#�gm��c�ǯЋEwF���,S����S�?F?��Nf��i�I�a'����M�z�Ӕŏ���U�ɳs?�XSS�qn4 4�|�+�.1ڟR����69�1�{h�9>�A�������6��b�T��Q�X�mg߃�X�5+{y��2���� s��׺�K���W׫���|F�P����I7�IJo�o�;���l��w|�}M��ߘ��b;P��ɚ3�}�lx�ԧ+T*($p	�
ܒ:�I��$��J�&*QE�����l��p���/}	�/������MQ�H��L䑄��[�tA��-�����Ŵ:Y�F�J���רTiƺ~+����0�!S��r��T����0�M�ܤ�U�6������(���h��Ơ���a�=W���m����_=����O5�#c�f��dè�q��[���'�k}�0����-J>5dWNjp�J���1oq"}31�SHA�d��o��2n[Tg�`�D�ю2eZ�.)�!�B,��42�̡e�)V����JD�v$�^���L�OK�%�i5��U��l�9�v�X�?���Sk ��Q7A=��0�{E��w��;5r8duD�<����V�b?�ֈd��JG��4�\qcM~<�%���W,,TL��?�>laavX���]c"��|���u�bz������Re�\������M藳5��F,}�������)\%�x;�~�_.����
��	�k
g����mC���<��L��o$� ����֜٘�<��(��y�	0�6[������~k8�Cr_\tMjI��I+�ʟK��OS�v�<�D
�X�T�u���#�Y�q`��r����,��u��=*VB�o|�g\��c5��*��Q���6�?�s�b�;�-4�V=�A{|���Ȗ�>�O� �&�Wf/������Z�d����K'1+�(�Q׷��;��g��d���bd�V d� 2%oĊeϐ�"-Y�G���Q��R�!�B�D����(ޔ��I�?N�
�R��
6���1��JKs9]j�]��%��kL���#\G�ީ��+��ҙ�/,CJ����tu)�K�%rv�0�<W[�:z��$_-�=�u��P�S4F��hs�l�2���KG��@@Z�&ٔR���gy�����o������1��z�Ճ��p��@�F�����jX�`h!�������ME�v'���3�+[G���cQ���}�0������� <8k��Ax�n�g�q��j�)0�Cn��]�[Rm�ç���TN��>�������ݣŊ�րPN�$�B&$����Y~�?�b,q�(m%`�e��R�Ա��zf���'���HrD{��
�9��؋��ٸ�bZ��vfWhO�MF����t�Bj����&L|x�s�G	n0�-	����&x��3�.>`�r״n
��ss�n\wϊ���r�V��� �,���n��6K'��:��Z2�wv���s4�L�-��)��CvU�(��J����+�X[�BU=^�N(����\��q=�Sfh�Z8{o�c��2�m��W����M�����I�:���������5r�𧷜W����[�O��hC�
�;}@`�J!U���J�7u����t�?�i-%8�t��N�V�&[�ià�E;���F+��۔A=+�c� ��I��N�Q�3�1���-���l��sz�v���S»l�~�Mx�_����_(IZ� _�I�u&�F��D�J���M�>m	Qdi�Z��v!�;����̤�Z��]�+��
�?� ��7��FŎ��o���Ką��|�3����AU��꽗�h�o��'�`N5��x~O��	��D��2�@ߣ� d�|Ce؎z���?�}������u�r1��D��?`�F>�X׸�;c�m_E�r�Im��$�eQ��� P� NI�㬦c�S���ct�
%_�gVs�/��{,��#���l6�/~v���c���0��ձ���4�E��hbچ�m�إ���3�jf	A�5�����i��.9�}�z�7���L�q-A���h�1�����۞��@I���.�A����H�/%��?/<0x�ǐ`ռx:��֨���5Myل�SS�*�o���_D����lCzM���N����C��֑��ȯ�+�����{DQ�:��a�j_DMĨj��YC����;�:*�:E$ȝ$�c����o��W0y
H���7;qЗ�$���Bf�o�娿n�nn0��O!}�C!NG�{,�y{�t�r�l���<��k�9�/�S�����jP��<�ܽ`�׶��!L@�~+�5�1	l1�loCC�s�ʟ.�^�D�2=�op�X�T<�$�&:�=��2���Ի�x�����O0a��:3���h�9�5��>����<��|�8��]B|�d�+�}
���-��kS)��g��B�O�10��݇5D�hّ��R
�p��,E�q���7lHdI4I~�3f�ǆ�����l�����ˇ��!X\c�PH�ׄ#Ͱ	�a�+0�O��|��KVܺ���T�K��,�d�#�=5(Pз�2V�-��W�^���1���׏�鶥�c�y����w��*�[��C�vB����,=��J��~y����|�L��gn-�.%jK�wu5�E)�(�� �����ǁ��Ŭ�cФ�P�1 M�ZNl*�i^lŏ�V�9�h��7����#���+ 0��2-j)�}�P�����8�S��_�F ��6�9
����AE�t`�;�e�͜��)y���y �!�;�t5E��O��8~]*��c��Xw�p:�v%��F��o�D��x�0�!QM�5��r�}I���b"C1},�q;�)'��Ha d�L�*x��d�	VR�V.�VN(-&�zcj��*���,$9|��Ee�Gc�K�ͻVuᝀy��؂Tq��xq�^�U�D�j���Ax&���k^d�L��Г�Q�@�r�"R
���}�k�+)3:�ڛf�z���#�QQ��$���.���]����VK���^5A򉶢�4mm����.ǃjlB��	��n�Ti����G���"�����QSw��B��u�;�ڴ�#�^=Z�[}5���;�?T��â�RP��PY��L'.	[���mr�~燑Z�z#u�.:�������/жU��	Ym�3�+G�E�����P?��x��n�
r��Q��1�0읭�J6E����u�D>����n�1��i�jEv�,�
������0F�w��3���)i���dh���
:jU4Hӄ듒�ՠ����������(�ʲ[m|�ڠ�lE|�Zk0ߡ�p�r'��#��_�Kb��.gc��x�l�v�Ũ[��*���qP�7�Q��O_�+�\�qخ�:�j'�Dv�R���&�h|�\��!��^#�Lw����08��gI=�V!��H��P�YV�S���Sg(�[�iY�X��=�Sw�k}<7G��V	^�J�×����`ea܎F)��z��v�����eY���l*|�Eg���(��L�"OgI�ۈ�KN�oO�-���-@��O�-A����K�	�	��b;`G�:�LU[D�����T�C?���Q�k�!!�u�U���m�k��I[}[��u��l�o'�B��Q�/��R�sM`$6� [)�v-ȀMZ��A\���U= ��yTY~����S���'�6��b52>����/�Bg�p��Yt�)1a�Œ
�����ѝxc�qR»Y����k��O�֡;�F�&��Ur����Y��'�S�7������5���hպ��_py��"�s#�ɳ�+��lԨ������3C��b��5A���AG���2(T��Y`�3i�ʷ@�_��w�
���(ن!��5�d�g��>V�+�����1/�+[�ϋl��N����(�L4��Ĳ@^��թ��9�CO�i,.d��2�� ��C�HgE�LmY�H���we"�F�����K_���J��S����[$�Y\r�D+P�bۼ!�k�lA�8~]���{�r�����0�NS�
�p�?8���1�J\i�M��6��Ƞ�h_Kq��QRUрk�����V��ǌѿ
[�o�an�S�9���X������Xȸ,�v�����~r�CC�לD�1fh3V�)�2��5Q!)zxTx!�;ʈS1޴P򘛛r�|��߮�IG�ڂp�:��(Ԁ$P���Hr��'�K�����ݩ=-�σ
��A ��B~��W�y;C(.��U���3tT� s�8�j���/��?tp/M@����S�cR�5}$�!	D�F�䬟T�6��p�7\g��d�~�ȥ!���yc�I7�&�x�`g�Z�nxc���=c�Z�f�#�m�a����SkE$cb>��IwEO��t��,�ԫ���n}건��.��a	�W��nd,�3���98���1��V�{t���­�!�AS�tk�����E����^�gIo���[�$��	���
�m7��c;�..�z��U�����+^��ʫl�G�_F�ֵ����.��I��R�m��f�