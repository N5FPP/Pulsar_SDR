��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0��`q�M�'���2&��Ȯ�W�4��д��|�6�K!b�'mY�`��L����Tr�AW��:��3����'�v�WM��=K*��1<��(t!�1�l�<M.�efvH�\��0V(&��2��j�P�cG���J8�|�ݦ5���'J��I��/���� 9�	q�Ϻ7����5������(����U1v����V���W91ƞ�3^:�)e���'qU)�j7#��ME!A�W���$?}��~I6�L�޾�v��}hK���) ��N�������65�n��ī��7�?|��q�a1@ͫ<W]�M�Q}�?��;�F�G�������E��F��Kz�;@H[�:SegD�2z��B������E�7k�l{r�d��aߪzr�PU���|�>~�!�֚ �ߖU�d6oOg ���	�:���fX�پ�����4��k(�ީ�*n'υn�	N�A��5��Ap&�28+�1�r�W���-�f�KYUs��a����qɛ���*N�Z<�
��l$�`P�M�P}j��@��b�Gx�yS;�,��'��yFB0?K%t�(��ڸ���"��c�8�<y��Ah_�č|~�>+S��hb�����J����.�`���ע�e�D���E�HY�L� `t��� 8�.�`[�ra����~��#�e�ݺ�/��s�	Hf��:�D��������gK��-'��������l�m26�׈ w�R[�?b���� ��=��i��T2é�3���ر� FW@�`�{��w�,�d�R���
�O��<O0t7��-�x!�'{�eQM�u�E������Tnh�w=�qd��^�>Q��a_�#3z�8�]�D?�zV��t0Y,Y�d^TG/��_�<CV��|�ӷ��;M+'z{b�e�ED��-tp;̔�*.	�j�{�Y"�b����-r��.k2�����Q:�A�J�$�����";��*%�����/2��V���YG�H�;�ƺ����+9�Dq�� r��1Q�jp�����t8�K�H��(j�+�{0H����;j4JR�+��W���ȃyPI�^)��{�<�͹��|��1Լ� �64�l���!c���'fa�AE�n��hh�(��<P�Zy(��E`-�0[I0��@��>5 �N@��%��:cj;[==�EM\&e����c���u�`� ���GJz��a|���n����c�UIQ����%3�>{�Kmq��8<
ȸ�M�]��~����8�K�(6j��u�s�t6���[��V����Ԗ��إ�^ul�C��a�4i�3>}�\x[sbTM��P��r<�v�� A�[&"W%�:�+���LY߀�V�������th��� _�J/V�uTD57�k���;|{�����+_/��o{͓��h�۹��"
��O_�\����)�?�)��" ��
��E	e�x�P�U[Cm����r�;C��%p\2*���,Y��l5�u��D�����:��ش�-�x�|g�@s��S| ���w��H$����^F�G/gv�=��Ҝ�K(��%�=�p �fB�s�&�u�;�y�8���"Eg���7��O&�|�����4-Қk�w��_^�D���g���A�,��� co���]������ާ���*@�ϹM�q���?�-?�P������i#ު}�.�\���50�|yx�]1/hX	j�����pG�M�2�<֙,���_w��5Ѝ�)�F����[���݉�&]��,���7�A�����P���j %��	����7HaDwwO�Hfc��kT*+��`���>����kl*0n��;��y� �J�d��������J��y��DUPI����c�a����-� ��m3p~9���լ��<�h)�a?����sL��ҵ���M��O�fS�
n83
�b���4ecƷ��V�\�;����~QK���nC�����C��&J]/*.=����w�:D�����q��+(�L�[F��J+	�s|��D�86s�At1XE�Y��2��q�� �P\26YSå��4/��VQR�����2�T�0�5`��W>s���2�I�G4~`J,�:K�2%Nn~��Pa��
sQ��#�A3�"
<���Bw�9 J�Z0U.�1�0g���@,2׼�[W�W�xVio�n�����A�u������',+ΊhѬ�++Ȍ{�'�%���,��[+,��ܶ��y��~�rc� q��I[-LF�X�4�s-)���m�0aTnL�����Mo�}�~bej�3���d���{�ӊ��y�̴����s���;[�̉�0F<���~y"��s�J�^�%Ѫ/�V5\���%c�L<�l��ºh���%ʖ��;�`�l���$ [8���YP�B)a���h"c*k^���K����TzrS���� $��}�I���t%�C�60L����Q�bd��������˯�P����n}�j+`����֗�v�f��Ֆ ��x���Q��;�ه��&o�� ՜n�O�ދ$���X�#�VlC�;!<z˔ ����,�ɵW�
���b�0K[-�'�	���9wq�Fg�|z�i��C #��x��P\��<�'B�f��&�p���Ab�̂롟zS.H�cY��4�nz� �-#2V+ȗ c�6�Y���BˆRJ2Pg��v��z�
;ѝ�.���Y?'N��Ll%���l���;Z��������5�3����bR��<5�Z�&	-"��#.`����i3���n�P贋���mfY�ݪg��'�L=-i)kLi��F�Uu�Oှ%�����e�*��kΎ�
(�KE琒����6|�֒�2�gk ��P<]�Ā�H��l���~r{+�����X�$�\� ���fsH��}%�0Y�Dh�����29��AgBUB�?{�+��)"�{�B�����~��g#�T�a�'G�G.������w*ƃM)��r'�(�½ИM�d�J*�_�L9jo�"��Nyw����w�R���Ժ���^�C�����Ov�+�d:�(�������rD����հ@��V��#�c�1���̑��W?��K7�+�&�_���u��\f�&���0�~y�7�=/l܊ak3�Hj��=(�M~na�4a�CG+t>Y�6g�F��d�جx�W�xfW�A�J𯽩mx�|C"o3&\�:Br��V�O�q�#A=�=G�@���K%1<�}v�2�?�%�
���EL���j�m��;,�Q��o*S���׏��a�*ܶ��'[}��K����} ���_iӤ��tPbHF���kƉ���:S�rz4Rb*4�4��"÷d2��^�Ro5�a��40<1H�ikU��K�}i#�1�KT^�j/&F�8+/;l�%��s�R�}o5HH��5���0��X��cd�ƹ��^3�j�ֻ��F��G<ܶ�Q���t���K�{n%t�j�u��Ie׼1,?����.�(3��<�i��^a3�~�#)�THV��WG>\��AM����.����i�8g�X����[�)�(�&j9�l,�H�Z�*���^$�58�������ȿ��@��)��IS1���5!u�R�K�c.���yB��k��"�Ԏ�YZ�^be�u�zW=�P� 3�U�J$^G���ka?�JUg��
�ᗓ��ޗQo=Ӝ��m'���}.��xM�'=cU�+kߘ��
Q�D qT��b�Ɣ�J���.e�gyD�0mGxL��Y0����`�}zgz����rIe�Ȑ�IR����ڇ0��{��i��"���w?)!f�]�[6u��s�^=L̘�U:�@s���/��IHJ�QP�P�t)*T�7��Pk�D4�^���2�6�]�h\��^����Zē.�UF9����&�O)sllƤ(�^
�FF����j�|m.��4!���{�_��P=C܁�����9�]�ILa��7�A�Z���ҽR�Q�>�pR����e� ���d�Z ��g�B�0��\jD�|ၔ�qCKu���lj8�\5�� 1���#(�]l lޤ�`s�Q���hb98P'���IF$I�����n�S/��}�Z�5�`��(�S����d����c���b�g����3��o"��j�>��u��t��3B��u�u"~|P^s@����8r[q��f �jh<�9t�Y1b��C��^	���M�VEW��Y4��!M{�������ܮ�H4�P��Jݸ�2�Mԗ]�/�x��u��.�"�0�.�>���7��G'�W;�Le�X��ua-M&�� ��UߝY�x]5ɋvq��n�H���!��X���±�ĕ��76����;�Xn��K���؇<#wQ�����mo�&|DSlL?&@�syLV^��Add�t�R?�7z��	i9Ŀ�nP�==z���82�r�xp�8��Q�"�y��:p�m���m �L]<\!���gY;�q��Fys�
C/�؇+�WC��ٯ���R2�<}#�J"���^����&����:	�*�b:�w@�Y��m2D� ���T'�~IX'���nd=��+��f(éx� ��� njM�����>���D��;J�cl罴�(���V"K��ؠ%Zt=��X��$J�xf7�QG����zf�������@ne'a��C��
<�P�R���8���Ks�Zi�/���V��:�/輿+8�Z�V���ELku����7ύ��}ד����=��g޲z�W_�4�U�(�Y�_�u�O�HPSp�0���	;���>Pe/+���tU�ᄴR�����J/@�;Ւ�@n�#D2ݤ�<�B'S$:�U���0MU��1XX�p@�Bcsl��n⣳�z��g�v�Gp�}s�T��a�
�������x����m�Qe��^�k�����ڨ�X�j��1���˪󇴭�|�	�1�Z�h*�ɂ#)l�8�ф0�b��pVT��;$rp�'.�����|�b���8{������$=�(~�2��<�8�C���7A���U���ez�'�4������F3�q�;Ӵٹ�7���7H�Q^�ʛxE�PL�a��M�� ������(����1��p�ԙ}Gf�ٟ52�s��W�����}�Qkn�����bz�/���vD�*Ia5��]��\��nb�����V&.ŰXP�;�/�(����z�-���rϮL�Yc0�(!F�ь��Ը���o�|3�~�V[+R�$�eO/R�^��:����?�� ���&|@���q,H����Kvkkq!|zڑ^؈��r��R��� �(m�B]�:e Һ��W�v�!|��U��X̿�����R?���Nߎ��|f���[��>��c�W��AL��m�A�������W.B���e�,���%��U.jz�5礗t&Qtԙ��(ʲ:�Z���bA8�ݳ���.��*B7 \����㶣7����$\- ����Yj`F�2�T��J�"���$tC�@oI/����a�1�B�#	���w���t��D�5����G��g>?a_%�S՗@�j%�:�����Y0M�s-��w�|.�Ѯg�vPqK�l�ۮرSH�K���kD��ay�wm�8�<����.���h��e�Z��]�cJ��N�ϙϞ�	�(��b��e�U�2�ɻ|i��p���1� �/���L�|9�\����?�`!_��^2%t�}\rb�EÅL.HkL+�f�,CA��.E��|�b�f��io=�2Y�{��0ܓQ�@����"v4׍�V��B�+:�X&d�a!�pF�=L��0]c��ms���"�Uz�y]�O���&y-PH�T�|����Ft"V�>�܌]�-�`t�g�P&�:�W���\/��Z68�#��x����(�����zC�������(���x�8��4b�\�-�!���ѕ�E|��*��s��dhc�x�I�:��� \�i�a��