��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞX�e�(����eZ�0 jY�%��{VY9?�C�><�f儧HJ#��� #�G��y���9T�3}��&�Ѝ���*��$��"�s�d^s;�n�BMg���FrQ���X��xa�ji�I.5ny>�P	��~�ͷ���|����_iD�\S�#�Ӹ�Y�M���4]�H9�@;T��e�S���pz�&:h���4(#��c!�ۗg��H��\x������p�񅑻�_���_�*fw���p���.��&����x��ª�zJڌ$��b~mѼ>)��V ��M�V%o��ٌ��gN��[j����-��m��o㵤(��Tַ�q8����?(�L��^�O�=�ii�l	����رQ1ⵊ��=�O4��rX_qNC9�c�1��O����7zi����E�;�ؙ'�5��ԗ�����Y�j�����K����%6��I�,h���\��9Ҭ/��pM��j �T�3�҄���gF�^ h�� ��TD� MT�">�v�t*�21ch�w�:l7��@����y?� J'9OpWBC��x�]DC����G[q۪�L�R�6Xz/�����ï�}e�>0�V&O�)�;�k�p��^?��,�ᰉ�=?���ǈ՛jњQM�J<H-����M)��ȹ��?�7�Z�� �K�
%H#� ���d�{$��"�\�𹰀�d��vt�s@�Un��� ٱ���at�/���%�]Q%8��89�n��6P�Qc��sL^��V$�����6w<�ᶬ+�yR�sO�S��Ie�q0�����k���S����=�#g�=ox���b�ў��+�J$	V�C�|��x��u���*�_8�;>������b������$��p�Y���VZ煨�����T��ṿ9\��&��D"���J�
9:��U$��Y&5G⻉�pQ��<	�Cm�"���Ώd�W��Y����f�o�ݾ�ظ���4�KylGo�I�Ň� �7�M��q���OFd�Nz�E�ԁ�ՅJq�t]�X@�r�cc�KpZ�P�z�2c�{g,��#�	wsS��qm�ce�b�t�Ë]���P��F1���~�g����!�ؘ7Br����PO h��p���H��r̈́�b~�{!���}�2�d.������1��ޞ�"�^�q��(��Y�_���>�3`����
�0�l���� c$0�{�gWר����E��bc�Yw�(���0�;9�d�v��ַgss���9\P~`�+��c1%f���ya����е��xRï?�[�b�\���:�!l2�Ժ�F�����kw��"�
٬2�R��T:*Bۮ*��aa�I�!#n7��/�#���t�Z9�|��`rZ����/��/��EiT�l��P�tvmȴ���� J�R@<�iCFm���9���^���L�v��R�!���f�DEw�&�H�'>5�|�{f[�j|_�{��_�R�F_�`1����{�����l�)H^�Klb�%�=�S�8H���(�>�Y��T�#�z��Fn}�?��a�$E����bzq f�Y��+����+��3.�Z��:M!�sj�D�l�T9�7��&�@˩Z�����8>�k����lC� �T��7e�3o���������_��Lp��?%ǽg��M����(�ɼjy�;~�ХPo�K�V�gh����Si.R�j~8�÷B`V�i%���Dm��m����B�aIA$M0Üc�r%Q�9���[�X:���:������E��z-���(�J���:Y%���]{�Cp���y�YSJx���pI�W��r�pD��U���9%���̷(�ٕ�8Y
���ů�:��S�$�)L!�W}oM���j��� �� tDc��$W�i`w�6P�m��~���%��"CU��Ja�O��͇��y��L�%��a���3��J�BO���