��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� f
���O�Q�h� 1[o���zp[ �c�p �2q�:�W�9)�t�(�����1�B�ps�n�ri�s�R�ng~r�t.��:���\�d�@������P�R�;^��42��i�i�h���71���e�9��9��X���z�]-��a�g�g���w�4��i	�p��� g���؎m/�/�1��~�8V�;�$�5��V�xo%Di�%J��� rA��/h�}�	&�+��;��+�����hs.��,��ӌ�*�:6 9N'{������+�q���a��6�hszx�ݒ}�����_��9���*C��x���P��r�*�C���¶"�[fJ�c�.M� �3�ls	^�I�i~_G�X,쳳�V�U>h������.`e+/�|i��U��=��dF+n�I{V�Y�����azڬ���_�r��7�}P;�}{��+��,��AN��'avVhO����V}����[�����.�*���Q4�VB��q߻$�	��
V���y��35>~~��9Ƹmn"��)yA׵X���~�TO*�ad�m^�J��
O��f�o���sM��?��@��] (9έ���.�Fr���	6D/���e�L��Z���t�k�'�`xK4���ܛ3�/�d-Ny����Z#ŧ��:%�Z"�R���U���^4r?��4��Z
s�	Ȼ�#��x�O��F�-�⋀��a��\�S�����*���̨������j$��ʨ�)��i
Uݳ
k�i�?]'+��I��hk��� b��=�qy�Ok)���&>W�Q��ˇ�͑�/��es~�;%֫S� �f_�n~f?���Ӏ&\��bU~���Nܳ֏�N"+OS�,�Q���g�\���Kۅ��G�`[Cx@���O�u����<1��+����w���00��.ɲ�sP?��47T!�[e7��r��f��@&�wT>��z��,�r*q��?����+'�i�{"����������eO% α8j����o�B�'���X�C׃x�Q�h�تb{��i'�>'��i��b+�b����>�t�\Ty���@}j�r�F�T�㻟�-l���_zmA�$>�R�*X�=�χ�6��o:g�O�P
V&(�"���Bp�(�K�a�ǰ�	4�4�=�Β�]`��� \g���D��N{����z�q����_�258�j���<8a0Y�i| ��z�<�>/)|�	W�䡯���,O��C��~�h�!�.��=l���=�y��y�ƫJ3(x��I�S='[����C��gߝ)/�PGek�d�.���Ng[���N�Tm�+[侮��#R�Pf�Dt$P�����0����+iٞC�\J�]�6`v)b1#S�\ԁEt�p�̖�L�-[�W��I�$�+oUYn�����;{@�%*�|�U�9�Tܲ�2IK���˝�"�'&�76�A܀w���d���PX *ǖ>�{==� _�4�]�`orӏ�l��i�RMT��'�s�qx)��ba��@SN�æ6cw�����t�M�Q���J�롰)ʮ4E��ޥk/CK4���\���XRXv)�g��z-u!�n�L p��{���=7��և<8�;�qX2A?���lQ�'�f"@ ��`�S�.Q,��S��X��:+�G4�jCEW��ܽW�k^9�Q��:+�ٟ�E��'��s������j��r�#���YB�sO:��"���X�����/Xtg��&*Wt�۪e���qb]�~�nw�S͡��/ ��Z!��`Xu���gI�����6Ŷ	V
���2��1�/�E�{���y�>K��K4�]��x��
�;L�/E�����ϳζ���o�0������k��ߥi�l,����R0��_�r՟e��RI��1��ۘ���FT��/G����{�CE
,b�喋��*���*�9��i�軃y�������*:}1Fך��)�dy(�g#�X���X�TO�-�����_�
La�MfU'�v�6(K�l�N��)�aG�^(��G?���&�s�|'�0T�)@��N�7hWHmR>�g���K����B�
�.7\���D�4���ux�>�M���(6��\ݹl���˺��.a��P�;�<_���w���q=������g�,F������)S�_x��pK�i_!5��D��.�}��k�d���C
��P�7!jf��M@H����!��?$ƒ�0b��Ůވ!u�*i;t�{��YF��+�Ɔ�̯=j���K�?�%$!�/�E��g߸c�
#q�f'�G_q󓮆D0W���i�9KB�|��I�� ���K����^6+9�ĸ���j�;L���Y�8�Y���Չ�r�j��.�����,�(�_�w��1cT1d��e���ƞF�iI�#���7v�Ux�?�+u�#i@E\���Pk\�kiZ�s���N�p�r?�}n �+�D�߽��mV��l4����"��~�/Wρ� "�u�B�|݁�d�╰v$q٤z��B��I}���/I_I��Uէ�w#�3\���S%[N�����CɎ��oLu�Ij��5eI>������C��/݋F����[< K���Ѱö�
�<�M:���a��h��t^ s�}��M�8�j�P-~>�������y)$.�rz9Z�W�#x�!c�~���<g+5S���wo�
�l��k�,s6���#<�6�]le~��]Wd�ir��:k�`���ƴc\���k��6�R"0�M�ch��Ɯ��+6�2H@��/9��NJ��橁�Ҽr�hZiK^O< m}\Y-��0ӧ��m r�7%G�*��9�_Q���B�EH�f��Ĝ:�QS�r���� ޚ92�-'��Vf:+_A�L��&*Їo���)t"ׅ��jfM���SYM���v�Ҳ&[����#��vpCkg#�Y{l@Qe֒�!y�&:4�Z쯃!��v�1y��\�E��G�2]�\Ss4�c�˘�ò@� J鵣Q)�0hw�$��dp���=�FX��d�NR�X�:�U�ϓ:;�ދ�k�ޞ����e��������u�h�o���Fx�m��TI���̄��Y�ι�2N^�y��C�|��YuUWK��arǋ*��:�uY��"��Sw�ma���k�]���`����%!�O�H�`ר����@��1Aq�F�ʿ�u�-�~z��YûL�Z\�oP߰w4��t0��ғ��9�lh���/�
����F���YD�.�3������+�5վ�?犡*��zeQ}�tqu�^�(�qq��
���{P�/�laq9b�q�F������gN���ݭ����?�C��3�IA^�:Xg�+�%��>�ti��Ay�	�Q?'��|~(O1�X$��M➫������H��%8q�d����ߡ�?�r��u��)n�C�C�G��A����l�[�2%���0̓IS蒧�̚b���<��w]���?X�hzC52�@~��<���^BJ`��\x[T�Ƭ�RC��3`�I� ���#c�->���Ʈf�:l��'��y˓5I
-Op�a-�B�ke��M|�2�F�ϣN衒�6~����٫�U{�V�l�6�-��R���VU+y�I�9`��פ�'D6�zg2%ρg%���'�H���������2�T�r�ᡥM����)����hXc}2s�\��r�G�Yۚ�n��(�x+����	�ɮ<©_H����AGK|� ض��oT�"J
]�Ęo����@A%��#������O�I�P���1��2�R�t�hhQ�8��U�t�t)XP� ��:!F���\?mI�UX	�ր(���L��iՂ4�6�TD��+2�zXjш����z���e�ʀd�No#����s�fP"��;�\�e���˯�_B>OSO�;O�
����Cd@Fj�f	��?�f�--Y�۩c\�]k��Luj�G	��v*���ZMU�v��S���o�I�ę�n�����'���;���k֩a*����A3
S���[�f�MU������_߆u��6�[��/$a�B>`J�&ށe�N8T� %1Vϣ�qD]}E\�SfR�{[��^ @=èK[�9���8��%n@C?0�WF�ul��J�S�:5d�U��h��Q�{P����#���V���
����������I玿��}e7���L������i�
�#��L���r���j9UF1GC�mas�N�&^ٍotH�Do~w���OQ�vh,R�;�̢��� 7���7�������B}j����Ǔ�d.#�=o��>ȅ�^A�[���t��H�.N� ()��:~�J�s喥�-�X��X�/
�2/ݨ����4ŷ��^R��
U��0@��{d5V3Wi>B> A��or�����8YuD����4d,1�@,.��A�b�p����s�i�6>�Z�~Ǐ�6b�p$˓�~�xE�DV�}p�)\w�`����NY^Q�m����t1�;�FZש�d1@���tGo�֢hx�1�I�]�
7I��m VqT�o�n.</�&�!��C㽼�����tQg��@ ?��=D�������K���qoQ��>�,�ǥF�{��-��YM��ߖL!��p�g���<��;���L�Nʗ�d�j��Ƈ��+[$U������hR��d�����>t����mV��G�=�͗����l�o��#��oi6���Bn0'�ԄபQ����$JϚF�!Uh��F��d6A K6�Mڵ ��U+�k�(\|��^�
�R1a�b�}G ���Q��2q�f'�� �W�:ı9�~�d��k��Ǔi��C�ߞH�����c��7;L�i��	%��� �ʮ4z� ��a5�!C5#Z����?M����X�k�[�`q�!�lrp��%:-�i�U'��6��+if��I�y���_|��]�z��y���_���&�bH|�6-�&՗�4��W����%��Qeb�þ��Dh�u����=$�k�-Pz���.0"�l�m�*������j�Cp0�3oR��gɈ�8�Ѫو#�y�(�H�麊n�'���D ��V��x0���e�GSu_1���Q���\�k7��0+|�ೋm��"(s
6��.�#�X�o���������e���WOO*��7�A<"��YV�Y'��H��C����b�4�<O`��'sf1g�p3O�o�i�ۜ,�X�)3I�Z^�����&��)���v� {S�=�:�#�?�mX��r�ͅ9���;٪@T�!B�A3+ͧ4N�\��C]�Q��p�g����Qj��Q|���E�8�A.`oᩁV��9�"��*���\��3>�2��#��iK�1��;E�\�������	����O�ʜ�W�s�`�d�\�w�5�7L��;۔�GR�(+�3��5z����/� ��I9�q�r�{A\wN�7.#G�Js
�j��~�FL����E��w�q�(D;u����<�u�7&�=U��}�I�|"0Dl�8����2l��΅�d�4��/��[���C6��_���
���eS�\x�D8����B��7�{$[䢚�����\�g��4oL�E��x��iz�lM��/G��W��v+��f`x�p��wF3��(X��m$�w�h?f�!�*�Ƚ�f����1��"���t+���z+�U�r,�u%G��i�_o0[V�7�4���Ϲ��
�$����u��
J���-�9���.D����i�h��A�3�B����W�S�}$��9JD/�y��jˁv�H�?;���Ӂ�hS���Ƕ���Ɇ��@Wv��D3��]d6���ѐ�����SKE��ΐ��pO�a�_Dc��2�L?֐\��ޥ_�&K�#�s��fZ�
�"�i�]��[��t���h�u���`S���f���&i�&�������{BX�[~g�ub�u�G�-��u�Eqy&�lWc��;빾�AJw:�q���;~��8�m���A�w���<W�
��L1��	�m�!0�J�Z���a����LbF]�Ul�t�y���U�<c�E��Ϝ����:CGi���*��AI���T�3��diEJ3��-�ǧ��B��mz%�zɄ�W�������F�pA��-���������L���WOU��0�9۲V�~
`�8T�P�p����]}��Ѱ#�
�O8P@�-� ���J�X/>��AkƲ�:ËUkF�ŪW��[)������+�U
�����fW������EL��u������C�"YiCi�Yq�P.�|V�=�o��:��n�f$��)ie�q�s��
*�rY����#�g�,pE��0/�c�1�����A6x�k��<T���̎�Kk¬��DªJ�Wi��p��@��p�����/�|��9����#R�{'%�>;��y0lIM5��Ȼ�����(}��w���U����N���v��MJ��z̸�䖜��ݔ�E�c��/$�M	��2����\"��ݥEt圇���B����f㬄'o�����ё�ze�E��M}��e�f����@wD��&����!o���at�	J(��q;��c�lq�ϧ��k��~ ��)�Sc���h�	�~����3=YŅ*Fy<TP����7�?���-A1�j6�?u-�D�=u���z_b<�3>����7s�Ư��«��v@��0V�Tq�z��!:׬=h#:^?~���:�*j���e���Z���]u����i
]�6��4q�\ӺY��I�ӎ؀�\6�a�C 
�	�Y�,���$U2�8!H�g��(���6z9ͬ� >M'K��9�4#>���2yBc�����]�֎�Ć+ռ��7Q}5$d�D�d�	�N�M�{�ND��T#�!��'�R���?����=�P됟�8�X�Xo\���5}x�t+�o�Y�/+w��&���߰�ި�����2`?��/cCD�?g��M����S{�we�L'���K���m��At���!�;|\�)��8cg
�%�Y"-V�.A#��K�kڼ; �Ic��?��r�f����"��QT���9�̮t� M�$�qN!��S
CSF�1J���*:ncH����t,�,;�N`���c<����M�o�U?_ �E��OP{s�idi��k���X�B5��.�֠�O��Z��������vko7�D�L�����+�¶h}����Da`�#=4߳���O7��D�}y@��M�
���ȳ�]��bj��t�ӈ��H����\�c��`�oW��_���IB;m��V�к���K��P|�&���2 F��Y�FoS(4̢f��OrJ�a�E/�?�S��c�)�x(y����i��\��{�64��0!��;Qk�g����O#�|oC����$_)x���OE�[9�g.-x,�xFk���X=LO��NT%%��IcS��a���B
63jҋ�|�d�1��b���w�$��c��E��VZ�j���~^KI�a�"�P�֋�#3[=uƘ~�rc�����Q��ǻ�&��L��"��74l��R������`�o�ez��NAt=r~��)m�	E�`ug���a�\F ��,T���vI��u������v��oQ���GT���&����{��]�+iD�T��VV�1���V#�KO(zL��T�s����[��"� o��j�:�#q�.[���HN�@���믿v�0CjMn��ʋ��y^ֿf4����d0X�X[���yB��-:����ZgS�'O^�41��%O�"L��
l��⽴/�� 7n�̗�����e�T�{l3<7��->S��
�@#VƃU�Cbi�������Q�	�K=tK��_Ɇ�Kp�Ҁ�%軞���,PD<�/lþ�,�̌� �G9b�����i�u
8��s2
���%p���PG{ h�໾���w�=&�&-v��NpW�5mX�a�t��$��zLL���@5%'��
���ڒY����gF�EۼV�3V��n���]�nL�8�����Bj�� �
/��5��j�E/�`R�l�@�>��"w��#/��8P���Bd��l�4̭D���B�Gn[�~�;N�b�45(�� �^ڒ�Ja-�EP ��o����oP�
�Tp��-��6��`����5��*��Wl��eg��1Nk���b@�������05x���{/�c�7`o>׸&5��)�W)��˧�8XS<&4��9�sW�	�~�c�q��&�'[�Z �z$����Wqb��ɭ��,���²=�vO�o�/�X zײ�\���CF{y��\�������#I�u�����y��Rq	��k�,]�X��/0?<����k��j�@V�s�Xqv��8@�E��&�]����-��d�	��6��P�<�&T��W��Ґe��I=W��l�f�g�D��n�\eq/߇SNѻ�g�aKH0O��f���6ĺ�f! ȶ����e�P�m��z�r�����Lh������Z��i,�1
1�T��n��aVyu�=��C��[�q[2o�.2�'8��l�*�jJg�ד��0�x�����q3e�{A'.%m,ؙ�H�Uar�Z��������V�P6�?\P�J
V�p7��_�[�,1���Mã{��ع��{��n{k�����l^>n�*�d�m��1��M��̇S-`�>���Ӱ}�}�"��EՅ���~�\�gϭFkk1���oFzI;�>�:�0L�O��g���T�#����ɿ�C���Do=k���it��6�.��ۢ7Φ��OVխE��X������^�¬���	�F?��BV�Na�T

�Ƹu�x��l�_��g%�/#ԾR��WO�#��*�c��_��D/L������Y���`,�z�~n�+��G�Ň��JW��x�G>)ݕʚ�Z�k�%�Bg��82* +��y�ᑘN#�w��~�p�%��J�=6/(����?�TR&���<sG�IZX�nڧQ�*��d.OP�L����@f��`��՛�> �68���+Tȋ�*(�|�{C��w�1>�b'r��*�k�bQ��^�E,��R�C�=m>d�������/��};��g0��Q��5u��Qaް�}]�Q�����鈹V>�#F����f`�3�ҌOÿABf��|�E��<f�� �����?*��&��B}{X�V���{����!빰�Eui�t��ۓ�s&�`����~���6�(������@��֠�:�-��y�⬫ِ�ﻟ~��~�Li^"��w1��.	������
�݉����ڥ� )��}��)(���9�M ;�w4�L޳�<d�T�����_z������\L��Ѷ��{$�����������:�C����S���F�F%ȭ�GL�e���b*9�D����k�_��wM�����(���I����Զ�P���u�ʭIA|�ڟ�\��b� C�h�g���^��*y��w�sܳ8%o�_���5�R��P뻎��%�E�)T<�NY����)�o�vu�{�ͼ�T�%P��D�PY���@[��;��7�)�M�!i}���[�f�!-z~���5�� �4f9DvJT�Qy�T�9����E�:9рYA}8�*�т�Y��R��R2�ѧ��oe���h��__r��0�&�d�w0^����]NK�?ԝ7b.�:7�ο�^���2Rx�3�;B����y�r�AA�����)���q��HiG���k`��nb'PeQ]T��̮�/g��(��)'�5u������>�HFd��$�_�8���v$��,��s�nGJ�������3,�UV?b�b�՛���/R¯&ȅ�8r����Xe�#_޼��h�l痸S)���; ��O�STlb��r��MW��[IS��f�y�ٸ�b~�oR�=��������:��}(!V�2-L|m��}>>��iX`��j��	�xw!;��1���<6�l��{��x���1��_�#��*j��BX���J���㱮�D�o[=�-�O+T3aF�GI�ի�~�+����헹�k않���#Ȍ*�[i���q{Q�͹1�Sq���LTFn�Й�5�J�AX�Q�Q�A�+j�dh�Vr��j	h�:�m(_�X���^�%a�v^���v$p�� �(1�M�dL~IMFJ0�u�����"6�׏X�;z�����Oc�KB���A�p"��CD���t\k�kbȱ�52H���MBbd�9&�^�3F�����`E��),m��㤯9Rby;�I�ܕn���^|6���W�������˨�z�>�Y��(T@�f<.��C6=?�&�s�=�ڝj8^er�i�+�����m�P�TI�bAm� �`;�U��K5�Gf{��F_���'��8�n��3��\Qf��^^�9LQϼQV/	D<^�����3�V�cpܨ5��Z�D>F襭�D�m�	����G 3Dp
��������%�+۹=i�o�}'�q��C�Uq2q���O�_�h�,SH�s2�ń�dT�3cM���>�"󉹋T��F�G}��!U�Wm��Ų�1�:�4�8�	���SG�S��c�E2�Ra��w��N��#���wy�_�{���e��r��^��f~��l��?������p�MO��X���ݤ�@��z�ç
�Ů���!I�=<��ȹ�$}�<\Ҍ�6E�BI$N��Mm�S�wh�Z���3&��@7Y-É�V����`*+���P�<�Y���u62�I����̩�i�#Gg���W]]��m�/��$$�1��e�� �v����J?|�Zς*J��_��Fu�=�-�N���gƌ�κ3T5�˲���Ӑ
�I&%��Â����'�vIo���7�;0r�'`�u;��Rݨ��r|�}�<�����9��ThE����FS�!y��@��f��Tb&u�0�^��c��f
�p�!1�UQUֵ��ED��+	����iY�rrqCQ@�8�/G��0>��#�s-<���:�4)h=�yq���T�9U���E��P���A��WtYқTy�F"d�3��$O��Ƅ����t��� ��Z�U��=���'�q�(�/�
�?WJ*�Ѵ��p�^M�1�0���b�^m?P�{m���-ڨx�Ae|��ѭ��D��2���j�)LD�ᬈ��Gv���gA��:-9i�g��F�ڃʳ��j탬ͯJ �^�� ���l^壍�h���ŢߔLan( k���Mk�1�X{�*Xo�Uٚ���i����������I�im)�K�*l���`�h�l�0T�p�TsB2o�����w��@
�.��+�9�q��@��8U�+��Q��hVq2�|����R��dzBi߶�&�˜2�:@�7^=�Lz���l�6�'��o��bgn���K����8<;�o�5^����R5��Ұ<,>[�MF�6�hK���<���xKHr�/�����[j��SVWM^��?tխc̅�0���;�/�C�)��GS�S/����P�N�;��v��'	WjA7��~�5ԫ��%���G���m��3��^���_�[�aw������y���^K��e� �98
��u��9^a����ර�<�}AX�;g�e��˰o*����� �v:�� M���7�}�،-LE��ӳd����Z�'�˙:㸠�O4�<M�d�F��uִ�9q*�7��_��d�/����=�Ȣ���\��cT6���k�����Y�!Z�+IK��k$ܢ�f0��}���{�'l�RkW;N�� ��}���x�{����߂s�ͅD\�`F��J4�t;u���@c�N��J��DL��%�hd�}юՓ�l�~t��c1P�>3�n�0E�Yؠͽ"U�t��$Q3�9���\H@�0((�h�	���,I#w��'�xs2�����V�yVj˥"�)��*����k��3�S�[��bWˑh��Fؚ�7ڭ���N*b���(�g�f�|�#��֣���ڎ#2�����	a�"
4�g��{]Z��9��4�u�_�	}%c� �b��6��
�, ��3���꛿�yG�^|<ŵ�f7ot{����2KEj��f͟�o9��D��P�ww�Ab�k�{���rX�H�G�\p�\���g���K��k*X�����60��)��	�<W�Z;c�V�	slk�j�t��l�����HQ���j�jn����{ػ�����{����.@c:-<�k'�=���eʑ|��!Scc��</f��F�2E�E���l7���nzЇ��pS�5�� ,�a�SX�綂t5d&w3ë�(�<�>�t��Rx���D���鑏� ����T�T�ɻ e��Y^��2��2}�Q��{���h��߸�]���y2֔��f�@q�s�~_�>'�M�H~��^9?�Z� �n�(�b���(dQ�+jZ�X�_��H|㶔!��-�OVx�+0��_'�{ {K_س蠇�U�Fɩ	�;B0�Q4��&n��y��I��?�LM�s����<iR"	�bo��qH���*�j�����AR��?-6D�^���OK�����	��p�N��ڻ������j�t�����>�n2>C����H�J*dD�q�q$Ng��x��:�����gGd�]neo�V)��ַu��	��=&���kj��m��?a��K�)�������╔�5��k:K\u�N-Auu@s�4� %���6dIvǛ��¶:.�>|��p����ݬ*��#��?���mP�Z��n|���j�n�Ͱ<Qe��5I=@m�Z��m~�,<����ߣu�z-E��xnؼ��O�=����Pr0�ŉ`��Y[�ˆ�T%�r'�_3�DI��;~�7�lE�w^�}�v�w�=:,w���y�ʋ �L)��(��1�x,7 2C��SSg�e�����H�W7���CU#�~��)����6���VQ��C�zM a��}�H]���[��7�ⴿ:�yQ�
(� �����m,���ՁG.��*�@�L�S$o�e"�9{����LA�۸��2�r��!����o�0�'0W
�&t(�>S�:"���<�6f�ql���r-�U�<�2�@�η�H\"+��#��d�1��}�1��'v�el�K�p�����%���!Mx�\����0� '���N^�� S-:`8lM:��P$��P� .s��~t��1��@$?^���}�@�*cc�&�cRc�o�vm0!-��#۲�>��e��²���*V��@4B,��R��ʼn�ZyC���Þ�++����WR ����t���e�D���^�~�،ê�m|�}�/0 ��,��6��[�&�wK�T�h�TrI�z�B�0{�C?9#� ���qU	"'�Y�վn9�VS;��W9�wEny;�/&q�c�7p����p�
C"Zu�S�Q8uLy$Žn�]�6u�:z�'?Hk�S���RŖn$"�*E��J�}�I�3�
�b3�&��_u����*�����D򘥀a��IT�w�:�^�Et���Aex��O��#�5�i{W/HI�J��*?�D���+�*����2a� �	��Fu�{c~���0f:\���u+ο2.,�i�)��	����6ƾK�G�Uakgѽ���u��Q�Q;�2���+�/�nmKL"$�J���@���b����Þ��L�?�Z��bN_5)�����à|�b�J�ŷ2�E���#r�����(Pe�0�L�)zӛ\ʊ�1����b4�����CLo�#���e�߅��e��f�(�{�������l��z0���L�0�$\�yQ�#v�o5h�:yJ۶S�Pe�Q�j��h���;~q��)�\�4���N��! �@t�ވ��ﶄ�T�Q�IՉy�Q������9�W���gK�
k�Y��$MC��V��꣨�}R�� 쥚�nT��K��3sk���l�K����f��A���*^��kP�O�|t��4���������<�yT�tv�?Par���	i���G����d\KB\�)X��7mh*�?i0��|w08�����-�Ѳ�L��p�u[ڧw ���h�<G4-yf*Ϊs��I/u!�#+�ۆ�qI���*�Wd����B�k�a���a6��.��N��ѳ�Aa7�����4x􊥝S���ڨ�\��5���C\Q�����ߖ�3�s�k�e�n(�/f��/�<�L��ɵ�<5�{u��7q���Hxf�!�횗)��'����,�:�π:zaO>�����V��-���qQ�g�R�DH;ؚ5Z������^���j��4��ή:N��?QW��<����F]tmC�.���5TUYѵJ�T�FF��TDyYNH�����e��~u�|�Xh.�HB�� ��kg�v���������Ef1�J��$9��\\Jp��u ��_J慞c$�@�|����F��㹊�LS��q�
Do��+}Gg/��"����i�ˎ�UT��O*L���כ�Gc�-P�?%t�V�nr>�)�A��d�VYmy��|D����|ܢ/?g@&gր����C�WRV�_D�lBKɺ���O�C�Atb=�����3����!�7 άJ>�0IQ�d/�� ��k�����=/��;.� �!%ӫ���ȹk�qI�z��Fm���'�j-S�0K3t��1v���3{Ns�F�C�d]z0��%�:��a��	x��<���F]|�����x���Ͻ�iV�S�0��E�%;5�^&kr�n�@�h��hB�H�$�ס�2�t�d�:��i�6!i��zl��!J��]�JweǙA�Ђ-Z d�Rb�����)7S%u�K[��z���~|y��plF���6~�Z�	��p�9q�'�[���ⷧ���C�qr�Yٙ2�*\�b�N��� �c�:���G��%���u�~Z!7ݱ @UrD�}��IOC�:5����F�>���z�9.�!�^��qD#<Z�n�+�v�4
�C����/%w��k�)�o���c1|����g�{����:+��;d�VY������c����q��MIX6a`�]���r���2���࿻�L��d@jh�o �)��)��S"��j��=@�!HF���a��.���:����5��?_��Nʑfa|uH$_7C�o�G1�,*qq4����҅ ��aw/�����
r���i��ZN�^�xp�߼@�/��mv�����.���غ��ko���s�9oۃ���.9>�e���K���*�VYDÜ{�qՇ����Q�\&�/��i1��MK6g�_E����J+YԌ.����W�Ohx���g��G��טoh]��Z�DZ��u�]��2T��1>q��5�t�`W����'ԕ����t����ɑ�Y_�\lK^���Z�̰��Q�fλ���k��	�r���@Śo���X+�z��w�#R�P�b����������(A�9I��R��{�HЅ�%�Z|��������j�����Y�.�C�;�9�-@���ˤC6|%����/X�\��y턈�Xإ���X"8�
�c��${�=1��l����R7)?v~8��h�^~����H ���S�����&@7�ШR�|y]^��lbU*б�}����ƍ�W{�Ó�3a|5���九�*;�}<oTS!�]�*�n�L�^�Q�"�8Ȧ��R4Gi^|zG�!h.�������}?]���[���4��JKv�.�{q�`!�0��CE�:a\�l�6���E��4���st.�+���Л�	1(��w�\O��҉wJ��]�h��l����">��ZOcԅ�0\p��hW�%bڙ�#,���"�)d���la��1��;03&���+$=���mvi��%��e;[���8Oq�����9ِ�s�����*�[w����7X��^l9�Q捪��F��s_������RM(��_N��`����3���1�[� �ߠsH�޽�Mr���-J���N��s�b�E���:QЋt$2�P��0���Q�#�����B�7
M�۾)[ҫW���'�ف���_��
`;v�(��E��@f׏Dl����:G����}f�?�0������q�~-��؁�:��:�ˢBVc��eC�&_�_t�luI����Ct���@�?���2ޝD���e��L��u�ㆺa��bK�#��d�W�j����"��i��Z>մ�y3���4����`81�����mbLZ�����a1�����W��gL)�b���3̜9|�Bԝ#����v���Ts�τ��l�1ܴE�r<$�u�'�PLʰJ�[.��j�J���r�Y>Q���6\'�bv�R��SP�!��lJ�1��Jˋ��o�/�FF�R(�,�~~�H5<�c1���~�~�C3{���gt/�q�A�#�ɿVu��8L"_ύ��(�J�99�~�"1@�����O���(�4�g�f��� ��5F��W��B��"�!c?B��w�S�ߞ�Z.	����p0o�ҷFu
�	��"�!�[�F�!21�s8b��3N-܋�Nc�U����~e�����q��J=/��N��y��6j*�`H�����p�'�'\b%��i�
�w��ԙ[�����9>p�m���ds�����,}�����\���ʂN#b���<����i� �����Q�~n��g*U��F\8�z%����'*>�`4�BUBy�*ԯm�X�V�!iEg�6� ��P��/XYU䘺1B�X��g	���Չ*�L�&.�_3��,1I>�O��A��_�^��P-K�P#<N�Z��
��]~\�
��6s���^Xpn�Vz8���L\?�����}����S2�RYI��M������5rE�P����mA"�4\�۬@�v����l�;d�2(��9����4�D�V#�h�ʳ6���	)Լ�Q�����f~���}@�J0~��8&����s�O;y\����L2���}vf����N��w�oe|.�s�=�,��)s&�k�f�y؈zp�Q�*<�m�9���Q%���|�5w@dA��l�j�C�JY̸��U<\z�W�~���|_�ZbК�UV�`K�$n59W��I:�[��:iLS���Π>l}�8A3�E<�f���t����P6UH8t�fT5{�F�Cf���5CN�~ef�P�	n�-@��i8��H��X#��#��X��T_;���Ԇ�(&���--:����r-,W&����ԣ�w\`�IȔ%M�c�;923�Q��O��us@�*�ȸ� f~B,�.� ���6-L��	�I�?.Բ�`��d
A/"��_��ԗ;C����jΏTK湆8Q�rF��Kj'eTW�EX�ʝ-�H�?�����})N�גt���"���v��,~Tx���ƠJ��	��$Ɋ��/��`<˯�\~,+[�"�b���{ՆS�̊z>������0��j��t������ZK7��U�241�/ �Q��S�m{��)�T�]�ZB�R� ���G�G�< &ļ0�'����.M�ʴ����1�έ��q��&��s�w�ω�Iu��Y����ogQ�0	��p���q���I��A�(*�'�O�^�#A�h`����"g��w�����᪯�x]�r��DOWM蠪 �C֤�!�Jo��N	EO0��g_
GgԚ	-V{x�n�`O�\_p���d|�5i�Ұ��0~P��j �Ȳ&�򻑋���TN��̌%
�o�e`}��`=vr�(�?�T#Ԫl�K�)��|�';��/eM+R�-�s��D2V2�耼�KGP���/�������5g�s2��W�фܔƄ;�!�gc�i�ڛ\hؐ#c�|\���xr�V:����J�⑕�3�]HHy��iv>蝕����6fO�����}�}�7��`L{%��9�Y#\�7�VI�J�ByK��c/R����n��f����g5� S�,��s
IW�Ɲa`-Js�L�<�
Y�7)XJ��UP�U'��ch��҅d�
��iI<�/�|�%֖��IV���u� ��r�MW݂�P��:�Y`�3�T�r��g{!_��:��Ӗp�c	��M���^I(Y�D� ��.�7�/�u������lE�A~Vj1ӵǊk�/Սq�R��ׯ�̠��J�%"OF���|����N"×9�W��*��Tdgb?�0ݧ^Fu�>�A`1J�=p{.�G�q2���
����n���/�����6�]�}`��}���"Wp�`���N[Ik'	wv�� c�gt�<��������O2�a|�!��x}w�z���/�`PO��ݵ�t�m43&�@:p�="3A6�T� ����o壚-e~�1OהE`���7b?;[LK�`H�x��u�bt��lN&0�������l��y���H���l�D�Ut���(�����>���A-U� �w�( ���2v���>`a�۔�u���P!Dtw�>���<n8|����A����բ��M�hp��H����bfE%I:�䷆z�n��9ş�D�+��5�����N��V�����Cp��]&|��%�b�R�7���d�� �R���OZ�⾅���.�&{����� c�,�e�6�h�+�?q�Y�x1�c��R
�J>���J_M�� D�GpJ]�Hy�q�ȓUq�oٮ�_�3���H�ᔺ�����%�3m���y/�Fx�v�M���-^������bҞ�w��u�z��/��R��Z��Td���)�Ou��Ǻ��&