��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|̪��q[�d����0��>�����@�Q�b\~�-�X3i��ī�D�M����|��Qyc�
4�HJ+⿕����=x=�;��_N��;�Z�g��0�1�Wl}���a�K1ǘP6�R�&a1qgVZUJ���ON�Rv�շ���z��}9��"䒢½P佸WS�y����=�a=^���N� ���m3z�_�1r�����40S�����on��[4��+.n/$��>�:�]I�-�%5���kh���&��N��2i�ef;��.�OKŵ�d��B\�{w.	ѻ��\X6��)�m^�~��n���k'��p��Kцd�ג�*a���
�i�k�8zH�`��u��0�P{�5�`�0�C��o�9V�W���\��x���ñ�����כ�t�OUbH^��n�����	����q��v�:���U-6?ֿ\)o: �T��e|Ḓ��ݺ�~R/}~DZa��l�08J���|��֐4;�����tb�9Y��!L{��3���(`����1>�ڔM%�6O�y���hn�JN:�j���[�p�g	�Ԅ��N�Uk�
�lq��c��eLM��{�E*�w�_�tbbjv��꽇 2���>�)��L��H�OSg�e�l�Ƭ�M�: �ѫ����~0/5�0�v/�ʲ�e��P���ҶUr����~\�R~CLX���_ăF�g��Qf@�ϰ�6���oar9��W 3����)z���s�&F�%����"f��F�p�ͨ��ΖȹQϫ�A�.�BhO�˹+	����#��Ƃf�C��u��:�C#A�C݊W�N��ݱ��ʃ�B�r[("rTC/��-��Ew�s*-���*$�@s��pv�jj�'l��7�%����w_�fC`�Mp/Xz�"�d���|����.	t�
x�K�zI�o��tj% g3K9I3����QC0P�����YX�ū��X� �N��}��!8i�'����Ջx����\e���D��E����%Nf�ы�����:\���b��E���"��&H�M$	�f��-I�p��<�$jT	n�ó�Z(���$�s�͛"��LX�oJ�R�uHh��sJ�\\~����J��J9��=4��?��
��$�&G�)~����Iy0���k���oi�����+�����J�Q4z�nnJ�ƌ������V&6�/~�}G��;�j��Xu@
��jӽ�>� �u8�|�X?tG$h	�J��İU�'��Eq�R��*'�<*�B&\��X�m�'e�s]�ic��F�	�N�Vx����~�d*��i;E�?��`M5E*�*�1 �p&D���f2���EY�&
m�pe��n��lj�(jo�� $`w��e�zJu����:]�����?8�%��Q���l���]�#��?'���[��I�Z�v�wX_�(��0�������,.u0<>o3gо�d�	Y�����<�2�6�L6��G9����MS'c{�*�&����P2�x\�X���u�[!���8��� �6�}N$z({Z3�9W��)��>ª�Ӈ��7v�u�K"��?�=sCH5��,�l� �׫g���@?\���#N]���29FC��A�[�{w'�����T���;�3�E(�Ӑ<�g��~+N{P�J��������P�8�,~W`J˕���$�f؊.T����!>�b7p�?\ԃ�;����'��A�^�QGd#���p2W�J>��u�붚���LPC]0v�EoFz�D7=�)X��a�m����Y����7K��ېH��7�Jȗ`	��3I��_��-[L��an}`���)4�-���uD��S�nUШW�I3��*��͋������^�f��n�v���(��y?&��MI�M�)�5�%��v�������#���@(��&i�xЖ�3(c^FO�t�yfj}�Sc��O��͝�((�V�<7�*�y�s�5� ����w��q�w?|y���|�.����,FN�����t�Ϭ�]z?Ó[ �cy-)D�����j���ת�p�I��qꝾ��W.	Wkӟ��@l�N����e�׵e�A��GpLH��'�:��C�pO�b�t\�WZ��P��VMZ��s�D�&�,9��Z=�u�%>����P��'����]E�Wqȡffչ!��R#&��5�3A'E��5[��3����ֈ��b��`����S���@�g�i��5t=d3|��RY�$OIׇ�nt�g^���%���%�rW�lX>�<�����<�ʕip��X`/�-n��wd3�����<��v��x���I�S1��ډ9JMC��8I��gx�N�� >�z)^>R�i��~�-��l`���r�1v���ǫ(��[�ճ��ϽȻ�gr�Q��v���U�f�P)�^��zY}�HG�b����z��]�^���	�Y� �z�2���Hǐ*�� Y�p�dڊU�ƌ���`O�f�nmߟ���>�~�jKO��mO��^���J;2gK%QP�6�A�ɏ3���]�O.�ݵ���
��h�ܗ �Qhpi�-�:���w�A/:�!���Ec���K��N�I����n����NvB��_�������b�w��1��h}E����� 1�'�P~}e�#���zD�ջ�B�������U���0��Et^]����Q��V�]x�#;�FC/-��G$��.�?#G#6FϨ��:�L���	}1��'C�_�,�Y^�[KuM�+C_L��s$tZ���	�r����u;9L@K��۽c�A]Ը��.TxE:�>!e�(r�k��W�"bb��}OT����ҵ��3%ᇶ�9�E��מ�ᐘ�hG�\9�|���)Fz?�
\�=���|İWlqO�
)��i����e��j�=e�s�V&P��<�F1�נc���I�E��L)� ��Q��c����3ꀟ�T�h����6p�4OX�xR�4yJ�4%�Ek%��.4�y!����/�!ʇ >��N���S�\r����R�A�̖�_O� 5��~��!�-^W������@�f���w��&���{kg���q|� ��3�E-�������.��Y�"ۚN��i<����;��M+�����Ҟ��H�I��7U#@�P�w�]�Y�����W �����Aj��ߜ/����{8m�%�z���6`����B��>�ҿa'fē�nU��.{YR�ߪd�t"�! ��uO�/���\pf���^��;�4�l��y� ���i�[��?�8ziY�uܝ8�c]=�E>�w�gs� �\����8��91R�$�I�n`ݟ~ �:^
�S'<#�2v,��1=��Wu}Ɍ���ybg8v����_�Q�P�������Ev�-�=?�-�$Ei�^����r��ݠ��-����1���7���p�u���M�.����o={qzE&��ҍ�,�qуJ�eUtn��fS�#J�l�($�E���6[�����!���|ԇ��&2p���6�S�	r��-�=P4A/_$d�:X{֨��ޛ��a�@�?�93ʼ�d����Z�V�C˯p��a�f�����H��q	��1��A A*bp�s~��w8���w�8��\�tXjae���`�����|�um�r2�nOw�"�Ƒ�D�k}RԳ٨��Cr�ᬔ��7���n�q!��ْI��_a�҆�ƛ�w˄&�SzBEݝߑI~��0�(2kȕ㟬V*+�&Y+��b�t:���ip<�Zţ��1P�����}H�����5ʱ��?{�'�3���OZ��j��lq&#��2�3�'FOX�3@@TW��ϲ�:�w���s~!��ԒJ[�R��R�U�Q�Oת-ރ�E'x���T��s�%x�^�l��]�r�.�AM����Qz��S)U&J��}F��=.�> ᶸ*���Z�XY�b7����\��u��»�b樯��Xd0kw�����e���RneM恶Mt��:GR��5�D��6u��h�}���m�F}C4�<�&�C��;~a)�cY�@=�?�������*��/����o�UyT O|���25M6f��'w�	Ue`�V��j�C������)3�1�B�*𮊹V�>��~Q9-�MicH�E�
��ߖ��5�]R'�hևhʮH/���W`�W\���	���8�(:��Z��HL�e�Cǅ6���1���ie��D �u�x��2P�||��,�O�+��u3K���`�s<p���Ywu{�НH"�	��!�����IŸ�$��0u;Cs��y�af3Ob��4jv��;A�+Fh�|��֓"X�Ի�2{�y�Uk]瑳>���;�ݨ�:�BR�wU����)+��{�ݼ�,���;@�h�;�u�j��'���ؖ!��ς����,�]?�M��u���N�R�;���ڄX Ҥ9b��j��"���`m	d�q�n��*���犀�H\�ww�M��#�'���o��X�.8�n]� ?��`�K��i�f��^���T=���ͰJ2ѕ��S��ŜX��٫���C�7�q���מ�EFzV��&L�!5nkG���	�Ci'/U���� hw�#���*���8��T,��I�=���d0�l_�X<r�k�q�}���/��r2:�I���|��4o	��w�F�n�#���N�ᗇ��r��i�h<9A .��c����u��	�1�@7"|5M�:������������;�'��� W�Np$��r�D�H�B�4�$�N4������E����ݵ|7�T	ھL_�T't��A�<��9�(��^ ��d/O�[\zw�K�/Ԑ����-"��XZ�f���#|QcW�>q:�ݪ�:��r���>b}��1��Q,hF�-6�C��MR��*B+cq� �QL��c�}�;�c�o_ʄ���Ri�&�+HF�t8��z���T�,-���r��Z$Bcs�3fft>p�8+�p�G,饻�
i�I�r�+�I�z!��b��ƈ3�H�M����f1��+���d�OJܙ4Vt�wgvs�HE��]���^�7ҏ�g�f2��~���B~�ŉr�gۅ�7��?ٖ˟�3�!;��=�!�� ��k�N���j������]�|�D&-�/"�'�p8�����ї3P��	t�n�q�SƱ��H�ը��b���j��3��]�`\�S�b�d�?ׁD��y6IB�s� 腶��|\H��P���~�e����<X